
// Include register initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for register randomization.

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_
module BitLevelMaskWrite(
  input         clock,
                reset,
                needWAR,
  input  [4:0]  vd,
  output        in_0_ready,
  input         in_0_valid,
  input  [31:0] in_0_bits_data,
                in_0_bits_bitMask,
  input  [3:0]  in_0_bits_mask,
  input  [5:0]  in_0_bits_groupCounter,
  input         in_0_bits_ffoByOther,
  output        in_1_ready,
  input         in_1_valid,
  input  [31:0] in_1_bits_data,
                in_1_bits_bitMask,
  input  [3:0]  in_1_bits_mask,
  input  [5:0]  in_1_bits_groupCounter,
  input         in_1_bits_ffoByOther,
  output        in_2_ready,
  input         in_2_valid,
  input  [31:0] in_2_bits_data,
                in_2_bits_bitMask,
  input  [3:0]  in_2_bits_mask,
  input  [5:0]  in_2_bits_groupCounter,
  input         in_2_bits_ffoByOther,
  output        in_3_ready,
  input         in_3_valid,
  input  [31:0] in_3_bits_data,
                in_3_bits_bitMask,
  input  [3:0]  in_3_bits_mask,
  input  [5:0]  in_3_bits_groupCounter,
  input         in_3_bits_ffoByOther,
  output        in_4_ready,
  input         in_4_valid,
  input  [31:0] in_4_bits_data,
                in_4_bits_bitMask,
  input  [3:0]  in_4_bits_mask,
  input  [5:0]  in_4_bits_groupCounter,
  input         in_4_bits_ffoByOther,
  output        in_5_ready,
  input         in_5_valid,
  input  [31:0] in_5_bits_data,
                in_5_bits_bitMask,
  input  [3:0]  in_5_bits_mask,
  input  [5:0]  in_5_bits_groupCounter,
  input         in_5_bits_ffoByOther,
  output        in_6_ready,
  input         in_6_valid,
  input  [31:0] in_6_bits_data,
                in_6_bits_bitMask,
  input  [3:0]  in_6_bits_mask,
  input  [5:0]  in_6_bits_groupCounter,
  input         in_6_bits_ffoByOther,
  output        in_7_ready,
  input         in_7_valid,
  input  [31:0] in_7_bits_data,
                in_7_bits_bitMask,
  input  [3:0]  in_7_bits_mask,
  input  [5:0]  in_7_bits_groupCounter,
  input         in_7_bits_ffoByOther,
  output        in_8_ready,
  input         in_8_valid,
  input  [31:0] in_8_bits_data,
                in_8_bits_bitMask,
  input  [3:0]  in_8_bits_mask,
  input  [5:0]  in_8_bits_groupCounter,
  input         in_8_bits_ffoByOther,
  output        in_9_ready,
  input         in_9_valid,
  input  [31:0] in_9_bits_data,
                in_9_bits_bitMask,
  input  [3:0]  in_9_bits_mask,
  input  [5:0]  in_9_bits_groupCounter,
  input         in_9_bits_ffoByOther,
  output        in_10_ready,
  input         in_10_valid,
  input  [31:0] in_10_bits_data,
                in_10_bits_bitMask,
  input  [3:0]  in_10_bits_mask,
  input  [5:0]  in_10_bits_groupCounter,
  input         in_10_bits_ffoByOther,
  output        in_11_ready,
  input         in_11_valid,
  input  [31:0] in_11_bits_data,
                in_11_bits_bitMask,
  input  [3:0]  in_11_bits_mask,
  input  [5:0]  in_11_bits_groupCounter,
  input         in_11_bits_ffoByOther,
  output        in_12_ready,
  input         in_12_valid,
  input  [31:0] in_12_bits_data,
                in_12_bits_bitMask,
  input  [3:0]  in_12_bits_mask,
  input  [5:0]  in_12_bits_groupCounter,
  input         in_12_bits_ffoByOther,
  output        in_13_ready,
  input         in_13_valid,
  input  [31:0] in_13_bits_data,
                in_13_bits_bitMask,
  input  [3:0]  in_13_bits_mask,
  input  [5:0]  in_13_bits_groupCounter,
  input         in_13_bits_ffoByOther,
  output        in_14_ready,
  input         in_14_valid,
  input  [31:0] in_14_bits_data,
                in_14_bits_bitMask,
  input  [3:0]  in_14_bits_mask,
  input  [5:0]  in_14_bits_groupCounter,
  input         in_14_bits_ffoByOther,
  output        in_15_ready,
  input         in_15_valid,
  input  [31:0] in_15_bits_data,
                in_15_bits_bitMask,
  input  [3:0]  in_15_bits_mask,
  input  [5:0]  in_15_bits_groupCounter,
  input         in_15_bits_ffoByOther,
  output        in_16_ready,
  input         in_16_valid,
  input  [31:0] in_16_bits_data,
                in_16_bits_bitMask,
  input  [3:0]  in_16_bits_mask,
  input  [5:0]  in_16_bits_groupCounter,
  input         in_16_bits_ffoByOther,
  output        in_17_ready,
  input         in_17_valid,
  input  [31:0] in_17_bits_data,
                in_17_bits_bitMask,
  input  [3:0]  in_17_bits_mask,
  input  [5:0]  in_17_bits_groupCounter,
  input         in_17_bits_ffoByOther,
  output        in_18_ready,
  input         in_18_valid,
  input  [31:0] in_18_bits_data,
                in_18_bits_bitMask,
  input  [3:0]  in_18_bits_mask,
  input  [5:0]  in_18_bits_groupCounter,
  input         in_18_bits_ffoByOther,
  output        in_19_ready,
  input         in_19_valid,
  input  [31:0] in_19_bits_data,
                in_19_bits_bitMask,
  input  [3:0]  in_19_bits_mask,
  input  [5:0]  in_19_bits_groupCounter,
  input         in_19_bits_ffoByOther,
  output        in_20_ready,
  input         in_20_valid,
  input  [31:0] in_20_bits_data,
                in_20_bits_bitMask,
  input  [3:0]  in_20_bits_mask,
  input  [5:0]  in_20_bits_groupCounter,
  input         in_20_bits_ffoByOther,
  output        in_21_ready,
  input         in_21_valid,
  input  [31:0] in_21_bits_data,
                in_21_bits_bitMask,
  input  [3:0]  in_21_bits_mask,
  input  [5:0]  in_21_bits_groupCounter,
  input         in_21_bits_ffoByOther,
  output        in_22_ready,
  input         in_22_valid,
  input  [31:0] in_22_bits_data,
                in_22_bits_bitMask,
  input  [3:0]  in_22_bits_mask,
  input  [5:0]  in_22_bits_groupCounter,
  input         in_22_bits_ffoByOther,
  output        in_23_ready,
  input         in_23_valid,
  input  [31:0] in_23_bits_data,
                in_23_bits_bitMask,
  input  [3:0]  in_23_bits_mask,
  input  [5:0]  in_23_bits_groupCounter,
  input         in_23_bits_ffoByOther,
  output        in_24_ready,
  input         in_24_valid,
  input  [31:0] in_24_bits_data,
                in_24_bits_bitMask,
  input  [3:0]  in_24_bits_mask,
  input  [5:0]  in_24_bits_groupCounter,
  input         in_24_bits_ffoByOther,
  output        in_25_ready,
  input         in_25_valid,
  input  [31:0] in_25_bits_data,
                in_25_bits_bitMask,
  input  [3:0]  in_25_bits_mask,
  input  [5:0]  in_25_bits_groupCounter,
  input         in_25_bits_ffoByOther,
  output        in_26_ready,
  input         in_26_valid,
  input  [31:0] in_26_bits_data,
                in_26_bits_bitMask,
  input  [3:0]  in_26_bits_mask,
  input  [5:0]  in_26_bits_groupCounter,
  input         in_26_bits_ffoByOther,
  output        in_27_ready,
  input         in_27_valid,
  input  [31:0] in_27_bits_data,
                in_27_bits_bitMask,
  input  [3:0]  in_27_bits_mask,
  input  [5:0]  in_27_bits_groupCounter,
  input         in_27_bits_ffoByOther,
  output        in_28_ready,
  input         in_28_valid,
  input  [31:0] in_28_bits_data,
                in_28_bits_bitMask,
  input  [3:0]  in_28_bits_mask,
  input  [5:0]  in_28_bits_groupCounter,
  input         in_28_bits_ffoByOther,
  output        in_29_ready,
  input         in_29_valid,
  input  [31:0] in_29_bits_data,
                in_29_bits_bitMask,
  input  [3:0]  in_29_bits_mask,
  input  [5:0]  in_29_bits_groupCounter,
  input         in_29_bits_ffoByOther,
  output        in_30_ready,
  input         in_30_valid,
  input  [31:0] in_30_bits_data,
                in_30_bits_bitMask,
  input  [3:0]  in_30_bits_mask,
  input  [5:0]  in_30_bits_groupCounter,
  input         in_30_bits_ffoByOther,
  output        in_31_ready,
  input         in_31_valid,
  input  [31:0] in_31_bits_data,
                in_31_bits_bitMask,
  input  [3:0]  in_31_bits_mask,
  input  [5:0]  in_31_bits_groupCounter,
  input         in_31_bits_ffoByOther,
                out_0_ready,
  output        out_0_valid,
                out_0_bits_ffoByOther,
  output [31:0] out_0_bits_writeData_data,
  output [3:0]  out_0_bits_writeData_mask,
  output [5:0]  out_0_bits_writeData_groupCounter,
  input         out_1_ready,
  output        out_1_valid,
                out_1_bits_ffoByOther,
  output [31:0] out_1_bits_writeData_data,
  output [3:0]  out_1_bits_writeData_mask,
  output [5:0]  out_1_bits_writeData_groupCounter,
  input         out_2_ready,
  output        out_2_valid,
                out_2_bits_ffoByOther,
  output [31:0] out_2_bits_writeData_data,
  output [3:0]  out_2_bits_writeData_mask,
  output [5:0]  out_2_bits_writeData_groupCounter,
  input         out_3_ready,
  output        out_3_valid,
                out_3_bits_ffoByOther,
  output [31:0] out_3_bits_writeData_data,
  output [3:0]  out_3_bits_writeData_mask,
  output [5:0]  out_3_bits_writeData_groupCounter,
  input         out_4_ready,
  output        out_4_valid,
                out_4_bits_ffoByOther,
  output [31:0] out_4_bits_writeData_data,
  output [3:0]  out_4_bits_writeData_mask,
  output [5:0]  out_4_bits_writeData_groupCounter,
  input         out_5_ready,
  output        out_5_valid,
                out_5_bits_ffoByOther,
  output [31:0] out_5_bits_writeData_data,
  output [3:0]  out_5_bits_writeData_mask,
  output [5:0]  out_5_bits_writeData_groupCounter,
  input         out_6_ready,
  output        out_6_valid,
                out_6_bits_ffoByOther,
  output [31:0] out_6_bits_writeData_data,
  output [3:0]  out_6_bits_writeData_mask,
  output [5:0]  out_6_bits_writeData_groupCounter,
  input         out_7_ready,
  output        out_7_valid,
                out_7_bits_ffoByOther,
  output [31:0] out_7_bits_writeData_data,
  output [3:0]  out_7_bits_writeData_mask,
  output [5:0]  out_7_bits_writeData_groupCounter,
  input         out_8_ready,
  output        out_8_valid,
                out_8_bits_ffoByOther,
  output [31:0] out_8_bits_writeData_data,
  output [3:0]  out_8_bits_writeData_mask,
  output [5:0]  out_8_bits_writeData_groupCounter,
  input         out_9_ready,
  output        out_9_valid,
                out_9_bits_ffoByOther,
  output [31:0] out_9_bits_writeData_data,
  output [3:0]  out_9_bits_writeData_mask,
  output [5:0]  out_9_bits_writeData_groupCounter,
  input         out_10_ready,
  output        out_10_valid,
                out_10_bits_ffoByOther,
  output [31:0] out_10_bits_writeData_data,
  output [3:0]  out_10_bits_writeData_mask,
  output [5:0]  out_10_bits_writeData_groupCounter,
  input         out_11_ready,
  output        out_11_valid,
                out_11_bits_ffoByOther,
  output [31:0] out_11_bits_writeData_data,
  output [3:0]  out_11_bits_writeData_mask,
  output [5:0]  out_11_bits_writeData_groupCounter,
  input         out_12_ready,
  output        out_12_valid,
                out_12_bits_ffoByOther,
  output [31:0] out_12_bits_writeData_data,
  output [3:0]  out_12_bits_writeData_mask,
  output [5:0]  out_12_bits_writeData_groupCounter,
  input         out_13_ready,
  output        out_13_valid,
                out_13_bits_ffoByOther,
  output [31:0] out_13_bits_writeData_data,
  output [3:0]  out_13_bits_writeData_mask,
  output [5:0]  out_13_bits_writeData_groupCounter,
  input         out_14_ready,
  output        out_14_valid,
                out_14_bits_ffoByOther,
  output [31:0] out_14_bits_writeData_data,
  output [3:0]  out_14_bits_writeData_mask,
  output [5:0]  out_14_bits_writeData_groupCounter,
  input         out_15_ready,
  output        out_15_valid,
                out_15_bits_ffoByOther,
  output [31:0] out_15_bits_writeData_data,
  output [3:0]  out_15_bits_writeData_mask,
  output [5:0]  out_15_bits_writeData_groupCounter,
  input         out_16_ready,
  output        out_16_valid,
                out_16_bits_ffoByOther,
  output [31:0] out_16_bits_writeData_data,
  output [3:0]  out_16_bits_writeData_mask,
  output [5:0]  out_16_bits_writeData_groupCounter,
  input         out_17_ready,
  output        out_17_valid,
                out_17_bits_ffoByOther,
  output [31:0] out_17_bits_writeData_data,
  output [3:0]  out_17_bits_writeData_mask,
  output [5:0]  out_17_bits_writeData_groupCounter,
  input         out_18_ready,
  output        out_18_valid,
                out_18_bits_ffoByOther,
  output [31:0] out_18_bits_writeData_data,
  output [3:0]  out_18_bits_writeData_mask,
  output [5:0]  out_18_bits_writeData_groupCounter,
  input         out_19_ready,
  output        out_19_valid,
                out_19_bits_ffoByOther,
  output [31:0] out_19_bits_writeData_data,
  output [3:0]  out_19_bits_writeData_mask,
  output [5:0]  out_19_bits_writeData_groupCounter,
  input         out_20_ready,
  output        out_20_valid,
                out_20_bits_ffoByOther,
  output [31:0] out_20_bits_writeData_data,
  output [3:0]  out_20_bits_writeData_mask,
  output [5:0]  out_20_bits_writeData_groupCounter,
  input         out_21_ready,
  output        out_21_valid,
                out_21_bits_ffoByOther,
  output [31:0] out_21_bits_writeData_data,
  output [3:0]  out_21_bits_writeData_mask,
  output [5:0]  out_21_bits_writeData_groupCounter,
  input         out_22_ready,
  output        out_22_valid,
                out_22_bits_ffoByOther,
  output [31:0] out_22_bits_writeData_data,
  output [3:0]  out_22_bits_writeData_mask,
  output [5:0]  out_22_bits_writeData_groupCounter,
  input         out_23_ready,
  output        out_23_valid,
                out_23_bits_ffoByOther,
  output [31:0] out_23_bits_writeData_data,
  output [3:0]  out_23_bits_writeData_mask,
  output [5:0]  out_23_bits_writeData_groupCounter,
  input         out_24_ready,
  output        out_24_valid,
                out_24_bits_ffoByOther,
  output [31:0] out_24_bits_writeData_data,
  output [3:0]  out_24_bits_writeData_mask,
  output [5:0]  out_24_bits_writeData_groupCounter,
  input         out_25_ready,
  output        out_25_valid,
                out_25_bits_ffoByOther,
  output [31:0] out_25_bits_writeData_data,
  output [3:0]  out_25_bits_writeData_mask,
  output [5:0]  out_25_bits_writeData_groupCounter,
  input         out_26_ready,
  output        out_26_valid,
                out_26_bits_ffoByOther,
  output [31:0] out_26_bits_writeData_data,
  output [3:0]  out_26_bits_writeData_mask,
  output [5:0]  out_26_bits_writeData_groupCounter,
  input         out_27_ready,
  output        out_27_valid,
                out_27_bits_ffoByOther,
  output [31:0] out_27_bits_writeData_data,
  output [3:0]  out_27_bits_writeData_mask,
  output [5:0]  out_27_bits_writeData_groupCounter,
  input         out_28_ready,
  output        out_28_valid,
                out_28_bits_ffoByOther,
  output [31:0] out_28_bits_writeData_data,
  output [3:0]  out_28_bits_writeData_mask,
  output [5:0]  out_28_bits_writeData_groupCounter,
  input         out_29_ready,
  output        out_29_valid,
                out_29_bits_ffoByOther,
  output [31:0] out_29_bits_writeData_data,
  output [3:0]  out_29_bits_writeData_mask,
  output [5:0]  out_29_bits_writeData_groupCounter,
  input         out_30_ready,
  output        out_30_valid,
                out_30_bits_ffoByOther,
  output [31:0] out_30_bits_writeData_data,
  output [3:0]  out_30_bits_writeData_mask,
  output [5:0]  out_30_bits_writeData_groupCounter,
  input         out_31_ready,
  output        out_31_valid,
                out_31_bits_ffoByOther,
  output [31:0] out_31_bits_writeData_data,
  output [3:0]  out_31_bits_writeData_mask,
  output [5:0]  out_31_bits_writeData_groupCounter,
  input         readChannel_0_ready,
  output        readChannel_0_valid,
  output [4:0]  readChannel_0_bits_vs,
  output [1:0]  readChannel_0_bits_offset,
  input         readChannel_1_ready,
  output        readChannel_1_valid,
  output [4:0]  readChannel_1_bits_vs,
  output [1:0]  readChannel_1_bits_offset,
  input         readChannel_2_ready,
  output        readChannel_2_valid,
  output [4:0]  readChannel_2_bits_vs,
  output [1:0]  readChannel_2_bits_offset,
  input         readChannel_3_ready,
  output        readChannel_3_valid,
  output [4:0]  readChannel_3_bits_vs,
  output [1:0]  readChannel_3_bits_offset,
  input         readChannel_4_ready,
  output        readChannel_4_valid,
  output [4:0]  readChannel_4_bits_vs,
  output [1:0]  readChannel_4_bits_offset,
  input         readChannel_5_ready,
  output        readChannel_5_valid,
  output [4:0]  readChannel_5_bits_vs,
  output [1:0]  readChannel_5_bits_offset,
  input         readChannel_6_ready,
  output        readChannel_6_valid,
  output [4:0]  readChannel_6_bits_vs,
  output [1:0]  readChannel_6_bits_offset,
  input         readChannel_7_ready,
  output        readChannel_7_valid,
  output [4:0]  readChannel_7_bits_vs,
  output [1:0]  readChannel_7_bits_offset,
  input         readChannel_8_ready,
  output        readChannel_8_valid,
  output [4:0]  readChannel_8_bits_vs,
  output [1:0]  readChannel_8_bits_offset,
  input         readChannel_9_ready,
  output        readChannel_9_valid,
  output [4:0]  readChannel_9_bits_vs,
  output [1:0]  readChannel_9_bits_offset,
  input         readChannel_10_ready,
  output        readChannel_10_valid,
  output [4:0]  readChannel_10_bits_vs,
  output [1:0]  readChannel_10_bits_offset,
  input         readChannel_11_ready,
  output        readChannel_11_valid,
  output [4:0]  readChannel_11_bits_vs,
  output [1:0]  readChannel_11_bits_offset,
  input         readChannel_12_ready,
  output        readChannel_12_valid,
  output [4:0]  readChannel_12_bits_vs,
  output [1:0]  readChannel_12_bits_offset,
  input         readChannel_13_ready,
  output        readChannel_13_valid,
  output [4:0]  readChannel_13_bits_vs,
  output [1:0]  readChannel_13_bits_offset,
  input         readChannel_14_ready,
  output        readChannel_14_valid,
  output [4:0]  readChannel_14_bits_vs,
  output [1:0]  readChannel_14_bits_offset,
  input         readChannel_15_ready,
  output        readChannel_15_valid,
  output [4:0]  readChannel_15_bits_vs,
  output [1:0]  readChannel_15_bits_offset,
  input         readChannel_16_ready,
  output        readChannel_16_valid,
  output [4:0]  readChannel_16_bits_vs,
  output [1:0]  readChannel_16_bits_offset,
  input         readChannel_17_ready,
  output        readChannel_17_valid,
  output [4:0]  readChannel_17_bits_vs,
  output [1:0]  readChannel_17_bits_offset,
  input         readChannel_18_ready,
  output        readChannel_18_valid,
  output [4:0]  readChannel_18_bits_vs,
  output [1:0]  readChannel_18_bits_offset,
  input         readChannel_19_ready,
  output        readChannel_19_valid,
  output [4:0]  readChannel_19_bits_vs,
  output [1:0]  readChannel_19_bits_offset,
  input         readChannel_20_ready,
  output        readChannel_20_valid,
  output [4:0]  readChannel_20_bits_vs,
  output [1:0]  readChannel_20_bits_offset,
  input         readChannel_21_ready,
  output        readChannel_21_valid,
  output [4:0]  readChannel_21_bits_vs,
  output [1:0]  readChannel_21_bits_offset,
  input         readChannel_22_ready,
  output        readChannel_22_valid,
  output [4:0]  readChannel_22_bits_vs,
  output [1:0]  readChannel_22_bits_offset,
  input         readChannel_23_ready,
  output        readChannel_23_valid,
  output [4:0]  readChannel_23_bits_vs,
  output [1:0]  readChannel_23_bits_offset,
  input         readChannel_24_ready,
  output        readChannel_24_valid,
  output [4:0]  readChannel_24_bits_vs,
  output [1:0]  readChannel_24_bits_offset,
  input         readChannel_25_ready,
  output        readChannel_25_valid,
  output [4:0]  readChannel_25_bits_vs,
  output [1:0]  readChannel_25_bits_offset,
  input         readChannel_26_ready,
  output        readChannel_26_valid,
  output [4:0]  readChannel_26_bits_vs,
  output [1:0]  readChannel_26_bits_offset,
  input         readChannel_27_ready,
  output        readChannel_27_valid,
  output [4:0]  readChannel_27_bits_vs,
  output [1:0]  readChannel_27_bits_offset,
  input         readChannel_28_ready,
  output        readChannel_28_valid,
  output [4:0]  readChannel_28_bits_vs,
  output [1:0]  readChannel_28_bits_offset,
  input         readChannel_29_ready,
  output        readChannel_29_valid,
  output [4:0]  readChannel_29_bits_vs,
  output [1:0]  readChannel_29_bits_offset,
  input         readChannel_30_ready,
  output        readChannel_30_valid,
  output [4:0]  readChannel_30_bits_vs,
  output [1:0]  readChannel_30_bits_offset,
  input         readChannel_31_ready,
  output        readChannel_31_valid,
  output [4:0]  readChannel_31_bits_vs,
  output [1:0]  readChannel_31_bits_offset,
  input         readResult_0_valid,
  input  [31:0] readResult_0_bits,
  input         readResult_1_valid,
  input  [31:0] readResult_1_bits,
  input         readResult_2_valid,
  input  [31:0] readResult_2_bits,
  input         readResult_3_valid,
  input  [31:0] readResult_3_bits,
  input         readResult_4_valid,
  input  [31:0] readResult_4_bits,
  input         readResult_5_valid,
  input  [31:0] readResult_5_bits,
  input         readResult_6_valid,
  input  [31:0] readResult_6_bits,
  input         readResult_7_valid,
  input  [31:0] readResult_7_bits,
  input         readResult_8_valid,
  input  [31:0] readResult_8_bits,
  input         readResult_9_valid,
  input  [31:0] readResult_9_bits,
  input         readResult_10_valid,
  input  [31:0] readResult_10_bits,
  input         readResult_11_valid,
  input  [31:0] readResult_11_bits,
  input         readResult_12_valid,
  input  [31:0] readResult_12_bits,
  input         readResult_13_valid,
  input  [31:0] readResult_13_bits,
  input         readResult_14_valid,
  input  [31:0] readResult_14_bits,
  input         readResult_15_valid,
  input  [31:0] readResult_15_bits,
  input         readResult_16_valid,
  input  [31:0] readResult_16_bits,
  input         readResult_17_valid,
  input  [31:0] readResult_17_bits,
  input         readResult_18_valid,
  input  [31:0] readResult_18_bits,
  input         readResult_19_valid,
  input  [31:0] readResult_19_bits,
  input         readResult_20_valid,
  input  [31:0] readResult_20_bits,
  input         readResult_21_valid,
  input  [31:0] readResult_21_bits,
  input         readResult_22_valid,
  input  [31:0] readResult_22_bits,
  input         readResult_23_valid,
  input  [31:0] readResult_23_bits,
  input         readResult_24_valid,
  input  [31:0] readResult_24_bits,
  input         readResult_25_valid,
  input  [31:0] readResult_25_bits,
  input         readResult_26_valid,
  input  [31:0] readResult_26_bits,
  input         readResult_27_valid,
  input  [31:0] readResult_27_bits,
  input         readResult_28_valid,
  input  [31:0] readResult_28_bits,
  input         readResult_29_valid,
  input  [31:0] readResult_29_bits,
  input         readResult_30_valid,
  input  [31:0] readResult_30_bits,
  input         readResult_31_valid,
  input  [31:0] readResult_31_bits,
  output        stageClear
);

  wire        _stageClearVec_WaitReadQueue_fifo_31_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_31_full;
  wire        _stageClearVec_WaitReadQueue_fifo_31_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_31_data_out;
  wire        _stageClearVec_reqQueue_fifo_31_empty;
  wire        _stageClearVec_reqQueue_fifo_31_full;
  wire        _stageClearVec_reqQueue_fifo_31_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_31_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_30_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_30_full;
  wire        _stageClearVec_WaitReadQueue_fifo_30_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_30_data_out;
  wire        _stageClearVec_reqQueue_fifo_30_empty;
  wire        _stageClearVec_reqQueue_fifo_30_full;
  wire        _stageClearVec_reqQueue_fifo_30_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_30_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_29_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_29_full;
  wire        _stageClearVec_WaitReadQueue_fifo_29_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_29_data_out;
  wire        _stageClearVec_reqQueue_fifo_29_empty;
  wire        _stageClearVec_reqQueue_fifo_29_full;
  wire        _stageClearVec_reqQueue_fifo_29_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_29_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_28_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_28_full;
  wire        _stageClearVec_WaitReadQueue_fifo_28_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_28_data_out;
  wire        _stageClearVec_reqQueue_fifo_28_empty;
  wire        _stageClearVec_reqQueue_fifo_28_full;
  wire        _stageClearVec_reqQueue_fifo_28_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_28_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_27_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_27_full;
  wire        _stageClearVec_WaitReadQueue_fifo_27_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_27_data_out;
  wire        _stageClearVec_reqQueue_fifo_27_empty;
  wire        _stageClearVec_reqQueue_fifo_27_full;
  wire        _stageClearVec_reqQueue_fifo_27_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_27_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_26_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_26_full;
  wire        _stageClearVec_WaitReadQueue_fifo_26_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_26_data_out;
  wire        _stageClearVec_reqQueue_fifo_26_empty;
  wire        _stageClearVec_reqQueue_fifo_26_full;
  wire        _stageClearVec_reqQueue_fifo_26_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_26_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_25_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_25_full;
  wire        _stageClearVec_WaitReadQueue_fifo_25_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_25_data_out;
  wire        _stageClearVec_reqQueue_fifo_25_empty;
  wire        _stageClearVec_reqQueue_fifo_25_full;
  wire        _stageClearVec_reqQueue_fifo_25_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_25_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_24_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_24_full;
  wire        _stageClearVec_WaitReadQueue_fifo_24_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_24_data_out;
  wire        _stageClearVec_reqQueue_fifo_24_empty;
  wire        _stageClearVec_reqQueue_fifo_24_full;
  wire        _stageClearVec_reqQueue_fifo_24_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_24_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_23_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_23_full;
  wire        _stageClearVec_WaitReadQueue_fifo_23_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_23_data_out;
  wire        _stageClearVec_reqQueue_fifo_23_empty;
  wire        _stageClearVec_reqQueue_fifo_23_full;
  wire        _stageClearVec_reqQueue_fifo_23_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_23_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_22_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_22_full;
  wire        _stageClearVec_WaitReadQueue_fifo_22_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_22_data_out;
  wire        _stageClearVec_reqQueue_fifo_22_empty;
  wire        _stageClearVec_reqQueue_fifo_22_full;
  wire        _stageClearVec_reqQueue_fifo_22_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_22_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_21_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_21_full;
  wire        _stageClearVec_WaitReadQueue_fifo_21_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_21_data_out;
  wire        _stageClearVec_reqQueue_fifo_21_empty;
  wire        _stageClearVec_reqQueue_fifo_21_full;
  wire        _stageClearVec_reqQueue_fifo_21_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_21_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_20_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_20_full;
  wire        _stageClearVec_WaitReadQueue_fifo_20_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_20_data_out;
  wire        _stageClearVec_reqQueue_fifo_20_empty;
  wire        _stageClearVec_reqQueue_fifo_20_full;
  wire        _stageClearVec_reqQueue_fifo_20_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_20_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_19_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_19_full;
  wire        _stageClearVec_WaitReadQueue_fifo_19_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_19_data_out;
  wire        _stageClearVec_reqQueue_fifo_19_empty;
  wire        _stageClearVec_reqQueue_fifo_19_full;
  wire        _stageClearVec_reqQueue_fifo_19_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_19_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_18_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_18_full;
  wire        _stageClearVec_WaitReadQueue_fifo_18_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_18_data_out;
  wire        _stageClearVec_reqQueue_fifo_18_empty;
  wire        _stageClearVec_reqQueue_fifo_18_full;
  wire        _stageClearVec_reqQueue_fifo_18_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_18_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_17_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_17_full;
  wire        _stageClearVec_WaitReadQueue_fifo_17_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_17_data_out;
  wire        _stageClearVec_reqQueue_fifo_17_empty;
  wire        _stageClearVec_reqQueue_fifo_17_full;
  wire        _stageClearVec_reqQueue_fifo_17_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_17_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_16_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_16_full;
  wire        _stageClearVec_WaitReadQueue_fifo_16_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_16_data_out;
  wire        _stageClearVec_reqQueue_fifo_16_empty;
  wire        _stageClearVec_reqQueue_fifo_16_full;
  wire        _stageClearVec_reqQueue_fifo_16_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_16_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_15_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_15_full;
  wire        _stageClearVec_WaitReadQueue_fifo_15_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_15_data_out;
  wire        _stageClearVec_reqQueue_fifo_15_empty;
  wire        _stageClearVec_reqQueue_fifo_15_full;
  wire        _stageClearVec_reqQueue_fifo_15_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_15_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_14_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_14_full;
  wire        _stageClearVec_WaitReadQueue_fifo_14_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_14_data_out;
  wire        _stageClearVec_reqQueue_fifo_14_empty;
  wire        _stageClearVec_reqQueue_fifo_14_full;
  wire        _stageClearVec_reqQueue_fifo_14_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_14_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_13_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_13_full;
  wire        _stageClearVec_WaitReadQueue_fifo_13_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_13_data_out;
  wire        _stageClearVec_reqQueue_fifo_13_empty;
  wire        _stageClearVec_reqQueue_fifo_13_full;
  wire        _stageClearVec_reqQueue_fifo_13_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_13_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_12_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_12_full;
  wire        _stageClearVec_WaitReadQueue_fifo_12_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_12_data_out;
  wire        _stageClearVec_reqQueue_fifo_12_empty;
  wire        _stageClearVec_reqQueue_fifo_12_full;
  wire        _stageClearVec_reqQueue_fifo_12_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_12_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_11_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_11_full;
  wire        _stageClearVec_WaitReadQueue_fifo_11_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_11_data_out;
  wire        _stageClearVec_reqQueue_fifo_11_empty;
  wire        _stageClearVec_reqQueue_fifo_11_full;
  wire        _stageClearVec_reqQueue_fifo_11_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_11_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_10_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_10_full;
  wire        _stageClearVec_WaitReadQueue_fifo_10_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_10_data_out;
  wire        _stageClearVec_reqQueue_fifo_10_empty;
  wire        _stageClearVec_reqQueue_fifo_10_full;
  wire        _stageClearVec_reqQueue_fifo_10_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_10_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_9_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_9_full;
  wire        _stageClearVec_WaitReadQueue_fifo_9_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_9_data_out;
  wire        _stageClearVec_reqQueue_fifo_9_empty;
  wire        _stageClearVec_reqQueue_fifo_9_full;
  wire        _stageClearVec_reqQueue_fifo_9_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_9_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_8_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_8_full;
  wire        _stageClearVec_WaitReadQueue_fifo_8_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_8_data_out;
  wire        _stageClearVec_reqQueue_fifo_8_empty;
  wire        _stageClearVec_reqQueue_fifo_8_full;
  wire        _stageClearVec_reqQueue_fifo_8_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_8_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_7_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_7_full;
  wire        _stageClearVec_WaitReadQueue_fifo_7_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_7_data_out;
  wire        _stageClearVec_reqQueue_fifo_7_empty;
  wire        _stageClearVec_reqQueue_fifo_7_full;
  wire        _stageClearVec_reqQueue_fifo_7_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_7_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_6_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_6_full;
  wire        _stageClearVec_WaitReadQueue_fifo_6_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_6_data_out;
  wire        _stageClearVec_reqQueue_fifo_6_empty;
  wire        _stageClearVec_reqQueue_fifo_6_full;
  wire        _stageClearVec_reqQueue_fifo_6_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_6_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_5_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_5_full;
  wire        _stageClearVec_WaitReadQueue_fifo_5_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_5_data_out;
  wire        _stageClearVec_reqQueue_fifo_5_empty;
  wire        _stageClearVec_reqQueue_fifo_5_full;
  wire        _stageClearVec_reqQueue_fifo_5_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_5_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_4_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_4_full;
  wire        _stageClearVec_WaitReadQueue_fifo_4_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_4_data_out;
  wire        _stageClearVec_reqQueue_fifo_4_empty;
  wire        _stageClearVec_reqQueue_fifo_4_full;
  wire        _stageClearVec_reqQueue_fifo_4_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_4_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_3_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_3_full;
  wire        _stageClearVec_WaitReadQueue_fifo_3_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_3_data_out;
  wire        _stageClearVec_reqQueue_fifo_3_empty;
  wire        _stageClearVec_reqQueue_fifo_3_full;
  wire        _stageClearVec_reqQueue_fifo_3_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_3_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_2_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_2_full;
  wire        _stageClearVec_WaitReadQueue_fifo_2_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_2_data_out;
  wire        _stageClearVec_reqQueue_fifo_2_empty;
  wire        _stageClearVec_reqQueue_fifo_2_full;
  wire        _stageClearVec_reqQueue_fifo_2_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_2_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_1_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_1_full;
  wire        _stageClearVec_WaitReadQueue_fifo_1_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_1_data_out;
  wire        _stageClearVec_reqQueue_fifo_1_empty;
  wire        _stageClearVec_reqQueue_fifo_1_full;
  wire        _stageClearVec_reqQueue_fifo_1_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_1_data_out;
  wire        _stageClearVec_WaitReadQueue_fifo_empty;
  wire        _stageClearVec_WaitReadQueue_fifo_full;
  wire        _stageClearVec_WaitReadQueue_fifo_error;
  wire [74:0] _stageClearVec_WaitReadQueue_fifo_data_out;
  wire        _stageClearVec_reqQueue_fifo_empty;
  wire        _stageClearVec_reqQueue_fifo_full;
  wire        _stageClearVec_reqQueue_fifo_error;
  wire [74:0] _stageClearVec_reqQueue_fifo_data_out;
  wire        stageClearVec_WaitReadQueue_31_almostFull;
  wire        stageClearVec_WaitReadQueue_31_almostEmpty;
  wire        stageClearVec_reqQueue_31_almostFull;
  wire        stageClearVec_reqQueue_31_almostEmpty;
  wire        stageClearVec_WaitReadQueue_30_almostFull;
  wire        stageClearVec_WaitReadQueue_30_almostEmpty;
  wire        stageClearVec_reqQueue_30_almostFull;
  wire        stageClearVec_reqQueue_30_almostEmpty;
  wire        stageClearVec_WaitReadQueue_29_almostFull;
  wire        stageClearVec_WaitReadQueue_29_almostEmpty;
  wire        stageClearVec_reqQueue_29_almostFull;
  wire        stageClearVec_reqQueue_29_almostEmpty;
  wire        stageClearVec_WaitReadQueue_28_almostFull;
  wire        stageClearVec_WaitReadQueue_28_almostEmpty;
  wire        stageClearVec_reqQueue_28_almostFull;
  wire        stageClearVec_reqQueue_28_almostEmpty;
  wire        stageClearVec_WaitReadQueue_27_almostFull;
  wire        stageClearVec_WaitReadQueue_27_almostEmpty;
  wire        stageClearVec_reqQueue_27_almostFull;
  wire        stageClearVec_reqQueue_27_almostEmpty;
  wire        stageClearVec_WaitReadQueue_26_almostFull;
  wire        stageClearVec_WaitReadQueue_26_almostEmpty;
  wire        stageClearVec_reqQueue_26_almostFull;
  wire        stageClearVec_reqQueue_26_almostEmpty;
  wire        stageClearVec_WaitReadQueue_25_almostFull;
  wire        stageClearVec_WaitReadQueue_25_almostEmpty;
  wire        stageClearVec_reqQueue_25_almostFull;
  wire        stageClearVec_reqQueue_25_almostEmpty;
  wire        stageClearVec_WaitReadQueue_24_almostFull;
  wire        stageClearVec_WaitReadQueue_24_almostEmpty;
  wire        stageClearVec_reqQueue_24_almostFull;
  wire        stageClearVec_reqQueue_24_almostEmpty;
  wire        stageClearVec_WaitReadQueue_23_almostFull;
  wire        stageClearVec_WaitReadQueue_23_almostEmpty;
  wire        stageClearVec_reqQueue_23_almostFull;
  wire        stageClearVec_reqQueue_23_almostEmpty;
  wire        stageClearVec_WaitReadQueue_22_almostFull;
  wire        stageClearVec_WaitReadQueue_22_almostEmpty;
  wire        stageClearVec_reqQueue_22_almostFull;
  wire        stageClearVec_reqQueue_22_almostEmpty;
  wire        stageClearVec_WaitReadQueue_21_almostFull;
  wire        stageClearVec_WaitReadQueue_21_almostEmpty;
  wire        stageClearVec_reqQueue_21_almostFull;
  wire        stageClearVec_reqQueue_21_almostEmpty;
  wire        stageClearVec_WaitReadQueue_20_almostFull;
  wire        stageClearVec_WaitReadQueue_20_almostEmpty;
  wire        stageClearVec_reqQueue_20_almostFull;
  wire        stageClearVec_reqQueue_20_almostEmpty;
  wire        stageClearVec_WaitReadQueue_19_almostFull;
  wire        stageClearVec_WaitReadQueue_19_almostEmpty;
  wire        stageClearVec_reqQueue_19_almostFull;
  wire        stageClearVec_reqQueue_19_almostEmpty;
  wire        stageClearVec_WaitReadQueue_18_almostFull;
  wire        stageClearVec_WaitReadQueue_18_almostEmpty;
  wire        stageClearVec_reqQueue_18_almostFull;
  wire        stageClearVec_reqQueue_18_almostEmpty;
  wire        stageClearVec_WaitReadQueue_17_almostFull;
  wire        stageClearVec_WaitReadQueue_17_almostEmpty;
  wire        stageClearVec_reqQueue_17_almostFull;
  wire        stageClearVec_reqQueue_17_almostEmpty;
  wire        stageClearVec_WaitReadQueue_16_almostFull;
  wire        stageClearVec_WaitReadQueue_16_almostEmpty;
  wire        stageClearVec_reqQueue_16_almostFull;
  wire        stageClearVec_reqQueue_16_almostEmpty;
  wire        stageClearVec_WaitReadQueue_15_almostFull;
  wire        stageClearVec_WaitReadQueue_15_almostEmpty;
  wire        stageClearVec_reqQueue_15_almostFull;
  wire        stageClearVec_reqQueue_15_almostEmpty;
  wire        stageClearVec_WaitReadQueue_14_almostFull;
  wire        stageClearVec_WaitReadQueue_14_almostEmpty;
  wire        stageClearVec_reqQueue_14_almostFull;
  wire        stageClearVec_reqQueue_14_almostEmpty;
  wire        stageClearVec_WaitReadQueue_13_almostFull;
  wire        stageClearVec_WaitReadQueue_13_almostEmpty;
  wire        stageClearVec_reqQueue_13_almostFull;
  wire        stageClearVec_reqQueue_13_almostEmpty;
  wire        stageClearVec_WaitReadQueue_12_almostFull;
  wire        stageClearVec_WaitReadQueue_12_almostEmpty;
  wire        stageClearVec_reqQueue_12_almostFull;
  wire        stageClearVec_reqQueue_12_almostEmpty;
  wire        stageClearVec_WaitReadQueue_11_almostFull;
  wire        stageClearVec_WaitReadQueue_11_almostEmpty;
  wire        stageClearVec_reqQueue_11_almostFull;
  wire        stageClearVec_reqQueue_11_almostEmpty;
  wire        stageClearVec_WaitReadQueue_10_almostFull;
  wire        stageClearVec_WaitReadQueue_10_almostEmpty;
  wire        stageClearVec_reqQueue_10_almostFull;
  wire        stageClearVec_reqQueue_10_almostEmpty;
  wire        stageClearVec_WaitReadQueue_9_almostFull;
  wire        stageClearVec_WaitReadQueue_9_almostEmpty;
  wire        stageClearVec_reqQueue_9_almostFull;
  wire        stageClearVec_reqQueue_9_almostEmpty;
  wire        stageClearVec_WaitReadQueue_8_almostFull;
  wire        stageClearVec_WaitReadQueue_8_almostEmpty;
  wire        stageClearVec_reqQueue_8_almostFull;
  wire        stageClearVec_reqQueue_8_almostEmpty;
  wire        stageClearVec_WaitReadQueue_7_almostFull;
  wire        stageClearVec_WaitReadQueue_7_almostEmpty;
  wire        stageClearVec_reqQueue_7_almostFull;
  wire        stageClearVec_reqQueue_7_almostEmpty;
  wire        stageClearVec_WaitReadQueue_6_almostFull;
  wire        stageClearVec_WaitReadQueue_6_almostEmpty;
  wire        stageClearVec_reqQueue_6_almostFull;
  wire        stageClearVec_reqQueue_6_almostEmpty;
  wire        stageClearVec_WaitReadQueue_5_almostFull;
  wire        stageClearVec_WaitReadQueue_5_almostEmpty;
  wire        stageClearVec_reqQueue_5_almostFull;
  wire        stageClearVec_reqQueue_5_almostEmpty;
  wire        stageClearVec_WaitReadQueue_4_almostFull;
  wire        stageClearVec_WaitReadQueue_4_almostEmpty;
  wire        stageClearVec_reqQueue_4_almostFull;
  wire        stageClearVec_reqQueue_4_almostEmpty;
  wire        stageClearVec_WaitReadQueue_3_almostFull;
  wire        stageClearVec_WaitReadQueue_3_almostEmpty;
  wire        stageClearVec_reqQueue_3_almostFull;
  wire        stageClearVec_reqQueue_3_almostEmpty;
  wire        stageClearVec_WaitReadQueue_2_almostFull;
  wire        stageClearVec_WaitReadQueue_2_almostEmpty;
  wire        stageClearVec_reqQueue_2_almostFull;
  wire        stageClearVec_reqQueue_2_almostEmpty;
  wire        stageClearVec_WaitReadQueue_1_almostFull;
  wire        stageClearVec_WaitReadQueue_1_almostEmpty;
  wire        stageClearVec_reqQueue_1_almostFull;
  wire        stageClearVec_reqQueue_1_almostEmpty;
  wire        stageClearVec_WaitReadQueue_almostFull;
  wire        stageClearVec_WaitReadQueue_almostEmpty;
  wire        stageClearVec_reqQueue_almostFull;
  wire        stageClearVec_reqQueue_almostEmpty;
  wire        stageClearVec_reqQueue_31_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_31_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_31_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_31_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_31_deq_bits_data;
  wire        stageClearVec_reqQueue_30_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_30_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_30_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_30_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_30_deq_bits_data;
  wire        stageClearVec_reqQueue_29_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_29_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_29_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_29_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_29_deq_bits_data;
  wire        stageClearVec_reqQueue_28_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_28_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_28_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_28_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_28_deq_bits_data;
  wire        stageClearVec_reqQueue_27_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_27_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_27_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_27_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_27_deq_bits_data;
  wire        stageClearVec_reqQueue_26_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_26_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_26_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_26_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_26_deq_bits_data;
  wire        stageClearVec_reqQueue_25_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_25_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_25_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_25_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_25_deq_bits_data;
  wire        stageClearVec_reqQueue_24_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_24_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_24_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_24_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_24_deq_bits_data;
  wire        stageClearVec_reqQueue_23_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_23_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_23_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_23_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_23_deq_bits_data;
  wire        stageClearVec_reqQueue_22_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_22_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_22_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_22_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_22_deq_bits_data;
  wire        stageClearVec_reqQueue_21_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_21_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_21_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_21_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_21_deq_bits_data;
  wire        stageClearVec_reqQueue_20_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_20_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_20_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_20_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_20_deq_bits_data;
  wire        stageClearVec_reqQueue_19_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_19_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_19_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_19_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_19_deq_bits_data;
  wire        stageClearVec_reqQueue_18_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_18_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_18_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_18_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_18_deq_bits_data;
  wire        stageClearVec_reqQueue_17_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_17_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_17_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_17_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_17_deq_bits_data;
  wire        stageClearVec_reqQueue_16_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_16_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_16_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_16_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_16_deq_bits_data;
  wire        stageClearVec_reqQueue_15_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_15_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_15_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_15_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_15_deq_bits_data;
  wire        stageClearVec_reqQueue_14_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_14_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_14_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_14_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_14_deq_bits_data;
  wire        stageClearVec_reqQueue_13_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_13_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_13_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_13_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_13_deq_bits_data;
  wire        stageClearVec_reqQueue_12_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_12_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_12_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_12_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_12_deq_bits_data;
  wire        stageClearVec_reqQueue_11_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_11_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_11_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_11_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_11_deq_bits_data;
  wire        stageClearVec_reqQueue_10_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_10_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_10_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_10_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_10_deq_bits_data;
  wire        stageClearVec_reqQueue_9_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_9_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_9_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_9_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_9_deq_bits_data;
  wire        stageClearVec_reqQueue_8_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_8_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_8_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_8_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_8_deq_bits_data;
  wire        stageClearVec_reqQueue_7_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_7_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_7_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_7_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_7_deq_bits_data;
  wire        stageClearVec_reqQueue_6_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_6_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_6_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_6_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_6_deq_bits_data;
  wire        stageClearVec_reqQueue_5_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_5_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_5_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_5_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_5_deq_bits_data;
  wire        stageClearVec_reqQueue_4_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_4_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_4_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_4_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_4_deq_bits_data;
  wire        stageClearVec_reqQueue_3_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_3_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_3_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_3_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_3_deq_bits_data;
  wire        stageClearVec_reqQueue_2_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_2_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_2_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_2_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_2_deq_bits_data;
  wire        stageClearVec_reqQueue_1_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_1_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_1_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_1_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_1_deq_bits_data;
  wire        stageClearVec_reqQueue_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_reqQueue_deq_bits_groupCounter;
  wire [3:0]  stageClearVec_reqQueue_deq_bits_mask;
  wire [31:0] stageClearVec_reqQueue_deq_bits_bitMask;
  wire [31:0] stageClearVec_reqQueue_deq_bits_data;
  wire        in_0_valid_0 = in_0_valid;
  wire [31:0] in_0_bits_data_0 = in_0_bits_data;
  wire [31:0] in_0_bits_bitMask_0 = in_0_bits_bitMask;
  wire [3:0]  in_0_bits_mask_0 = in_0_bits_mask;
  wire [5:0]  in_0_bits_groupCounter_0 = in_0_bits_groupCounter;
  wire        in_0_bits_ffoByOther_0 = in_0_bits_ffoByOther;
  wire        in_1_valid_0 = in_1_valid;
  wire [31:0] in_1_bits_data_0 = in_1_bits_data;
  wire [31:0] in_1_bits_bitMask_0 = in_1_bits_bitMask;
  wire [3:0]  in_1_bits_mask_0 = in_1_bits_mask;
  wire [5:0]  in_1_bits_groupCounter_0 = in_1_bits_groupCounter;
  wire        in_1_bits_ffoByOther_0 = in_1_bits_ffoByOther;
  wire        in_2_valid_0 = in_2_valid;
  wire [31:0] in_2_bits_data_0 = in_2_bits_data;
  wire [31:0] in_2_bits_bitMask_0 = in_2_bits_bitMask;
  wire [3:0]  in_2_bits_mask_0 = in_2_bits_mask;
  wire [5:0]  in_2_bits_groupCounter_0 = in_2_bits_groupCounter;
  wire        in_2_bits_ffoByOther_0 = in_2_bits_ffoByOther;
  wire        in_3_valid_0 = in_3_valid;
  wire [31:0] in_3_bits_data_0 = in_3_bits_data;
  wire [31:0] in_3_bits_bitMask_0 = in_3_bits_bitMask;
  wire [3:0]  in_3_bits_mask_0 = in_3_bits_mask;
  wire [5:0]  in_3_bits_groupCounter_0 = in_3_bits_groupCounter;
  wire        in_3_bits_ffoByOther_0 = in_3_bits_ffoByOther;
  wire        in_4_valid_0 = in_4_valid;
  wire [31:0] in_4_bits_data_0 = in_4_bits_data;
  wire [31:0] in_4_bits_bitMask_0 = in_4_bits_bitMask;
  wire [3:0]  in_4_bits_mask_0 = in_4_bits_mask;
  wire [5:0]  in_4_bits_groupCounter_0 = in_4_bits_groupCounter;
  wire        in_4_bits_ffoByOther_0 = in_4_bits_ffoByOther;
  wire        in_5_valid_0 = in_5_valid;
  wire [31:0] in_5_bits_data_0 = in_5_bits_data;
  wire [31:0] in_5_bits_bitMask_0 = in_5_bits_bitMask;
  wire [3:0]  in_5_bits_mask_0 = in_5_bits_mask;
  wire [5:0]  in_5_bits_groupCounter_0 = in_5_bits_groupCounter;
  wire        in_5_bits_ffoByOther_0 = in_5_bits_ffoByOther;
  wire        in_6_valid_0 = in_6_valid;
  wire [31:0] in_6_bits_data_0 = in_6_bits_data;
  wire [31:0] in_6_bits_bitMask_0 = in_6_bits_bitMask;
  wire [3:0]  in_6_bits_mask_0 = in_6_bits_mask;
  wire [5:0]  in_6_bits_groupCounter_0 = in_6_bits_groupCounter;
  wire        in_6_bits_ffoByOther_0 = in_6_bits_ffoByOther;
  wire        in_7_valid_0 = in_7_valid;
  wire [31:0] in_7_bits_data_0 = in_7_bits_data;
  wire [31:0] in_7_bits_bitMask_0 = in_7_bits_bitMask;
  wire [3:0]  in_7_bits_mask_0 = in_7_bits_mask;
  wire [5:0]  in_7_bits_groupCounter_0 = in_7_bits_groupCounter;
  wire        in_7_bits_ffoByOther_0 = in_7_bits_ffoByOther;
  wire        in_8_valid_0 = in_8_valid;
  wire [31:0] in_8_bits_data_0 = in_8_bits_data;
  wire [31:0] in_8_bits_bitMask_0 = in_8_bits_bitMask;
  wire [3:0]  in_8_bits_mask_0 = in_8_bits_mask;
  wire [5:0]  in_8_bits_groupCounter_0 = in_8_bits_groupCounter;
  wire        in_8_bits_ffoByOther_0 = in_8_bits_ffoByOther;
  wire        in_9_valid_0 = in_9_valid;
  wire [31:0] in_9_bits_data_0 = in_9_bits_data;
  wire [31:0] in_9_bits_bitMask_0 = in_9_bits_bitMask;
  wire [3:0]  in_9_bits_mask_0 = in_9_bits_mask;
  wire [5:0]  in_9_bits_groupCounter_0 = in_9_bits_groupCounter;
  wire        in_9_bits_ffoByOther_0 = in_9_bits_ffoByOther;
  wire        in_10_valid_0 = in_10_valid;
  wire [31:0] in_10_bits_data_0 = in_10_bits_data;
  wire [31:0] in_10_bits_bitMask_0 = in_10_bits_bitMask;
  wire [3:0]  in_10_bits_mask_0 = in_10_bits_mask;
  wire [5:0]  in_10_bits_groupCounter_0 = in_10_bits_groupCounter;
  wire        in_10_bits_ffoByOther_0 = in_10_bits_ffoByOther;
  wire        in_11_valid_0 = in_11_valid;
  wire [31:0] in_11_bits_data_0 = in_11_bits_data;
  wire [31:0] in_11_bits_bitMask_0 = in_11_bits_bitMask;
  wire [3:0]  in_11_bits_mask_0 = in_11_bits_mask;
  wire [5:0]  in_11_bits_groupCounter_0 = in_11_bits_groupCounter;
  wire        in_11_bits_ffoByOther_0 = in_11_bits_ffoByOther;
  wire        in_12_valid_0 = in_12_valid;
  wire [31:0] in_12_bits_data_0 = in_12_bits_data;
  wire [31:0] in_12_bits_bitMask_0 = in_12_bits_bitMask;
  wire [3:0]  in_12_bits_mask_0 = in_12_bits_mask;
  wire [5:0]  in_12_bits_groupCounter_0 = in_12_bits_groupCounter;
  wire        in_12_bits_ffoByOther_0 = in_12_bits_ffoByOther;
  wire        in_13_valid_0 = in_13_valid;
  wire [31:0] in_13_bits_data_0 = in_13_bits_data;
  wire [31:0] in_13_bits_bitMask_0 = in_13_bits_bitMask;
  wire [3:0]  in_13_bits_mask_0 = in_13_bits_mask;
  wire [5:0]  in_13_bits_groupCounter_0 = in_13_bits_groupCounter;
  wire        in_13_bits_ffoByOther_0 = in_13_bits_ffoByOther;
  wire        in_14_valid_0 = in_14_valid;
  wire [31:0] in_14_bits_data_0 = in_14_bits_data;
  wire [31:0] in_14_bits_bitMask_0 = in_14_bits_bitMask;
  wire [3:0]  in_14_bits_mask_0 = in_14_bits_mask;
  wire [5:0]  in_14_bits_groupCounter_0 = in_14_bits_groupCounter;
  wire        in_14_bits_ffoByOther_0 = in_14_bits_ffoByOther;
  wire        in_15_valid_0 = in_15_valid;
  wire [31:0] in_15_bits_data_0 = in_15_bits_data;
  wire [31:0] in_15_bits_bitMask_0 = in_15_bits_bitMask;
  wire [3:0]  in_15_bits_mask_0 = in_15_bits_mask;
  wire [5:0]  in_15_bits_groupCounter_0 = in_15_bits_groupCounter;
  wire        in_15_bits_ffoByOther_0 = in_15_bits_ffoByOther;
  wire        in_16_valid_0 = in_16_valid;
  wire [31:0] in_16_bits_data_0 = in_16_bits_data;
  wire [31:0] in_16_bits_bitMask_0 = in_16_bits_bitMask;
  wire [3:0]  in_16_bits_mask_0 = in_16_bits_mask;
  wire [5:0]  in_16_bits_groupCounter_0 = in_16_bits_groupCounter;
  wire        in_16_bits_ffoByOther_0 = in_16_bits_ffoByOther;
  wire        in_17_valid_0 = in_17_valid;
  wire [31:0] in_17_bits_data_0 = in_17_bits_data;
  wire [31:0] in_17_bits_bitMask_0 = in_17_bits_bitMask;
  wire [3:0]  in_17_bits_mask_0 = in_17_bits_mask;
  wire [5:0]  in_17_bits_groupCounter_0 = in_17_bits_groupCounter;
  wire        in_17_bits_ffoByOther_0 = in_17_bits_ffoByOther;
  wire        in_18_valid_0 = in_18_valid;
  wire [31:0] in_18_bits_data_0 = in_18_bits_data;
  wire [31:0] in_18_bits_bitMask_0 = in_18_bits_bitMask;
  wire [3:0]  in_18_bits_mask_0 = in_18_bits_mask;
  wire [5:0]  in_18_bits_groupCounter_0 = in_18_bits_groupCounter;
  wire        in_18_bits_ffoByOther_0 = in_18_bits_ffoByOther;
  wire        in_19_valid_0 = in_19_valid;
  wire [31:0] in_19_bits_data_0 = in_19_bits_data;
  wire [31:0] in_19_bits_bitMask_0 = in_19_bits_bitMask;
  wire [3:0]  in_19_bits_mask_0 = in_19_bits_mask;
  wire [5:0]  in_19_bits_groupCounter_0 = in_19_bits_groupCounter;
  wire        in_19_bits_ffoByOther_0 = in_19_bits_ffoByOther;
  wire        in_20_valid_0 = in_20_valid;
  wire [31:0] in_20_bits_data_0 = in_20_bits_data;
  wire [31:0] in_20_bits_bitMask_0 = in_20_bits_bitMask;
  wire [3:0]  in_20_bits_mask_0 = in_20_bits_mask;
  wire [5:0]  in_20_bits_groupCounter_0 = in_20_bits_groupCounter;
  wire        in_20_bits_ffoByOther_0 = in_20_bits_ffoByOther;
  wire        in_21_valid_0 = in_21_valid;
  wire [31:0] in_21_bits_data_0 = in_21_bits_data;
  wire [31:0] in_21_bits_bitMask_0 = in_21_bits_bitMask;
  wire [3:0]  in_21_bits_mask_0 = in_21_bits_mask;
  wire [5:0]  in_21_bits_groupCounter_0 = in_21_bits_groupCounter;
  wire        in_21_bits_ffoByOther_0 = in_21_bits_ffoByOther;
  wire        in_22_valid_0 = in_22_valid;
  wire [31:0] in_22_bits_data_0 = in_22_bits_data;
  wire [31:0] in_22_bits_bitMask_0 = in_22_bits_bitMask;
  wire [3:0]  in_22_bits_mask_0 = in_22_bits_mask;
  wire [5:0]  in_22_bits_groupCounter_0 = in_22_bits_groupCounter;
  wire        in_22_bits_ffoByOther_0 = in_22_bits_ffoByOther;
  wire        in_23_valid_0 = in_23_valid;
  wire [31:0] in_23_bits_data_0 = in_23_bits_data;
  wire [31:0] in_23_bits_bitMask_0 = in_23_bits_bitMask;
  wire [3:0]  in_23_bits_mask_0 = in_23_bits_mask;
  wire [5:0]  in_23_bits_groupCounter_0 = in_23_bits_groupCounter;
  wire        in_23_bits_ffoByOther_0 = in_23_bits_ffoByOther;
  wire        in_24_valid_0 = in_24_valid;
  wire [31:0] in_24_bits_data_0 = in_24_bits_data;
  wire [31:0] in_24_bits_bitMask_0 = in_24_bits_bitMask;
  wire [3:0]  in_24_bits_mask_0 = in_24_bits_mask;
  wire [5:0]  in_24_bits_groupCounter_0 = in_24_bits_groupCounter;
  wire        in_24_bits_ffoByOther_0 = in_24_bits_ffoByOther;
  wire        in_25_valid_0 = in_25_valid;
  wire [31:0] in_25_bits_data_0 = in_25_bits_data;
  wire [31:0] in_25_bits_bitMask_0 = in_25_bits_bitMask;
  wire [3:0]  in_25_bits_mask_0 = in_25_bits_mask;
  wire [5:0]  in_25_bits_groupCounter_0 = in_25_bits_groupCounter;
  wire        in_25_bits_ffoByOther_0 = in_25_bits_ffoByOther;
  wire        in_26_valid_0 = in_26_valid;
  wire [31:0] in_26_bits_data_0 = in_26_bits_data;
  wire [31:0] in_26_bits_bitMask_0 = in_26_bits_bitMask;
  wire [3:0]  in_26_bits_mask_0 = in_26_bits_mask;
  wire [5:0]  in_26_bits_groupCounter_0 = in_26_bits_groupCounter;
  wire        in_26_bits_ffoByOther_0 = in_26_bits_ffoByOther;
  wire        in_27_valid_0 = in_27_valid;
  wire [31:0] in_27_bits_data_0 = in_27_bits_data;
  wire [31:0] in_27_bits_bitMask_0 = in_27_bits_bitMask;
  wire [3:0]  in_27_bits_mask_0 = in_27_bits_mask;
  wire [5:0]  in_27_bits_groupCounter_0 = in_27_bits_groupCounter;
  wire        in_27_bits_ffoByOther_0 = in_27_bits_ffoByOther;
  wire        in_28_valid_0 = in_28_valid;
  wire [31:0] in_28_bits_data_0 = in_28_bits_data;
  wire [31:0] in_28_bits_bitMask_0 = in_28_bits_bitMask;
  wire [3:0]  in_28_bits_mask_0 = in_28_bits_mask;
  wire [5:0]  in_28_bits_groupCounter_0 = in_28_bits_groupCounter;
  wire        in_28_bits_ffoByOther_0 = in_28_bits_ffoByOther;
  wire        in_29_valid_0 = in_29_valid;
  wire [31:0] in_29_bits_data_0 = in_29_bits_data;
  wire [31:0] in_29_bits_bitMask_0 = in_29_bits_bitMask;
  wire [3:0]  in_29_bits_mask_0 = in_29_bits_mask;
  wire [5:0]  in_29_bits_groupCounter_0 = in_29_bits_groupCounter;
  wire        in_29_bits_ffoByOther_0 = in_29_bits_ffoByOther;
  wire        in_30_valid_0 = in_30_valid;
  wire [31:0] in_30_bits_data_0 = in_30_bits_data;
  wire [31:0] in_30_bits_bitMask_0 = in_30_bits_bitMask;
  wire [3:0]  in_30_bits_mask_0 = in_30_bits_mask;
  wire [5:0]  in_30_bits_groupCounter_0 = in_30_bits_groupCounter;
  wire        in_30_bits_ffoByOther_0 = in_30_bits_ffoByOther;
  wire        in_31_valid_0 = in_31_valid;
  wire [31:0] in_31_bits_data_0 = in_31_bits_data;
  wire [31:0] in_31_bits_bitMask_0 = in_31_bits_bitMask;
  wire [3:0]  in_31_bits_mask_0 = in_31_bits_mask;
  wire [5:0]  in_31_bits_groupCounter_0 = in_31_bits_groupCounter;
  wire        in_31_bits_ffoByOther_0 = in_31_bits_ffoByOther;
  wire        out_0_ready_0 = out_0_ready;
  wire        out_1_ready_0 = out_1_ready;
  wire        out_2_ready_0 = out_2_ready;
  wire        out_3_ready_0 = out_3_ready;
  wire        out_4_ready_0 = out_4_ready;
  wire        out_5_ready_0 = out_5_ready;
  wire        out_6_ready_0 = out_6_ready;
  wire        out_7_ready_0 = out_7_ready;
  wire        out_8_ready_0 = out_8_ready;
  wire        out_9_ready_0 = out_9_ready;
  wire        out_10_ready_0 = out_10_ready;
  wire        out_11_ready_0 = out_11_ready;
  wire        out_12_ready_0 = out_12_ready;
  wire        out_13_ready_0 = out_13_ready;
  wire        out_14_ready_0 = out_14_ready;
  wire        out_15_ready_0 = out_15_ready;
  wire        out_16_ready_0 = out_16_ready;
  wire        out_17_ready_0 = out_17_ready;
  wire        out_18_ready_0 = out_18_ready;
  wire        out_19_ready_0 = out_19_ready;
  wire        out_20_ready_0 = out_20_ready;
  wire        out_21_ready_0 = out_21_ready;
  wire        out_22_ready_0 = out_22_ready;
  wire        out_23_ready_0 = out_23_ready;
  wire        out_24_ready_0 = out_24_ready;
  wire        out_25_ready_0 = out_25_ready;
  wire        out_26_ready_0 = out_26_ready;
  wire        out_27_ready_0 = out_27_ready;
  wire        out_28_ready_0 = out_28_ready;
  wire        out_29_ready_0 = out_29_ready;
  wire        out_30_ready_0 = out_30_ready;
  wire        out_31_ready_0 = out_31_ready;
  wire        readChannel_0_ready_0 = readChannel_0_ready;
  wire        readChannel_1_ready_0 = readChannel_1_ready;
  wire        readChannel_2_ready_0 = readChannel_2_ready;
  wire        readChannel_3_ready_0 = readChannel_3_ready;
  wire        readChannel_4_ready_0 = readChannel_4_ready;
  wire        readChannel_5_ready_0 = readChannel_5_ready;
  wire        readChannel_6_ready_0 = readChannel_6_ready;
  wire        readChannel_7_ready_0 = readChannel_7_ready;
  wire        readChannel_8_ready_0 = readChannel_8_ready;
  wire        readChannel_9_ready_0 = readChannel_9_ready;
  wire        readChannel_10_ready_0 = readChannel_10_ready;
  wire        readChannel_11_ready_0 = readChannel_11_ready;
  wire        readChannel_12_ready_0 = readChannel_12_ready;
  wire        readChannel_13_ready_0 = readChannel_13_ready;
  wire        readChannel_14_ready_0 = readChannel_14_ready;
  wire        readChannel_15_ready_0 = readChannel_15_ready;
  wire        readChannel_16_ready_0 = readChannel_16_ready;
  wire        readChannel_17_ready_0 = readChannel_17_ready;
  wire        readChannel_18_ready_0 = readChannel_18_ready;
  wire        readChannel_19_ready_0 = readChannel_19_ready;
  wire        readChannel_20_ready_0 = readChannel_20_ready;
  wire        readChannel_21_ready_0 = readChannel_21_ready;
  wire        readChannel_22_ready_0 = readChannel_22_ready;
  wire        readChannel_23_ready_0 = readChannel_23_ready;
  wire        readChannel_24_ready_0 = readChannel_24_ready;
  wire        readChannel_25_ready_0 = readChannel_25_ready;
  wire        readChannel_26_ready_0 = readChannel_26_ready;
  wire        readChannel_27_ready_0 = readChannel_27_ready;
  wire        readChannel_28_ready_0 = readChannel_28_ready;
  wire        readChannel_29_ready_0 = readChannel_29_ready;
  wire        readChannel_30_ready_0 = readChannel_30_ready;
  wire        readChannel_31_ready_0 = readChannel_31_ready;
  wire [1:0]  readChannel_0_bits_readSource = 2'h0;
  wire [1:0]  readChannel_1_bits_readSource = 2'h0;
  wire [1:0]  readChannel_2_bits_readSource = 2'h0;
  wire [1:0]  readChannel_3_bits_readSource = 2'h0;
  wire [1:0]  readChannel_4_bits_readSource = 2'h0;
  wire [1:0]  readChannel_5_bits_readSource = 2'h0;
  wire [1:0]  readChannel_6_bits_readSource = 2'h0;
  wire [1:0]  readChannel_7_bits_readSource = 2'h0;
  wire [1:0]  readChannel_8_bits_readSource = 2'h0;
  wire [1:0]  readChannel_9_bits_readSource = 2'h0;
  wire [1:0]  readChannel_10_bits_readSource = 2'h0;
  wire [1:0]  readChannel_11_bits_readSource = 2'h0;
  wire [1:0]  readChannel_12_bits_readSource = 2'h0;
  wire [1:0]  readChannel_13_bits_readSource = 2'h0;
  wire [1:0]  readChannel_14_bits_readSource = 2'h0;
  wire [1:0]  readChannel_15_bits_readSource = 2'h0;
  wire [1:0]  readChannel_16_bits_readSource = 2'h0;
  wire [1:0]  readChannel_17_bits_readSource = 2'h0;
  wire [1:0]  readChannel_18_bits_readSource = 2'h0;
  wire [1:0]  readChannel_19_bits_readSource = 2'h0;
  wire [1:0]  readChannel_20_bits_readSource = 2'h0;
  wire [1:0]  readChannel_21_bits_readSource = 2'h0;
  wire [1:0]  readChannel_22_bits_readSource = 2'h0;
  wire [1:0]  readChannel_23_bits_readSource = 2'h0;
  wire [1:0]  readChannel_24_bits_readSource = 2'h0;
  wire [1:0]  readChannel_25_bits_readSource = 2'h0;
  wire [1:0]  readChannel_26_bits_readSource = 2'h0;
  wire [1:0]  readChannel_27_bits_readSource = 2'h0;
  wire [1:0]  readChannel_28_bits_readSource = 2'h0;
  wire [1:0]  readChannel_29_bits_readSource = 2'h0;
  wire [1:0]  readChannel_30_bits_readSource = 2'h0;
  wire [1:0]  readChannel_31_bits_readSource = 2'h0;
  wire [2:0]  out_0_bits_index = 3'h0;
  wire [2:0]  out_1_bits_index = 3'h0;
  wire [2:0]  out_2_bits_index = 3'h0;
  wire [2:0]  out_3_bits_index = 3'h0;
  wire [2:0]  out_4_bits_index = 3'h0;
  wire [2:0]  out_5_bits_index = 3'h0;
  wire [2:0]  out_6_bits_index = 3'h0;
  wire [2:0]  out_7_bits_index = 3'h0;
  wire [2:0]  out_8_bits_index = 3'h0;
  wire [2:0]  out_9_bits_index = 3'h0;
  wire [2:0]  out_10_bits_index = 3'h0;
  wire [2:0]  out_11_bits_index = 3'h0;
  wire [2:0]  out_12_bits_index = 3'h0;
  wire [2:0]  out_13_bits_index = 3'h0;
  wire [2:0]  out_14_bits_index = 3'h0;
  wire [2:0]  out_15_bits_index = 3'h0;
  wire [2:0]  out_16_bits_index = 3'h0;
  wire [2:0]  out_17_bits_index = 3'h0;
  wire [2:0]  out_18_bits_index = 3'h0;
  wire [2:0]  out_19_bits_index = 3'h0;
  wire [2:0]  out_20_bits_index = 3'h0;
  wire [2:0]  out_21_bits_index = 3'h0;
  wire [2:0]  out_22_bits_index = 3'h0;
  wire [2:0]  out_23_bits_index = 3'h0;
  wire [2:0]  out_24_bits_index = 3'h0;
  wire [2:0]  out_25_bits_index = 3'h0;
  wire [2:0]  out_26_bits_index = 3'h0;
  wire [2:0]  out_27_bits_index = 3'h0;
  wire [2:0]  out_28_bits_index = 3'h0;
  wire [2:0]  out_29_bits_index = 3'h0;
  wire [2:0]  out_30_bits_index = 3'h0;
  wire [2:0]  out_31_bits_index = 3'h0;
  wire [2:0]  readChannel_0_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_1_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_2_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_3_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_4_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_5_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_6_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_7_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_8_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_9_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_10_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_11_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_12_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_13_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_14_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_15_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_16_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_17_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_18_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_19_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_20_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_21_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_22_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_23_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_24_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_25_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_26_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_27_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_28_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_29_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_30_bits_instructionIndex = 3'h0;
  wire [2:0]  readChannel_31_bits_instructionIndex = 3'h0;
  wire [4:0]  out_0_bits_writeData_vd = 5'h0;
  wire [4:0]  out_1_bits_writeData_vd = 5'h0;
  wire [4:0]  out_2_bits_writeData_vd = 5'h0;
  wire [4:0]  out_3_bits_writeData_vd = 5'h0;
  wire [4:0]  out_4_bits_writeData_vd = 5'h0;
  wire [4:0]  out_5_bits_writeData_vd = 5'h0;
  wire [4:0]  out_6_bits_writeData_vd = 5'h0;
  wire [4:0]  out_7_bits_writeData_vd = 5'h0;
  wire [4:0]  out_8_bits_writeData_vd = 5'h0;
  wire [4:0]  out_9_bits_writeData_vd = 5'h0;
  wire [4:0]  out_10_bits_writeData_vd = 5'h0;
  wire [4:0]  out_11_bits_writeData_vd = 5'h0;
  wire [4:0]  out_12_bits_writeData_vd = 5'h0;
  wire [4:0]  out_13_bits_writeData_vd = 5'h0;
  wire [4:0]  out_14_bits_writeData_vd = 5'h0;
  wire [4:0]  out_15_bits_writeData_vd = 5'h0;
  wire [4:0]  out_16_bits_writeData_vd = 5'h0;
  wire [4:0]  out_17_bits_writeData_vd = 5'h0;
  wire [4:0]  out_18_bits_writeData_vd = 5'h0;
  wire [4:0]  out_19_bits_writeData_vd = 5'h0;
  wire [4:0]  out_20_bits_writeData_vd = 5'h0;
  wire [4:0]  out_21_bits_writeData_vd = 5'h0;
  wire [4:0]  out_22_bits_writeData_vd = 5'h0;
  wire [4:0]  out_23_bits_writeData_vd = 5'h0;
  wire [4:0]  out_24_bits_writeData_vd = 5'h0;
  wire [4:0]  out_25_bits_writeData_vd = 5'h0;
  wire [4:0]  out_26_bits_writeData_vd = 5'h0;
  wire [4:0]  out_27_bits_writeData_vd = 5'h0;
  wire [4:0]  out_28_bits_writeData_vd = 5'h0;
  wire [4:0]  out_29_bits_writeData_vd = 5'h0;
  wire [4:0]  out_30_bits_writeData_vd = 5'h0;
  wire [4:0]  out_31_bits_writeData_vd = 5'h0;
  wire        stageClearVec_reqQueue_enq_ready;
  wire        stageClearVec_reqQueue_enq_valid = in_0_valid_0;
  wire [31:0] stageClearVec_reqQueue_enq_bits_data = in_0_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_enq_bits_bitMask = in_0_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_enq_bits_mask = in_0_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_enq_bits_groupCounter = in_0_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_enq_bits_ffoByOther = in_0_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_1_enq_ready;
  wire        stageClearVec_reqQueue_1_enq_valid = in_1_valid_0;
  wire [31:0] stageClearVec_reqQueue_1_enq_bits_data = in_1_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_1_enq_bits_bitMask = in_1_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_1_enq_bits_mask = in_1_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_1_enq_bits_groupCounter = in_1_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_1_enq_bits_ffoByOther = in_1_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_2_enq_ready;
  wire        stageClearVec_reqQueue_2_enq_valid = in_2_valid_0;
  wire [31:0] stageClearVec_reqQueue_2_enq_bits_data = in_2_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_2_enq_bits_bitMask = in_2_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_2_enq_bits_mask = in_2_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_2_enq_bits_groupCounter = in_2_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_2_enq_bits_ffoByOther = in_2_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_3_enq_ready;
  wire        stageClearVec_reqQueue_3_enq_valid = in_3_valid_0;
  wire [31:0] stageClearVec_reqQueue_3_enq_bits_data = in_3_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_3_enq_bits_bitMask = in_3_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_3_enq_bits_mask = in_3_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_3_enq_bits_groupCounter = in_3_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_3_enq_bits_ffoByOther = in_3_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_4_enq_ready;
  wire        stageClearVec_reqQueue_4_enq_valid = in_4_valid_0;
  wire [31:0] stageClearVec_reqQueue_4_enq_bits_data = in_4_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_4_enq_bits_bitMask = in_4_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_4_enq_bits_mask = in_4_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_4_enq_bits_groupCounter = in_4_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_4_enq_bits_ffoByOther = in_4_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_5_enq_ready;
  wire        stageClearVec_reqQueue_5_enq_valid = in_5_valid_0;
  wire [31:0] stageClearVec_reqQueue_5_enq_bits_data = in_5_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_5_enq_bits_bitMask = in_5_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_5_enq_bits_mask = in_5_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_5_enq_bits_groupCounter = in_5_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_5_enq_bits_ffoByOther = in_5_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_6_enq_ready;
  wire        stageClearVec_reqQueue_6_enq_valid = in_6_valid_0;
  wire [31:0] stageClearVec_reqQueue_6_enq_bits_data = in_6_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_6_enq_bits_bitMask = in_6_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_6_enq_bits_mask = in_6_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_6_enq_bits_groupCounter = in_6_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_6_enq_bits_ffoByOther = in_6_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_7_enq_ready;
  wire        stageClearVec_reqQueue_7_enq_valid = in_7_valid_0;
  wire [31:0] stageClearVec_reqQueue_7_enq_bits_data = in_7_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_7_enq_bits_bitMask = in_7_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_7_enq_bits_mask = in_7_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_7_enq_bits_groupCounter = in_7_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_7_enq_bits_ffoByOther = in_7_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_8_enq_ready;
  wire        stageClearVec_reqQueue_8_enq_valid = in_8_valid_0;
  wire [31:0] stageClearVec_reqQueue_8_enq_bits_data = in_8_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_8_enq_bits_bitMask = in_8_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_8_enq_bits_mask = in_8_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_8_enq_bits_groupCounter = in_8_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_8_enq_bits_ffoByOther = in_8_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_9_enq_ready;
  wire        stageClearVec_reqQueue_9_enq_valid = in_9_valid_0;
  wire [31:0] stageClearVec_reqQueue_9_enq_bits_data = in_9_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_9_enq_bits_bitMask = in_9_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_9_enq_bits_mask = in_9_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_9_enq_bits_groupCounter = in_9_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_9_enq_bits_ffoByOther = in_9_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_10_enq_ready;
  wire        stageClearVec_reqQueue_10_enq_valid = in_10_valid_0;
  wire [31:0] stageClearVec_reqQueue_10_enq_bits_data = in_10_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_10_enq_bits_bitMask = in_10_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_10_enq_bits_mask = in_10_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_10_enq_bits_groupCounter = in_10_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_10_enq_bits_ffoByOther = in_10_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_11_enq_ready;
  wire        stageClearVec_reqQueue_11_enq_valid = in_11_valid_0;
  wire [31:0] stageClearVec_reqQueue_11_enq_bits_data = in_11_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_11_enq_bits_bitMask = in_11_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_11_enq_bits_mask = in_11_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_11_enq_bits_groupCounter = in_11_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_11_enq_bits_ffoByOther = in_11_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_12_enq_ready;
  wire        stageClearVec_reqQueue_12_enq_valid = in_12_valid_0;
  wire [31:0] stageClearVec_reqQueue_12_enq_bits_data = in_12_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_12_enq_bits_bitMask = in_12_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_12_enq_bits_mask = in_12_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_12_enq_bits_groupCounter = in_12_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_12_enq_bits_ffoByOther = in_12_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_13_enq_ready;
  wire        stageClearVec_reqQueue_13_enq_valid = in_13_valid_0;
  wire [31:0] stageClearVec_reqQueue_13_enq_bits_data = in_13_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_13_enq_bits_bitMask = in_13_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_13_enq_bits_mask = in_13_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_13_enq_bits_groupCounter = in_13_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_13_enq_bits_ffoByOther = in_13_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_14_enq_ready;
  wire        stageClearVec_reqQueue_14_enq_valid = in_14_valid_0;
  wire [31:0] stageClearVec_reqQueue_14_enq_bits_data = in_14_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_14_enq_bits_bitMask = in_14_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_14_enq_bits_mask = in_14_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_14_enq_bits_groupCounter = in_14_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_14_enq_bits_ffoByOther = in_14_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_15_enq_ready;
  wire        stageClearVec_reqQueue_15_enq_valid = in_15_valid_0;
  wire [31:0] stageClearVec_reqQueue_15_enq_bits_data = in_15_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_15_enq_bits_bitMask = in_15_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_15_enq_bits_mask = in_15_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_15_enq_bits_groupCounter = in_15_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_15_enq_bits_ffoByOther = in_15_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_16_enq_ready;
  wire        stageClearVec_reqQueue_16_enq_valid = in_16_valid_0;
  wire [31:0] stageClearVec_reqQueue_16_enq_bits_data = in_16_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_16_enq_bits_bitMask = in_16_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_16_enq_bits_mask = in_16_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_16_enq_bits_groupCounter = in_16_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_16_enq_bits_ffoByOther = in_16_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_17_enq_ready;
  wire        stageClearVec_reqQueue_17_enq_valid = in_17_valid_0;
  wire [31:0] stageClearVec_reqQueue_17_enq_bits_data = in_17_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_17_enq_bits_bitMask = in_17_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_17_enq_bits_mask = in_17_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_17_enq_bits_groupCounter = in_17_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_17_enq_bits_ffoByOther = in_17_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_18_enq_ready;
  wire        stageClearVec_reqQueue_18_enq_valid = in_18_valid_0;
  wire [31:0] stageClearVec_reqQueue_18_enq_bits_data = in_18_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_18_enq_bits_bitMask = in_18_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_18_enq_bits_mask = in_18_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_18_enq_bits_groupCounter = in_18_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_18_enq_bits_ffoByOther = in_18_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_19_enq_ready;
  wire        stageClearVec_reqQueue_19_enq_valid = in_19_valid_0;
  wire [31:0] stageClearVec_reqQueue_19_enq_bits_data = in_19_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_19_enq_bits_bitMask = in_19_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_19_enq_bits_mask = in_19_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_19_enq_bits_groupCounter = in_19_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_19_enq_bits_ffoByOther = in_19_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_20_enq_ready;
  wire        stageClearVec_reqQueue_20_enq_valid = in_20_valid_0;
  wire [31:0] stageClearVec_reqQueue_20_enq_bits_data = in_20_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_20_enq_bits_bitMask = in_20_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_20_enq_bits_mask = in_20_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_20_enq_bits_groupCounter = in_20_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_20_enq_bits_ffoByOther = in_20_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_21_enq_ready;
  wire        stageClearVec_reqQueue_21_enq_valid = in_21_valid_0;
  wire [31:0] stageClearVec_reqQueue_21_enq_bits_data = in_21_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_21_enq_bits_bitMask = in_21_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_21_enq_bits_mask = in_21_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_21_enq_bits_groupCounter = in_21_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_21_enq_bits_ffoByOther = in_21_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_22_enq_ready;
  wire        stageClearVec_reqQueue_22_enq_valid = in_22_valid_0;
  wire [31:0] stageClearVec_reqQueue_22_enq_bits_data = in_22_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_22_enq_bits_bitMask = in_22_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_22_enq_bits_mask = in_22_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_22_enq_bits_groupCounter = in_22_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_22_enq_bits_ffoByOther = in_22_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_23_enq_ready;
  wire        stageClearVec_reqQueue_23_enq_valid = in_23_valid_0;
  wire [31:0] stageClearVec_reqQueue_23_enq_bits_data = in_23_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_23_enq_bits_bitMask = in_23_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_23_enq_bits_mask = in_23_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_23_enq_bits_groupCounter = in_23_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_23_enq_bits_ffoByOther = in_23_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_24_enq_ready;
  wire        stageClearVec_reqQueue_24_enq_valid = in_24_valid_0;
  wire [31:0] stageClearVec_reqQueue_24_enq_bits_data = in_24_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_24_enq_bits_bitMask = in_24_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_24_enq_bits_mask = in_24_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_24_enq_bits_groupCounter = in_24_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_24_enq_bits_ffoByOther = in_24_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_25_enq_ready;
  wire        stageClearVec_reqQueue_25_enq_valid = in_25_valid_0;
  wire [31:0] stageClearVec_reqQueue_25_enq_bits_data = in_25_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_25_enq_bits_bitMask = in_25_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_25_enq_bits_mask = in_25_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_25_enq_bits_groupCounter = in_25_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_25_enq_bits_ffoByOther = in_25_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_26_enq_ready;
  wire        stageClearVec_reqQueue_26_enq_valid = in_26_valid_0;
  wire [31:0] stageClearVec_reqQueue_26_enq_bits_data = in_26_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_26_enq_bits_bitMask = in_26_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_26_enq_bits_mask = in_26_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_26_enq_bits_groupCounter = in_26_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_26_enq_bits_ffoByOther = in_26_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_27_enq_ready;
  wire        stageClearVec_reqQueue_27_enq_valid = in_27_valid_0;
  wire [31:0] stageClearVec_reqQueue_27_enq_bits_data = in_27_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_27_enq_bits_bitMask = in_27_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_27_enq_bits_mask = in_27_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_27_enq_bits_groupCounter = in_27_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_27_enq_bits_ffoByOther = in_27_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_28_enq_ready;
  wire        stageClearVec_reqQueue_28_enq_valid = in_28_valid_0;
  wire [31:0] stageClearVec_reqQueue_28_enq_bits_data = in_28_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_28_enq_bits_bitMask = in_28_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_28_enq_bits_mask = in_28_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_28_enq_bits_groupCounter = in_28_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_28_enq_bits_ffoByOther = in_28_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_29_enq_ready;
  wire        stageClearVec_reqQueue_29_enq_valid = in_29_valid_0;
  wire [31:0] stageClearVec_reqQueue_29_enq_bits_data = in_29_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_29_enq_bits_bitMask = in_29_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_29_enq_bits_mask = in_29_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_29_enq_bits_groupCounter = in_29_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_29_enq_bits_ffoByOther = in_29_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_30_enq_ready;
  wire        stageClearVec_reqQueue_30_enq_valid = in_30_valid_0;
  wire [31:0] stageClearVec_reqQueue_30_enq_bits_data = in_30_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_30_enq_bits_bitMask = in_30_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_30_enq_bits_mask = in_30_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_30_enq_bits_groupCounter = in_30_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_30_enq_bits_ffoByOther = in_30_bits_ffoByOther_0;
  wire        stageClearVec_reqQueue_31_enq_ready;
  wire        stageClearVec_reqQueue_31_enq_valid = in_31_valid_0;
  wire [31:0] stageClearVec_reqQueue_31_enq_bits_data = in_31_bits_data_0;
  wire [31:0] stageClearVec_reqQueue_31_enq_bits_bitMask = in_31_bits_bitMask_0;
  wire [3:0]  stageClearVec_reqQueue_31_enq_bits_mask = in_31_bits_mask_0;
  wire [5:0]  stageClearVec_reqQueue_31_enq_bits_groupCounter = in_31_bits_groupCounter_0;
  wire        stageClearVec_reqQueue_31_enq_bits_ffoByOther = in_31_bits_ffoByOther_0;
  wire        stageClearVec_WaitReadQueue_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_1_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_1_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_2_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_2_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_3_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_3_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_4_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_4_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_5_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_5_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_6_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_6_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_7_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_7_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_8_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_8_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_9_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_9_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_10_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_10_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_11_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_11_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_12_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_12_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_13_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_13_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_14_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_14_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_15_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_15_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_16_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_16_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_17_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_17_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_18_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_18_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_19_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_19_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_20_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_20_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_21_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_21_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_22_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_22_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_23_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_23_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_24_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_24_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_25_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_25_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_26_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_26_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_27_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_27_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_28_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_28_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_29_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_29_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_30_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_30_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_31_deq_bits_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_31_deq_bits_groupCounter;
  wire        in_0_ready_0 = stageClearVec_reqQueue_enq_ready;
  wire        stageClearVec_reqQueue_deq_valid;
  assign stageClearVec_reqQueue_deq_valid = ~_stageClearVec_reqQueue_fifo_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_enq_bits_data = stageClearVec_reqQueue_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_mask;
  wire [31:0] stageClearVec_WaitReadQueue_enq_bits_bitMask = stageClearVec_reqQueue_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_enq_bits_mask = stageClearVec_reqQueue_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_enq_bits_groupCounter = stageClearVec_reqQueue_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_enq_bits_ffoByOther = stageClearVec_reqQueue_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo = {stageClearVec_reqQueue_enq_bits_groupCounter, stageClearVec_reqQueue_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi = {stageClearVec_reqQueue_enq_bits_data, stageClearVec_reqQueue_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi = {stageClearVec_reqQueue_dataIn_hi_hi, stageClearVec_reqQueue_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn = {stageClearVec_reqQueue_dataIn_hi, stageClearVec_reqQueue_dataIn_lo};
  assign stageClearVec_reqQueue_dataOut_ffoByOther = _stageClearVec_reqQueue_fifo_data_out[0];
  assign stageClearVec_reqQueue_dataOut_groupCounter = _stageClearVec_reqQueue_fifo_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_mask = _stageClearVec_reqQueue_fifo_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_bitMask = _stageClearVec_reqQueue_fifo_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_data = _stageClearVec_reqQueue_fifo_data_out[74:43];
  assign stageClearVec_reqQueue_deq_bits_data = stageClearVec_reqQueue_dataOut_data;
  assign stageClearVec_reqQueue_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_bitMask;
  assign stageClearVec_reqQueue_deq_bits_mask = stageClearVec_reqQueue_dataOut_mask;
  assign stageClearVec_reqQueue_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_groupCounter;
  assign stageClearVec_reqQueue_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_ffoByOther;
  assign stageClearVec_reqQueue_enq_ready = ~_stageClearVec_reqQueue_fifo_full;
  wire        stageClearVec_reqQueue_deq_ready;
  wire        stageClearVec_WaitReadQueue_deq_valid;
  assign stageClearVec_WaitReadQueue_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_groupCounter;
  wire [5:0]  out_0_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_ffoByOther;
  wire        out_0_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo = {stageClearVec_WaitReadQueue_enq_bits_groupCounter, stageClearVec_WaitReadQueue_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi = {stageClearVec_WaitReadQueue_enq_bits_data, stageClearVec_WaitReadQueue_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi = {stageClearVec_WaitReadQueue_dataIn_hi_hi, stageClearVec_WaitReadQueue_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn = {stageClearVec_WaitReadQueue_dataIn_hi, stageClearVec_WaitReadQueue_dataIn_lo};
  assign stageClearVec_WaitReadQueue_dataOut_ffoByOther = _stageClearVec_WaitReadQueue_fifo_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_groupCounter = _stageClearVec_WaitReadQueue_fifo_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_mask = _stageClearVec_WaitReadQueue_fifo_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_bitMask = _stageClearVec_WaitReadQueue_fifo_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_data = _stageClearVec_WaitReadQueue_fifo_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_data;
  wire [31:0] stageClearVec_WaitReadQueue_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_mask;
  assign stageClearVec_WaitReadQueue_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_groupCounter;
  assign stageClearVec_WaitReadQueue_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_ffoByOther;
  wire        stageClearVec_WaitReadQueue_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_full;
  wire        stageClearVec_WaitReadQueue_enq_valid;
  wire        stageClearVec_WaitReadQueue_deq_ready;
  wire        stageClearVec_readReady = ~needWAR | readChannel_0_ready_0;
  assign stageClearVec_WaitReadQueue_enq_valid = stageClearVec_reqQueue_deq_valid & stageClearVec_readReady;
  assign stageClearVec_reqQueue_deq_ready = stageClearVec_WaitReadQueue_enq_ready & stageClearVec_readReady;
  wire        readChannel_0_valid_0 = stageClearVec_reqQueue_deq_valid & needWAR & stageClearVec_WaitReadQueue_enq_ready;
  wire [4:0]  readChannel_0_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_0_bits_offset_0 = stageClearVec_reqQueue_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid = ~needWAR | readResult_0_valid;
  wire [31:0] stageClearVec_WARData = stageClearVec_WaitReadQueue_deq_bits_data & stageClearVec_WaitReadQueue_deq_bits_bitMask | readResult_0_bits & ~stageClearVec_WaitReadQueue_deq_bits_bitMask;
  wire        out_0_valid_0 = stageClearVec_WaitReadQueue_deq_valid & stageClearVec_readResultValid;
  assign stageClearVec_WaitReadQueue_deq_ready = out_0_ready_0 & stageClearVec_readResultValid;
  wire [31:0] out_0_bits_writeData_data_0 = needWAR ? stageClearVec_WARData : stageClearVec_WaitReadQueue_deq_bits_data;
  wire [3:0]  out_0_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter;
  wire        _stageClearVec_T = in_0_ready_0 & in_0_valid_0;
  wire [2:0]  stageClearVec_counterChange = _stageClearVec_T ? 3'h1 : 3'h7;
  wire        stageClearVec_0 = stageClearVec_counter == 3'h0;
  wire        in_1_ready_0 = stageClearVec_reqQueue_1_enq_ready;
  wire        stageClearVec_reqQueue_1_deq_valid;
  assign stageClearVec_reqQueue_1_deq_valid = ~_stageClearVec_reqQueue_fifo_1_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_1_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_1_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_1_enq_bits_data = stageClearVec_reqQueue_1_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_1_mask;
  wire [31:0] stageClearVec_WaitReadQueue_1_enq_bits_bitMask = stageClearVec_reqQueue_1_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_1_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_1_enq_bits_mask = stageClearVec_reqQueue_1_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_1_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_1_enq_bits_groupCounter = stageClearVec_reqQueue_1_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_1_enq_bits_ffoByOther = stageClearVec_reqQueue_1_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_1 = {stageClearVec_reqQueue_1_enq_bits_groupCounter, stageClearVec_reqQueue_1_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_1 = {stageClearVec_reqQueue_1_enq_bits_data, stageClearVec_reqQueue_1_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_1 = {stageClearVec_reqQueue_dataIn_hi_hi_1, stageClearVec_reqQueue_1_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_1 = {stageClearVec_reqQueue_dataIn_hi_1, stageClearVec_reqQueue_dataIn_lo_1};
  assign stageClearVec_reqQueue_dataOut_1_ffoByOther = _stageClearVec_reqQueue_fifo_1_data_out[0];
  assign stageClearVec_reqQueue_dataOut_1_groupCounter = _stageClearVec_reqQueue_fifo_1_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_1_mask = _stageClearVec_reqQueue_fifo_1_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_1_bitMask = _stageClearVec_reqQueue_fifo_1_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_1_data = _stageClearVec_reqQueue_fifo_1_data_out[74:43];
  assign stageClearVec_reqQueue_1_deq_bits_data = stageClearVec_reqQueue_dataOut_1_data;
  assign stageClearVec_reqQueue_1_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_1_bitMask;
  assign stageClearVec_reqQueue_1_deq_bits_mask = stageClearVec_reqQueue_dataOut_1_mask;
  assign stageClearVec_reqQueue_1_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_1_groupCounter;
  assign stageClearVec_reqQueue_1_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_1_ffoByOther;
  assign stageClearVec_reqQueue_1_enq_ready = ~_stageClearVec_reqQueue_fifo_1_full;
  wire        stageClearVec_reqQueue_1_deq_ready;
  wire        stageClearVec_WaitReadQueue_1_deq_valid;
  assign stageClearVec_WaitReadQueue_1_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_1_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_1_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_1_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_1_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_1_groupCounter;
  wire [5:0]  out_1_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_1_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_1_ffoByOther;
  wire        out_1_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_1_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_1 = {stageClearVec_WaitReadQueue_1_enq_bits_groupCounter, stageClearVec_WaitReadQueue_1_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_1 = {stageClearVec_WaitReadQueue_1_enq_bits_data, stageClearVec_WaitReadQueue_1_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_1 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_1, stageClearVec_WaitReadQueue_1_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_1 = {stageClearVec_WaitReadQueue_dataIn_hi_1, stageClearVec_WaitReadQueue_dataIn_lo_1};
  assign stageClearVec_WaitReadQueue_dataOut_1_ffoByOther = _stageClearVec_WaitReadQueue_fifo_1_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_1_groupCounter = _stageClearVec_WaitReadQueue_fifo_1_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_1_mask = _stageClearVec_WaitReadQueue_fifo_1_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_1_bitMask = _stageClearVec_WaitReadQueue_fifo_1_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_1_data = _stageClearVec_WaitReadQueue_fifo_1_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_1_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_1_data;
  wire [31:0] stageClearVec_WaitReadQueue_1_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_1_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_1_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_1_mask;
  assign stageClearVec_WaitReadQueue_1_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_1_groupCounter;
  assign stageClearVec_WaitReadQueue_1_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_1_ffoByOther;
  wire        stageClearVec_WaitReadQueue_1_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_1_full;
  wire        stageClearVec_WaitReadQueue_1_enq_valid;
  wire        stageClearVec_WaitReadQueue_1_deq_ready;
  wire        stageClearVec_readReady_1 = ~needWAR | readChannel_1_ready_0;
  assign stageClearVec_WaitReadQueue_1_enq_valid = stageClearVec_reqQueue_1_deq_valid & stageClearVec_readReady_1;
  assign stageClearVec_reqQueue_1_deq_ready = stageClearVec_WaitReadQueue_1_enq_ready & stageClearVec_readReady_1;
  wire        readChannel_1_valid_0 = stageClearVec_reqQueue_1_deq_valid & needWAR & stageClearVec_WaitReadQueue_1_enq_ready;
  wire [4:0]  readChannel_1_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_1_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_1_bits_offset_0 = stageClearVec_reqQueue_1_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_1 = ~needWAR | readResult_1_valid;
  wire [31:0] stageClearVec_WARData_1 = stageClearVec_WaitReadQueue_1_deq_bits_data & stageClearVec_WaitReadQueue_1_deq_bits_bitMask | readResult_1_bits & ~stageClearVec_WaitReadQueue_1_deq_bits_bitMask;
  wire        out_1_valid_0 = stageClearVec_WaitReadQueue_1_deq_valid & stageClearVec_readResultValid_1;
  assign stageClearVec_WaitReadQueue_1_deq_ready = out_1_ready_0 & stageClearVec_readResultValid_1;
  wire [31:0] out_1_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_1 : stageClearVec_WaitReadQueue_1_deq_bits_data;
  wire [3:0]  out_1_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_1_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_1;
  wire        _stageClearVec_T_3 = in_1_ready_0 & in_1_valid_0;
  wire [2:0]  stageClearVec_counterChange_1 = _stageClearVec_T_3 ? 3'h1 : 3'h7;
  wire        stageClearVec_1 = stageClearVec_counter_1 == 3'h0;
  wire        in_2_ready_0 = stageClearVec_reqQueue_2_enq_ready;
  wire        stageClearVec_reqQueue_2_deq_valid;
  assign stageClearVec_reqQueue_2_deq_valid = ~_stageClearVec_reqQueue_fifo_2_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_2_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_2_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_2_enq_bits_data = stageClearVec_reqQueue_2_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_2_mask;
  wire [31:0] stageClearVec_WaitReadQueue_2_enq_bits_bitMask = stageClearVec_reqQueue_2_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_2_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_2_enq_bits_mask = stageClearVec_reqQueue_2_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_2_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_2_enq_bits_groupCounter = stageClearVec_reqQueue_2_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_2_enq_bits_ffoByOther = stageClearVec_reqQueue_2_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_2 = {stageClearVec_reqQueue_2_enq_bits_groupCounter, stageClearVec_reqQueue_2_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_2 = {stageClearVec_reqQueue_2_enq_bits_data, stageClearVec_reqQueue_2_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_2 = {stageClearVec_reqQueue_dataIn_hi_hi_2, stageClearVec_reqQueue_2_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_2 = {stageClearVec_reqQueue_dataIn_hi_2, stageClearVec_reqQueue_dataIn_lo_2};
  assign stageClearVec_reqQueue_dataOut_2_ffoByOther = _stageClearVec_reqQueue_fifo_2_data_out[0];
  assign stageClearVec_reqQueue_dataOut_2_groupCounter = _stageClearVec_reqQueue_fifo_2_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_2_mask = _stageClearVec_reqQueue_fifo_2_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_2_bitMask = _stageClearVec_reqQueue_fifo_2_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_2_data = _stageClearVec_reqQueue_fifo_2_data_out[74:43];
  assign stageClearVec_reqQueue_2_deq_bits_data = stageClearVec_reqQueue_dataOut_2_data;
  assign stageClearVec_reqQueue_2_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_2_bitMask;
  assign stageClearVec_reqQueue_2_deq_bits_mask = stageClearVec_reqQueue_dataOut_2_mask;
  assign stageClearVec_reqQueue_2_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_2_groupCounter;
  assign stageClearVec_reqQueue_2_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_2_ffoByOther;
  assign stageClearVec_reqQueue_2_enq_ready = ~_stageClearVec_reqQueue_fifo_2_full;
  wire        stageClearVec_reqQueue_2_deq_ready;
  wire        stageClearVec_WaitReadQueue_2_deq_valid;
  assign stageClearVec_WaitReadQueue_2_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_2_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_2_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_2_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_2_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_2_groupCounter;
  wire [5:0]  out_2_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_2_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_2_ffoByOther;
  wire        out_2_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_2_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_2 = {stageClearVec_WaitReadQueue_2_enq_bits_groupCounter, stageClearVec_WaitReadQueue_2_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_2 = {stageClearVec_WaitReadQueue_2_enq_bits_data, stageClearVec_WaitReadQueue_2_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_2 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_2, stageClearVec_WaitReadQueue_2_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_2 = {stageClearVec_WaitReadQueue_dataIn_hi_2, stageClearVec_WaitReadQueue_dataIn_lo_2};
  assign stageClearVec_WaitReadQueue_dataOut_2_ffoByOther = _stageClearVec_WaitReadQueue_fifo_2_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_2_groupCounter = _stageClearVec_WaitReadQueue_fifo_2_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_2_mask = _stageClearVec_WaitReadQueue_fifo_2_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_2_bitMask = _stageClearVec_WaitReadQueue_fifo_2_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_2_data = _stageClearVec_WaitReadQueue_fifo_2_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_2_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_2_data;
  wire [31:0] stageClearVec_WaitReadQueue_2_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_2_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_2_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_2_mask;
  assign stageClearVec_WaitReadQueue_2_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_2_groupCounter;
  assign stageClearVec_WaitReadQueue_2_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_2_ffoByOther;
  wire        stageClearVec_WaitReadQueue_2_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_2_full;
  wire        stageClearVec_WaitReadQueue_2_enq_valid;
  wire        stageClearVec_WaitReadQueue_2_deq_ready;
  wire        stageClearVec_readReady_2 = ~needWAR | readChannel_2_ready_0;
  assign stageClearVec_WaitReadQueue_2_enq_valid = stageClearVec_reqQueue_2_deq_valid & stageClearVec_readReady_2;
  assign stageClearVec_reqQueue_2_deq_ready = stageClearVec_WaitReadQueue_2_enq_ready & stageClearVec_readReady_2;
  wire        readChannel_2_valid_0 = stageClearVec_reqQueue_2_deq_valid & needWAR & stageClearVec_WaitReadQueue_2_enq_ready;
  wire [4:0]  readChannel_2_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_2_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_2_bits_offset_0 = stageClearVec_reqQueue_2_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_2 = ~needWAR | readResult_2_valid;
  wire [31:0] stageClearVec_WARData_2 = stageClearVec_WaitReadQueue_2_deq_bits_data & stageClearVec_WaitReadQueue_2_deq_bits_bitMask | readResult_2_bits & ~stageClearVec_WaitReadQueue_2_deq_bits_bitMask;
  wire        out_2_valid_0 = stageClearVec_WaitReadQueue_2_deq_valid & stageClearVec_readResultValid_2;
  assign stageClearVec_WaitReadQueue_2_deq_ready = out_2_ready_0 & stageClearVec_readResultValid_2;
  wire [31:0] out_2_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_2 : stageClearVec_WaitReadQueue_2_deq_bits_data;
  wire [3:0]  out_2_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_2_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_2;
  wire        _stageClearVec_T_6 = in_2_ready_0 & in_2_valid_0;
  wire [2:0]  stageClearVec_counterChange_2 = _stageClearVec_T_6 ? 3'h1 : 3'h7;
  wire        stageClearVec_2 = stageClearVec_counter_2 == 3'h0;
  wire        in_3_ready_0 = stageClearVec_reqQueue_3_enq_ready;
  wire        stageClearVec_reqQueue_3_deq_valid;
  assign stageClearVec_reqQueue_3_deq_valid = ~_stageClearVec_reqQueue_fifo_3_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_3_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_3_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_3_enq_bits_data = stageClearVec_reqQueue_3_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_3_mask;
  wire [31:0] stageClearVec_WaitReadQueue_3_enq_bits_bitMask = stageClearVec_reqQueue_3_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_3_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_3_enq_bits_mask = stageClearVec_reqQueue_3_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_3_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_3_enq_bits_groupCounter = stageClearVec_reqQueue_3_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_3_enq_bits_ffoByOther = stageClearVec_reqQueue_3_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_3 = {stageClearVec_reqQueue_3_enq_bits_groupCounter, stageClearVec_reqQueue_3_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_3 = {stageClearVec_reqQueue_3_enq_bits_data, stageClearVec_reqQueue_3_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_3 = {stageClearVec_reqQueue_dataIn_hi_hi_3, stageClearVec_reqQueue_3_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_3 = {stageClearVec_reqQueue_dataIn_hi_3, stageClearVec_reqQueue_dataIn_lo_3};
  assign stageClearVec_reqQueue_dataOut_3_ffoByOther = _stageClearVec_reqQueue_fifo_3_data_out[0];
  assign stageClearVec_reqQueue_dataOut_3_groupCounter = _stageClearVec_reqQueue_fifo_3_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_3_mask = _stageClearVec_reqQueue_fifo_3_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_3_bitMask = _stageClearVec_reqQueue_fifo_3_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_3_data = _stageClearVec_reqQueue_fifo_3_data_out[74:43];
  assign stageClearVec_reqQueue_3_deq_bits_data = stageClearVec_reqQueue_dataOut_3_data;
  assign stageClearVec_reqQueue_3_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_3_bitMask;
  assign stageClearVec_reqQueue_3_deq_bits_mask = stageClearVec_reqQueue_dataOut_3_mask;
  assign stageClearVec_reqQueue_3_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_3_groupCounter;
  assign stageClearVec_reqQueue_3_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_3_ffoByOther;
  assign stageClearVec_reqQueue_3_enq_ready = ~_stageClearVec_reqQueue_fifo_3_full;
  wire        stageClearVec_reqQueue_3_deq_ready;
  wire        stageClearVec_WaitReadQueue_3_deq_valid;
  assign stageClearVec_WaitReadQueue_3_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_3_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_3_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_3_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_3_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_3_groupCounter;
  wire [5:0]  out_3_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_3_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_3_ffoByOther;
  wire        out_3_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_3_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_3 = {stageClearVec_WaitReadQueue_3_enq_bits_groupCounter, stageClearVec_WaitReadQueue_3_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_3 = {stageClearVec_WaitReadQueue_3_enq_bits_data, stageClearVec_WaitReadQueue_3_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_3 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_3, stageClearVec_WaitReadQueue_3_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_3 = {stageClearVec_WaitReadQueue_dataIn_hi_3, stageClearVec_WaitReadQueue_dataIn_lo_3};
  assign stageClearVec_WaitReadQueue_dataOut_3_ffoByOther = _stageClearVec_WaitReadQueue_fifo_3_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_3_groupCounter = _stageClearVec_WaitReadQueue_fifo_3_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_3_mask = _stageClearVec_WaitReadQueue_fifo_3_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_3_bitMask = _stageClearVec_WaitReadQueue_fifo_3_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_3_data = _stageClearVec_WaitReadQueue_fifo_3_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_3_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_3_data;
  wire [31:0] stageClearVec_WaitReadQueue_3_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_3_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_3_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_3_mask;
  assign stageClearVec_WaitReadQueue_3_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_3_groupCounter;
  assign stageClearVec_WaitReadQueue_3_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_3_ffoByOther;
  wire        stageClearVec_WaitReadQueue_3_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_3_full;
  wire        stageClearVec_WaitReadQueue_3_enq_valid;
  wire        stageClearVec_WaitReadQueue_3_deq_ready;
  wire        stageClearVec_readReady_3 = ~needWAR | readChannel_3_ready_0;
  assign stageClearVec_WaitReadQueue_3_enq_valid = stageClearVec_reqQueue_3_deq_valid & stageClearVec_readReady_3;
  assign stageClearVec_reqQueue_3_deq_ready = stageClearVec_WaitReadQueue_3_enq_ready & stageClearVec_readReady_3;
  wire        readChannel_3_valid_0 = stageClearVec_reqQueue_3_deq_valid & needWAR & stageClearVec_WaitReadQueue_3_enq_ready;
  wire [4:0]  readChannel_3_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_3_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_3_bits_offset_0 = stageClearVec_reqQueue_3_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_3 = ~needWAR | readResult_3_valid;
  wire [31:0] stageClearVec_WARData_3 = stageClearVec_WaitReadQueue_3_deq_bits_data & stageClearVec_WaitReadQueue_3_deq_bits_bitMask | readResult_3_bits & ~stageClearVec_WaitReadQueue_3_deq_bits_bitMask;
  wire        out_3_valid_0 = stageClearVec_WaitReadQueue_3_deq_valid & stageClearVec_readResultValid_3;
  assign stageClearVec_WaitReadQueue_3_deq_ready = out_3_ready_0 & stageClearVec_readResultValid_3;
  wire [31:0] out_3_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_3 : stageClearVec_WaitReadQueue_3_deq_bits_data;
  wire [3:0]  out_3_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_3_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_3;
  wire        _stageClearVec_T_9 = in_3_ready_0 & in_3_valid_0;
  wire [2:0]  stageClearVec_counterChange_3 = _stageClearVec_T_9 ? 3'h1 : 3'h7;
  wire        stageClearVec_3 = stageClearVec_counter_3 == 3'h0;
  wire        in_4_ready_0 = stageClearVec_reqQueue_4_enq_ready;
  wire        stageClearVec_reqQueue_4_deq_valid;
  assign stageClearVec_reqQueue_4_deq_valid = ~_stageClearVec_reqQueue_fifo_4_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_4_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_4_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_4_enq_bits_data = stageClearVec_reqQueue_4_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_4_mask;
  wire [31:0] stageClearVec_WaitReadQueue_4_enq_bits_bitMask = stageClearVec_reqQueue_4_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_4_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_4_enq_bits_mask = stageClearVec_reqQueue_4_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_4_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_4_enq_bits_groupCounter = stageClearVec_reqQueue_4_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_4_enq_bits_ffoByOther = stageClearVec_reqQueue_4_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_4 = {stageClearVec_reqQueue_4_enq_bits_groupCounter, stageClearVec_reqQueue_4_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_4 = {stageClearVec_reqQueue_4_enq_bits_data, stageClearVec_reqQueue_4_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_4 = {stageClearVec_reqQueue_dataIn_hi_hi_4, stageClearVec_reqQueue_4_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_4 = {stageClearVec_reqQueue_dataIn_hi_4, stageClearVec_reqQueue_dataIn_lo_4};
  assign stageClearVec_reqQueue_dataOut_4_ffoByOther = _stageClearVec_reqQueue_fifo_4_data_out[0];
  assign stageClearVec_reqQueue_dataOut_4_groupCounter = _stageClearVec_reqQueue_fifo_4_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_4_mask = _stageClearVec_reqQueue_fifo_4_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_4_bitMask = _stageClearVec_reqQueue_fifo_4_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_4_data = _stageClearVec_reqQueue_fifo_4_data_out[74:43];
  assign stageClearVec_reqQueue_4_deq_bits_data = stageClearVec_reqQueue_dataOut_4_data;
  assign stageClearVec_reqQueue_4_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_4_bitMask;
  assign stageClearVec_reqQueue_4_deq_bits_mask = stageClearVec_reqQueue_dataOut_4_mask;
  assign stageClearVec_reqQueue_4_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_4_groupCounter;
  assign stageClearVec_reqQueue_4_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_4_ffoByOther;
  assign stageClearVec_reqQueue_4_enq_ready = ~_stageClearVec_reqQueue_fifo_4_full;
  wire        stageClearVec_reqQueue_4_deq_ready;
  wire        stageClearVec_WaitReadQueue_4_deq_valid;
  assign stageClearVec_WaitReadQueue_4_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_4_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_4_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_4_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_4_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_4_groupCounter;
  wire [5:0]  out_4_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_4_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_4_ffoByOther;
  wire        out_4_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_4_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_4 = {stageClearVec_WaitReadQueue_4_enq_bits_groupCounter, stageClearVec_WaitReadQueue_4_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_4 = {stageClearVec_WaitReadQueue_4_enq_bits_data, stageClearVec_WaitReadQueue_4_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_4 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_4, stageClearVec_WaitReadQueue_4_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_4 = {stageClearVec_WaitReadQueue_dataIn_hi_4, stageClearVec_WaitReadQueue_dataIn_lo_4};
  assign stageClearVec_WaitReadQueue_dataOut_4_ffoByOther = _stageClearVec_WaitReadQueue_fifo_4_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_4_groupCounter = _stageClearVec_WaitReadQueue_fifo_4_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_4_mask = _stageClearVec_WaitReadQueue_fifo_4_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_4_bitMask = _stageClearVec_WaitReadQueue_fifo_4_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_4_data = _stageClearVec_WaitReadQueue_fifo_4_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_4_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_4_data;
  wire [31:0] stageClearVec_WaitReadQueue_4_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_4_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_4_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_4_mask;
  assign stageClearVec_WaitReadQueue_4_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_4_groupCounter;
  assign stageClearVec_WaitReadQueue_4_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_4_ffoByOther;
  wire        stageClearVec_WaitReadQueue_4_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_4_full;
  wire        stageClearVec_WaitReadQueue_4_enq_valid;
  wire        stageClearVec_WaitReadQueue_4_deq_ready;
  wire        stageClearVec_readReady_4 = ~needWAR | readChannel_4_ready_0;
  assign stageClearVec_WaitReadQueue_4_enq_valid = stageClearVec_reqQueue_4_deq_valid & stageClearVec_readReady_4;
  assign stageClearVec_reqQueue_4_deq_ready = stageClearVec_WaitReadQueue_4_enq_ready & stageClearVec_readReady_4;
  wire        readChannel_4_valid_0 = stageClearVec_reqQueue_4_deq_valid & needWAR & stageClearVec_WaitReadQueue_4_enq_ready;
  wire [4:0]  readChannel_4_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_4_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_4_bits_offset_0 = stageClearVec_reqQueue_4_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_4 = ~needWAR | readResult_4_valid;
  wire [31:0] stageClearVec_WARData_4 = stageClearVec_WaitReadQueue_4_deq_bits_data & stageClearVec_WaitReadQueue_4_deq_bits_bitMask | readResult_4_bits & ~stageClearVec_WaitReadQueue_4_deq_bits_bitMask;
  wire        out_4_valid_0 = stageClearVec_WaitReadQueue_4_deq_valid & stageClearVec_readResultValid_4;
  assign stageClearVec_WaitReadQueue_4_deq_ready = out_4_ready_0 & stageClearVec_readResultValid_4;
  wire [31:0] out_4_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_4 : stageClearVec_WaitReadQueue_4_deq_bits_data;
  wire [3:0]  out_4_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_4_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_4;
  wire        _stageClearVec_T_12 = in_4_ready_0 & in_4_valid_0;
  wire [2:0]  stageClearVec_counterChange_4 = _stageClearVec_T_12 ? 3'h1 : 3'h7;
  wire        stageClearVec_4 = stageClearVec_counter_4 == 3'h0;
  wire        in_5_ready_0 = stageClearVec_reqQueue_5_enq_ready;
  wire        stageClearVec_reqQueue_5_deq_valid;
  assign stageClearVec_reqQueue_5_deq_valid = ~_stageClearVec_reqQueue_fifo_5_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_5_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_5_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_5_enq_bits_data = stageClearVec_reqQueue_5_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_5_mask;
  wire [31:0] stageClearVec_WaitReadQueue_5_enq_bits_bitMask = stageClearVec_reqQueue_5_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_5_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_5_enq_bits_mask = stageClearVec_reqQueue_5_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_5_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_5_enq_bits_groupCounter = stageClearVec_reqQueue_5_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_5_enq_bits_ffoByOther = stageClearVec_reqQueue_5_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_5 = {stageClearVec_reqQueue_5_enq_bits_groupCounter, stageClearVec_reqQueue_5_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_5 = {stageClearVec_reqQueue_5_enq_bits_data, stageClearVec_reqQueue_5_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_5 = {stageClearVec_reqQueue_dataIn_hi_hi_5, stageClearVec_reqQueue_5_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_5 = {stageClearVec_reqQueue_dataIn_hi_5, stageClearVec_reqQueue_dataIn_lo_5};
  assign stageClearVec_reqQueue_dataOut_5_ffoByOther = _stageClearVec_reqQueue_fifo_5_data_out[0];
  assign stageClearVec_reqQueue_dataOut_5_groupCounter = _stageClearVec_reqQueue_fifo_5_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_5_mask = _stageClearVec_reqQueue_fifo_5_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_5_bitMask = _stageClearVec_reqQueue_fifo_5_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_5_data = _stageClearVec_reqQueue_fifo_5_data_out[74:43];
  assign stageClearVec_reqQueue_5_deq_bits_data = stageClearVec_reqQueue_dataOut_5_data;
  assign stageClearVec_reqQueue_5_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_5_bitMask;
  assign stageClearVec_reqQueue_5_deq_bits_mask = stageClearVec_reqQueue_dataOut_5_mask;
  assign stageClearVec_reqQueue_5_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_5_groupCounter;
  assign stageClearVec_reqQueue_5_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_5_ffoByOther;
  assign stageClearVec_reqQueue_5_enq_ready = ~_stageClearVec_reqQueue_fifo_5_full;
  wire        stageClearVec_reqQueue_5_deq_ready;
  wire        stageClearVec_WaitReadQueue_5_deq_valid;
  assign stageClearVec_WaitReadQueue_5_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_5_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_5_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_5_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_5_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_5_groupCounter;
  wire [5:0]  out_5_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_5_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_5_ffoByOther;
  wire        out_5_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_5_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_5 = {stageClearVec_WaitReadQueue_5_enq_bits_groupCounter, stageClearVec_WaitReadQueue_5_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_5 = {stageClearVec_WaitReadQueue_5_enq_bits_data, stageClearVec_WaitReadQueue_5_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_5 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_5, stageClearVec_WaitReadQueue_5_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_5 = {stageClearVec_WaitReadQueue_dataIn_hi_5, stageClearVec_WaitReadQueue_dataIn_lo_5};
  assign stageClearVec_WaitReadQueue_dataOut_5_ffoByOther = _stageClearVec_WaitReadQueue_fifo_5_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_5_groupCounter = _stageClearVec_WaitReadQueue_fifo_5_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_5_mask = _stageClearVec_WaitReadQueue_fifo_5_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_5_bitMask = _stageClearVec_WaitReadQueue_fifo_5_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_5_data = _stageClearVec_WaitReadQueue_fifo_5_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_5_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_5_data;
  wire [31:0] stageClearVec_WaitReadQueue_5_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_5_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_5_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_5_mask;
  assign stageClearVec_WaitReadQueue_5_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_5_groupCounter;
  assign stageClearVec_WaitReadQueue_5_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_5_ffoByOther;
  wire        stageClearVec_WaitReadQueue_5_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_5_full;
  wire        stageClearVec_WaitReadQueue_5_enq_valid;
  wire        stageClearVec_WaitReadQueue_5_deq_ready;
  wire        stageClearVec_readReady_5 = ~needWAR | readChannel_5_ready_0;
  assign stageClearVec_WaitReadQueue_5_enq_valid = stageClearVec_reqQueue_5_deq_valid & stageClearVec_readReady_5;
  assign stageClearVec_reqQueue_5_deq_ready = stageClearVec_WaitReadQueue_5_enq_ready & stageClearVec_readReady_5;
  wire        readChannel_5_valid_0 = stageClearVec_reqQueue_5_deq_valid & needWAR & stageClearVec_WaitReadQueue_5_enq_ready;
  wire [4:0]  readChannel_5_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_5_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_5_bits_offset_0 = stageClearVec_reqQueue_5_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_5 = ~needWAR | readResult_5_valid;
  wire [31:0] stageClearVec_WARData_5 = stageClearVec_WaitReadQueue_5_deq_bits_data & stageClearVec_WaitReadQueue_5_deq_bits_bitMask | readResult_5_bits & ~stageClearVec_WaitReadQueue_5_deq_bits_bitMask;
  wire        out_5_valid_0 = stageClearVec_WaitReadQueue_5_deq_valid & stageClearVec_readResultValid_5;
  assign stageClearVec_WaitReadQueue_5_deq_ready = out_5_ready_0 & stageClearVec_readResultValid_5;
  wire [31:0] out_5_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_5 : stageClearVec_WaitReadQueue_5_deq_bits_data;
  wire [3:0]  out_5_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_5_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_5;
  wire        _stageClearVec_T_15 = in_5_ready_0 & in_5_valid_0;
  wire [2:0]  stageClearVec_counterChange_5 = _stageClearVec_T_15 ? 3'h1 : 3'h7;
  wire        stageClearVec_5 = stageClearVec_counter_5 == 3'h0;
  wire        in_6_ready_0 = stageClearVec_reqQueue_6_enq_ready;
  wire        stageClearVec_reqQueue_6_deq_valid;
  assign stageClearVec_reqQueue_6_deq_valid = ~_stageClearVec_reqQueue_fifo_6_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_6_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_6_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_6_enq_bits_data = stageClearVec_reqQueue_6_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_6_mask;
  wire [31:0] stageClearVec_WaitReadQueue_6_enq_bits_bitMask = stageClearVec_reqQueue_6_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_6_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_6_enq_bits_mask = stageClearVec_reqQueue_6_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_6_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_6_enq_bits_groupCounter = stageClearVec_reqQueue_6_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_6_enq_bits_ffoByOther = stageClearVec_reqQueue_6_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_6 = {stageClearVec_reqQueue_6_enq_bits_groupCounter, stageClearVec_reqQueue_6_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_6 = {stageClearVec_reqQueue_6_enq_bits_data, stageClearVec_reqQueue_6_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_6 = {stageClearVec_reqQueue_dataIn_hi_hi_6, stageClearVec_reqQueue_6_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_6 = {stageClearVec_reqQueue_dataIn_hi_6, stageClearVec_reqQueue_dataIn_lo_6};
  assign stageClearVec_reqQueue_dataOut_6_ffoByOther = _stageClearVec_reqQueue_fifo_6_data_out[0];
  assign stageClearVec_reqQueue_dataOut_6_groupCounter = _stageClearVec_reqQueue_fifo_6_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_6_mask = _stageClearVec_reqQueue_fifo_6_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_6_bitMask = _stageClearVec_reqQueue_fifo_6_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_6_data = _stageClearVec_reqQueue_fifo_6_data_out[74:43];
  assign stageClearVec_reqQueue_6_deq_bits_data = stageClearVec_reqQueue_dataOut_6_data;
  assign stageClearVec_reqQueue_6_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_6_bitMask;
  assign stageClearVec_reqQueue_6_deq_bits_mask = stageClearVec_reqQueue_dataOut_6_mask;
  assign stageClearVec_reqQueue_6_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_6_groupCounter;
  assign stageClearVec_reqQueue_6_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_6_ffoByOther;
  assign stageClearVec_reqQueue_6_enq_ready = ~_stageClearVec_reqQueue_fifo_6_full;
  wire        stageClearVec_reqQueue_6_deq_ready;
  wire        stageClearVec_WaitReadQueue_6_deq_valid;
  assign stageClearVec_WaitReadQueue_6_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_6_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_6_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_6_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_6_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_6_groupCounter;
  wire [5:0]  out_6_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_6_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_6_ffoByOther;
  wire        out_6_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_6_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_6 = {stageClearVec_WaitReadQueue_6_enq_bits_groupCounter, stageClearVec_WaitReadQueue_6_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_6 = {stageClearVec_WaitReadQueue_6_enq_bits_data, stageClearVec_WaitReadQueue_6_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_6 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_6, stageClearVec_WaitReadQueue_6_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_6 = {stageClearVec_WaitReadQueue_dataIn_hi_6, stageClearVec_WaitReadQueue_dataIn_lo_6};
  assign stageClearVec_WaitReadQueue_dataOut_6_ffoByOther = _stageClearVec_WaitReadQueue_fifo_6_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_6_groupCounter = _stageClearVec_WaitReadQueue_fifo_6_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_6_mask = _stageClearVec_WaitReadQueue_fifo_6_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_6_bitMask = _stageClearVec_WaitReadQueue_fifo_6_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_6_data = _stageClearVec_WaitReadQueue_fifo_6_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_6_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_6_data;
  wire [31:0] stageClearVec_WaitReadQueue_6_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_6_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_6_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_6_mask;
  assign stageClearVec_WaitReadQueue_6_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_6_groupCounter;
  assign stageClearVec_WaitReadQueue_6_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_6_ffoByOther;
  wire        stageClearVec_WaitReadQueue_6_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_6_full;
  wire        stageClearVec_WaitReadQueue_6_enq_valid;
  wire        stageClearVec_WaitReadQueue_6_deq_ready;
  wire        stageClearVec_readReady_6 = ~needWAR | readChannel_6_ready_0;
  assign stageClearVec_WaitReadQueue_6_enq_valid = stageClearVec_reqQueue_6_deq_valid & stageClearVec_readReady_6;
  assign stageClearVec_reqQueue_6_deq_ready = stageClearVec_WaitReadQueue_6_enq_ready & stageClearVec_readReady_6;
  wire        readChannel_6_valid_0 = stageClearVec_reqQueue_6_deq_valid & needWAR & stageClearVec_WaitReadQueue_6_enq_ready;
  wire [4:0]  readChannel_6_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_6_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_6_bits_offset_0 = stageClearVec_reqQueue_6_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_6 = ~needWAR | readResult_6_valid;
  wire [31:0] stageClearVec_WARData_6 = stageClearVec_WaitReadQueue_6_deq_bits_data & stageClearVec_WaitReadQueue_6_deq_bits_bitMask | readResult_6_bits & ~stageClearVec_WaitReadQueue_6_deq_bits_bitMask;
  wire        out_6_valid_0 = stageClearVec_WaitReadQueue_6_deq_valid & stageClearVec_readResultValid_6;
  assign stageClearVec_WaitReadQueue_6_deq_ready = out_6_ready_0 & stageClearVec_readResultValid_6;
  wire [31:0] out_6_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_6 : stageClearVec_WaitReadQueue_6_deq_bits_data;
  wire [3:0]  out_6_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_6_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_6;
  wire        _stageClearVec_T_18 = in_6_ready_0 & in_6_valid_0;
  wire [2:0]  stageClearVec_counterChange_6 = _stageClearVec_T_18 ? 3'h1 : 3'h7;
  wire        stageClearVec_6 = stageClearVec_counter_6 == 3'h0;
  wire        in_7_ready_0 = stageClearVec_reqQueue_7_enq_ready;
  wire        stageClearVec_reqQueue_7_deq_valid;
  assign stageClearVec_reqQueue_7_deq_valid = ~_stageClearVec_reqQueue_fifo_7_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_7_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_7_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_7_enq_bits_data = stageClearVec_reqQueue_7_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_7_mask;
  wire [31:0] stageClearVec_WaitReadQueue_7_enq_bits_bitMask = stageClearVec_reqQueue_7_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_7_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_7_enq_bits_mask = stageClearVec_reqQueue_7_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_7_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_7_enq_bits_groupCounter = stageClearVec_reqQueue_7_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_7_enq_bits_ffoByOther = stageClearVec_reqQueue_7_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_7 = {stageClearVec_reqQueue_7_enq_bits_groupCounter, stageClearVec_reqQueue_7_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_7 = {stageClearVec_reqQueue_7_enq_bits_data, stageClearVec_reqQueue_7_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_7 = {stageClearVec_reqQueue_dataIn_hi_hi_7, stageClearVec_reqQueue_7_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_7 = {stageClearVec_reqQueue_dataIn_hi_7, stageClearVec_reqQueue_dataIn_lo_7};
  assign stageClearVec_reqQueue_dataOut_7_ffoByOther = _stageClearVec_reqQueue_fifo_7_data_out[0];
  assign stageClearVec_reqQueue_dataOut_7_groupCounter = _stageClearVec_reqQueue_fifo_7_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_7_mask = _stageClearVec_reqQueue_fifo_7_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_7_bitMask = _stageClearVec_reqQueue_fifo_7_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_7_data = _stageClearVec_reqQueue_fifo_7_data_out[74:43];
  assign stageClearVec_reqQueue_7_deq_bits_data = stageClearVec_reqQueue_dataOut_7_data;
  assign stageClearVec_reqQueue_7_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_7_bitMask;
  assign stageClearVec_reqQueue_7_deq_bits_mask = stageClearVec_reqQueue_dataOut_7_mask;
  assign stageClearVec_reqQueue_7_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_7_groupCounter;
  assign stageClearVec_reqQueue_7_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_7_ffoByOther;
  assign stageClearVec_reqQueue_7_enq_ready = ~_stageClearVec_reqQueue_fifo_7_full;
  wire        stageClearVec_reqQueue_7_deq_ready;
  wire        stageClearVec_WaitReadQueue_7_deq_valid;
  assign stageClearVec_WaitReadQueue_7_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_7_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_7_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_7_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_7_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_7_groupCounter;
  wire [5:0]  out_7_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_7_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_7_ffoByOther;
  wire        out_7_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_7_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_7 = {stageClearVec_WaitReadQueue_7_enq_bits_groupCounter, stageClearVec_WaitReadQueue_7_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_7 = {stageClearVec_WaitReadQueue_7_enq_bits_data, stageClearVec_WaitReadQueue_7_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_7 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_7, stageClearVec_WaitReadQueue_7_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_7 = {stageClearVec_WaitReadQueue_dataIn_hi_7, stageClearVec_WaitReadQueue_dataIn_lo_7};
  assign stageClearVec_WaitReadQueue_dataOut_7_ffoByOther = _stageClearVec_WaitReadQueue_fifo_7_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_7_groupCounter = _stageClearVec_WaitReadQueue_fifo_7_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_7_mask = _stageClearVec_WaitReadQueue_fifo_7_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_7_bitMask = _stageClearVec_WaitReadQueue_fifo_7_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_7_data = _stageClearVec_WaitReadQueue_fifo_7_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_7_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_7_data;
  wire [31:0] stageClearVec_WaitReadQueue_7_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_7_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_7_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_7_mask;
  assign stageClearVec_WaitReadQueue_7_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_7_groupCounter;
  assign stageClearVec_WaitReadQueue_7_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_7_ffoByOther;
  wire        stageClearVec_WaitReadQueue_7_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_7_full;
  wire        stageClearVec_WaitReadQueue_7_enq_valid;
  wire        stageClearVec_WaitReadQueue_7_deq_ready;
  wire        stageClearVec_readReady_7 = ~needWAR | readChannel_7_ready_0;
  assign stageClearVec_WaitReadQueue_7_enq_valid = stageClearVec_reqQueue_7_deq_valid & stageClearVec_readReady_7;
  assign stageClearVec_reqQueue_7_deq_ready = stageClearVec_WaitReadQueue_7_enq_ready & stageClearVec_readReady_7;
  wire        readChannel_7_valid_0 = stageClearVec_reqQueue_7_deq_valid & needWAR & stageClearVec_WaitReadQueue_7_enq_ready;
  wire [4:0]  readChannel_7_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_7_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_7_bits_offset_0 = stageClearVec_reqQueue_7_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_7 = ~needWAR | readResult_7_valid;
  wire [31:0] stageClearVec_WARData_7 = stageClearVec_WaitReadQueue_7_deq_bits_data & stageClearVec_WaitReadQueue_7_deq_bits_bitMask | readResult_7_bits & ~stageClearVec_WaitReadQueue_7_deq_bits_bitMask;
  wire        out_7_valid_0 = stageClearVec_WaitReadQueue_7_deq_valid & stageClearVec_readResultValid_7;
  assign stageClearVec_WaitReadQueue_7_deq_ready = out_7_ready_0 & stageClearVec_readResultValid_7;
  wire [31:0] out_7_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_7 : stageClearVec_WaitReadQueue_7_deq_bits_data;
  wire [3:0]  out_7_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_7_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_7;
  wire        _stageClearVec_T_21 = in_7_ready_0 & in_7_valid_0;
  wire [2:0]  stageClearVec_counterChange_7 = _stageClearVec_T_21 ? 3'h1 : 3'h7;
  wire        stageClearVec_7 = stageClearVec_counter_7 == 3'h0;
  wire        in_8_ready_0 = stageClearVec_reqQueue_8_enq_ready;
  wire        stageClearVec_reqQueue_8_deq_valid;
  assign stageClearVec_reqQueue_8_deq_valid = ~_stageClearVec_reqQueue_fifo_8_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_8_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_8_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_8_enq_bits_data = stageClearVec_reqQueue_8_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_8_mask;
  wire [31:0] stageClearVec_WaitReadQueue_8_enq_bits_bitMask = stageClearVec_reqQueue_8_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_8_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_8_enq_bits_mask = stageClearVec_reqQueue_8_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_8_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_8_enq_bits_groupCounter = stageClearVec_reqQueue_8_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_8_enq_bits_ffoByOther = stageClearVec_reqQueue_8_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_8 = {stageClearVec_reqQueue_8_enq_bits_groupCounter, stageClearVec_reqQueue_8_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_8 = {stageClearVec_reqQueue_8_enq_bits_data, stageClearVec_reqQueue_8_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_8 = {stageClearVec_reqQueue_dataIn_hi_hi_8, stageClearVec_reqQueue_8_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_8 = {stageClearVec_reqQueue_dataIn_hi_8, stageClearVec_reqQueue_dataIn_lo_8};
  assign stageClearVec_reqQueue_dataOut_8_ffoByOther = _stageClearVec_reqQueue_fifo_8_data_out[0];
  assign stageClearVec_reqQueue_dataOut_8_groupCounter = _stageClearVec_reqQueue_fifo_8_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_8_mask = _stageClearVec_reqQueue_fifo_8_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_8_bitMask = _stageClearVec_reqQueue_fifo_8_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_8_data = _stageClearVec_reqQueue_fifo_8_data_out[74:43];
  assign stageClearVec_reqQueue_8_deq_bits_data = stageClearVec_reqQueue_dataOut_8_data;
  assign stageClearVec_reqQueue_8_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_8_bitMask;
  assign stageClearVec_reqQueue_8_deq_bits_mask = stageClearVec_reqQueue_dataOut_8_mask;
  assign stageClearVec_reqQueue_8_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_8_groupCounter;
  assign stageClearVec_reqQueue_8_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_8_ffoByOther;
  assign stageClearVec_reqQueue_8_enq_ready = ~_stageClearVec_reqQueue_fifo_8_full;
  wire        stageClearVec_reqQueue_8_deq_ready;
  wire        stageClearVec_WaitReadQueue_8_deq_valid;
  assign stageClearVec_WaitReadQueue_8_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_8_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_8_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_8_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_8_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_8_groupCounter;
  wire [5:0]  out_8_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_8_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_8_ffoByOther;
  wire        out_8_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_8_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_8 = {stageClearVec_WaitReadQueue_8_enq_bits_groupCounter, stageClearVec_WaitReadQueue_8_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_8 = {stageClearVec_WaitReadQueue_8_enq_bits_data, stageClearVec_WaitReadQueue_8_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_8 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_8, stageClearVec_WaitReadQueue_8_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_8 = {stageClearVec_WaitReadQueue_dataIn_hi_8, stageClearVec_WaitReadQueue_dataIn_lo_8};
  assign stageClearVec_WaitReadQueue_dataOut_8_ffoByOther = _stageClearVec_WaitReadQueue_fifo_8_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_8_groupCounter = _stageClearVec_WaitReadQueue_fifo_8_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_8_mask = _stageClearVec_WaitReadQueue_fifo_8_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_8_bitMask = _stageClearVec_WaitReadQueue_fifo_8_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_8_data = _stageClearVec_WaitReadQueue_fifo_8_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_8_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_8_data;
  wire [31:0] stageClearVec_WaitReadQueue_8_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_8_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_8_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_8_mask;
  assign stageClearVec_WaitReadQueue_8_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_8_groupCounter;
  assign stageClearVec_WaitReadQueue_8_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_8_ffoByOther;
  wire        stageClearVec_WaitReadQueue_8_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_8_full;
  wire        stageClearVec_WaitReadQueue_8_enq_valid;
  wire        stageClearVec_WaitReadQueue_8_deq_ready;
  wire        stageClearVec_readReady_8 = ~needWAR | readChannel_8_ready_0;
  assign stageClearVec_WaitReadQueue_8_enq_valid = stageClearVec_reqQueue_8_deq_valid & stageClearVec_readReady_8;
  assign stageClearVec_reqQueue_8_deq_ready = stageClearVec_WaitReadQueue_8_enq_ready & stageClearVec_readReady_8;
  wire        readChannel_8_valid_0 = stageClearVec_reqQueue_8_deq_valid & needWAR & stageClearVec_WaitReadQueue_8_enq_ready;
  wire [4:0]  readChannel_8_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_8_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_8_bits_offset_0 = stageClearVec_reqQueue_8_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_8 = ~needWAR | readResult_8_valid;
  wire [31:0] stageClearVec_WARData_8 = stageClearVec_WaitReadQueue_8_deq_bits_data & stageClearVec_WaitReadQueue_8_deq_bits_bitMask | readResult_8_bits & ~stageClearVec_WaitReadQueue_8_deq_bits_bitMask;
  wire        out_8_valid_0 = stageClearVec_WaitReadQueue_8_deq_valid & stageClearVec_readResultValid_8;
  assign stageClearVec_WaitReadQueue_8_deq_ready = out_8_ready_0 & stageClearVec_readResultValid_8;
  wire [31:0] out_8_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_8 : stageClearVec_WaitReadQueue_8_deq_bits_data;
  wire [3:0]  out_8_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_8_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_8;
  wire        _stageClearVec_T_24 = in_8_ready_0 & in_8_valid_0;
  wire [2:0]  stageClearVec_counterChange_8 = _stageClearVec_T_24 ? 3'h1 : 3'h7;
  wire        stageClearVec_8 = stageClearVec_counter_8 == 3'h0;
  wire        in_9_ready_0 = stageClearVec_reqQueue_9_enq_ready;
  wire        stageClearVec_reqQueue_9_deq_valid;
  assign stageClearVec_reqQueue_9_deq_valid = ~_stageClearVec_reqQueue_fifo_9_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_9_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_9_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_9_enq_bits_data = stageClearVec_reqQueue_9_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_9_mask;
  wire [31:0] stageClearVec_WaitReadQueue_9_enq_bits_bitMask = stageClearVec_reqQueue_9_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_9_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_9_enq_bits_mask = stageClearVec_reqQueue_9_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_9_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_9_enq_bits_groupCounter = stageClearVec_reqQueue_9_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_9_enq_bits_ffoByOther = stageClearVec_reqQueue_9_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_9 = {stageClearVec_reqQueue_9_enq_bits_groupCounter, stageClearVec_reqQueue_9_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_9 = {stageClearVec_reqQueue_9_enq_bits_data, stageClearVec_reqQueue_9_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_9 = {stageClearVec_reqQueue_dataIn_hi_hi_9, stageClearVec_reqQueue_9_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_9 = {stageClearVec_reqQueue_dataIn_hi_9, stageClearVec_reqQueue_dataIn_lo_9};
  assign stageClearVec_reqQueue_dataOut_9_ffoByOther = _stageClearVec_reqQueue_fifo_9_data_out[0];
  assign stageClearVec_reqQueue_dataOut_9_groupCounter = _stageClearVec_reqQueue_fifo_9_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_9_mask = _stageClearVec_reqQueue_fifo_9_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_9_bitMask = _stageClearVec_reqQueue_fifo_9_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_9_data = _stageClearVec_reqQueue_fifo_9_data_out[74:43];
  assign stageClearVec_reqQueue_9_deq_bits_data = stageClearVec_reqQueue_dataOut_9_data;
  assign stageClearVec_reqQueue_9_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_9_bitMask;
  assign stageClearVec_reqQueue_9_deq_bits_mask = stageClearVec_reqQueue_dataOut_9_mask;
  assign stageClearVec_reqQueue_9_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_9_groupCounter;
  assign stageClearVec_reqQueue_9_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_9_ffoByOther;
  assign stageClearVec_reqQueue_9_enq_ready = ~_stageClearVec_reqQueue_fifo_9_full;
  wire        stageClearVec_reqQueue_9_deq_ready;
  wire        stageClearVec_WaitReadQueue_9_deq_valid;
  assign stageClearVec_WaitReadQueue_9_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_9_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_9_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_9_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_9_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_9_groupCounter;
  wire [5:0]  out_9_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_9_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_9_ffoByOther;
  wire        out_9_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_9_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_9 = {stageClearVec_WaitReadQueue_9_enq_bits_groupCounter, stageClearVec_WaitReadQueue_9_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_9 = {stageClearVec_WaitReadQueue_9_enq_bits_data, stageClearVec_WaitReadQueue_9_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_9 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_9, stageClearVec_WaitReadQueue_9_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_9 = {stageClearVec_WaitReadQueue_dataIn_hi_9, stageClearVec_WaitReadQueue_dataIn_lo_9};
  assign stageClearVec_WaitReadQueue_dataOut_9_ffoByOther = _stageClearVec_WaitReadQueue_fifo_9_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_9_groupCounter = _stageClearVec_WaitReadQueue_fifo_9_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_9_mask = _stageClearVec_WaitReadQueue_fifo_9_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_9_bitMask = _stageClearVec_WaitReadQueue_fifo_9_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_9_data = _stageClearVec_WaitReadQueue_fifo_9_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_9_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_9_data;
  wire [31:0] stageClearVec_WaitReadQueue_9_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_9_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_9_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_9_mask;
  assign stageClearVec_WaitReadQueue_9_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_9_groupCounter;
  assign stageClearVec_WaitReadQueue_9_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_9_ffoByOther;
  wire        stageClearVec_WaitReadQueue_9_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_9_full;
  wire        stageClearVec_WaitReadQueue_9_enq_valid;
  wire        stageClearVec_WaitReadQueue_9_deq_ready;
  wire        stageClearVec_readReady_9 = ~needWAR | readChannel_9_ready_0;
  assign stageClearVec_WaitReadQueue_9_enq_valid = stageClearVec_reqQueue_9_deq_valid & stageClearVec_readReady_9;
  assign stageClearVec_reqQueue_9_deq_ready = stageClearVec_WaitReadQueue_9_enq_ready & stageClearVec_readReady_9;
  wire        readChannel_9_valid_0 = stageClearVec_reqQueue_9_deq_valid & needWAR & stageClearVec_WaitReadQueue_9_enq_ready;
  wire [4:0]  readChannel_9_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_9_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_9_bits_offset_0 = stageClearVec_reqQueue_9_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_9 = ~needWAR | readResult_9_valid;
  wire [31:0] stageClearVec_WARData_9 = stageClearVec_WaitReadQueue_9_deq_bits_data & stageClearVec_WaitReadQueue_9_deq_bits_bitMask | readResult_9_bits & ~stageClearVec_WaitReadQueue_9_deq_bits_bitMask;
  wire        out_9_valid_0 = stageClearVec_WaitReadQueue_9_deq_valid & stageClearVec_readResultValid_9;
  assign stageClearVec_WaitReadQueue_9_deq_ready = out_9_ready_0 & stageClearVec_readResultValid_9;
  wire [31:0] out_9_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_9 : stageClearVec_WaitReadQueue_9_deq_bits_data;
  wire [3:0]  out_9_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_9_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_9;
  wire        _stageClearVec_T_27 = in_9_ready_0 & in_9_valid_0;
  wire [2:0]  stageClearVec_counterChange_9 = _stageClearVec_T_27 ? 3'h1 : 3'h7;
  wire        stageClearVec_9 = stageClearVec_counter_9 == 3'h0;
  wire        in_10_ready_0 = stageClearVec_reqQueue_10_enq_ready;
  wire        stageClearVec_reqQueue_10_deq_valid;
  assign stageClearVec_reqQueue_10_deq_valid = ~_stageClearVec_reqQueue_fifo_10_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_10_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_10_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_10_enq_bits_data = stageClearVec_reqQueue_10_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_10_mask;
  wire [31:0] stageClearVec_WaitReadQueue_10_enq_bits_bitMask = stageClearVec_reqQueue_10_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_10_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_10_enq_bits_mask = stageClearVec_reqQueue_10_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_10_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_10_enq_bits_groupCounter = stageClearVec_reqQueue_10_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_10_enq_bits_ffoByOther = stageClearVec_reqQueue_10_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_10 = {stageClearVec_reqQueue_10_enq_bits_groupCounter, stageClearVec_reqQueue_10_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_10 = {stageClearVec_reqQueue_10_enq_bits_data, stageClearVec_reqQueue_10_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_10 = {stageClearVec_reqQueue_dataIn_hi_hi_10, stageClearVec_reqQueue_10_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_10 = {stageClearVec_reqQueue_dataIn_hi_10, stageClearVec_reqQueue_dataIn_lo_10};
  assign stageClearVec_reqQueue_dataOut_10_ffoByOther = _stageClearVec_reqQueue_fifo_10_data_out[0];
  assign stageClearVec_reqQueue_dataOut_10_groupCounter = _stageClearVec_reqQueue_fifo_10_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_10_mask = _stageClearVec_reqQueue_fifo_10_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_10_bitMask = _stageClearVec_reqQueue_fifo_10_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_10_data = _stageClearVec_reqQueue_fifo_10_data_out[74:43];
  assign stageClearVec_reqQueue_10_deq_bits_data = stageClearVec_reqQueue_dataOut_10_data;
  assign stageClearVec_reqQueue_10_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_10_bitMask;
  assign stageClearVec_reqQueue_10_deq_bits_mask = stageClearVec_reqQueue_dataOut_10_mask;
  assign stageClearVec_reqQueue_10_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_10_groupCounter;
  assign stageClearVec_reqQueue_10_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_10_ffoByOther;
  assign stageClearVec_reqQueue_10_enq_ready = ~_stageClearVec_reqQueue_fifo_10_full;
  wire        stageClearVec_reqQueue_10_deq_ready;
  wire        stageClearVec_WaitReadQueue_10_deq_valid;
  assign stageClearVec_WaitReadQueue_10_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_10_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_10_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_10_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_10_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_10_groupCounter;
  wire [5:0]  out_10_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_10_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_10_ffoByOther;
  wire        out_10_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_10_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_10 = {stageClearVec_WaitReadQueue_10_enq_bits_groupCounter, stageClearVec_WaitReadQueue_10_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_10 = {stageClearVec_WaitReadQueue_10_enq_bits_data, stageClearVec_WaitReadQueue_10_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_10 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_10, stageClearVec_WaitReadQueue_10_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_10 = {stageClearVec_WaitReadQueue_dataIn_hi_10, stageClearVec_WaitReadQueue_dataIn_lo_10};
  assign stageClearVec_WaitReadQueue_dataOut_10_ffoByOther = _stageClearVec_WaitReadQueue_fifo_10_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_10_groupCounter = _stageClearVec_WaitReadQueue_fifo_10_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_10_mask = _stageClearVec_WaitReadQueue_fifo_10_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_10_bitMask = _stageClearVec_WaitReadQueue_fifo_10_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_10_data = _stageClearVec_WaitReadQueue_fifo_10_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_10_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_10_data;
  wire [31:0] stageClearVec_WaitReadQueue_10_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_10_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_10_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_10_mask;
  assign stageClearVec_WaitReadQueue_10_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_10_groupCounter;
  assign stageClearVec_WaitReadQueue_10_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_10_ffoByOther;
  wire        stageClearVec_WaitReadQueue_10_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_10_full;
  wire        stageClearVec_WaitReadQueue_10_enq_valid;
  wire        stageClearVec_WaitReadQueue_10_deq_ready;
  wire        stageClearVec_readReady_10 = ~needWAR | readChannel_10_ready_0;
  assign stageClearVec_WaitReadQueue_10_enq_valid = stageClearVec_reqQueue_10_deq_valid & stageClearVec_readReady_10;
  assign stageClearVec_reqQueue_10_deq_ready = stageClearVec_WaitReadQueue_10_enq_ready & stageClearVec_readReady_10;
  wire        readChannel_10_valid_0 = stageClearVec_reqQueue_10_deq_valid & needWAR & stageClearVec_WaitReadQueue_10_enq_ready;
  wire [4:0]  readChannel_10_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_10_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_10_bits_offset_0 = stageClearVec_reqQueue_10_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_10 = ~needWAR | readResult_10_valid;
  wire [31:0] stageClearVec_WARData_10 = stageClearVec_WaitReadQueue_10_deq_bits_data & stageClearVec_WaitReadQueue_10_deq_bits_bitMask | readResult_10_bits & ~stageClearVec_WaitReadQueue_10_deq_bits_bitMask;
  wire        out_10_valid_0 = stageClearVec_WaitReadQueue_10_deq_valid & stageClearVec_readResultValid_10;
  assign stageClearVec_WaitReadQueue_10_deq_ready = out_10_ready_0 & stageClearVec_readResultValid_10;
  wire [31:0] out_10_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_10 : stageClearVec_WaitReadQueue_10_deq_bits_data;
  wire [3:0]  out_10_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_10_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_10;
  wire        _stageClearVec_T_30 = in_10_ready_0 & in_10_valid_0;
  wire [2:0]  stageClearVec_counterChange_10 = _stageClearVec_T_30 ? 3'h1 : 3'h7;
  wire        stageClearVec_10 = stageClearVec_counter_10 == 3'h0;
  wire        in_11_ready_0 = stageClearVec_reqQueue_11_enq_ready;
  wire        stageClearVec_reqQueue_11_deq_valid;
  assign stageClearVec_reqQueue_11_deq_valid = ~_stageClearVec_reqQueue_fifo_11_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_11_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_11_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_11_enq_bits_data = stageClearVec_reqQueue_11_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_11_mask;
  wire [31:0] stageClearVec_WaitReadQueue_11_enq_bits_bitMask = stageClearVec_reqQueue_11_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_11_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_11_enq_bits_mask = stageClearVec_reqQueue_11_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_11_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_11_enq_bits_groupCounter = stageClearVec_reqQueue_11_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_11_enq_bits_ffoByOther = stageClearVec_reqQueue_11_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_11 = {stageClearVec_reqQueue_11_enq_bits_groupCounter, stageClearVec_reqQueue_11_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_11 = {stageClearVec_reqQueue_11_enq_bits_data, stageClearVec_reqQueue_11_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_11 = {stageClearVec_reqQueue_dataIn_hi_hi_11, stageClearVec_reqQueue_11_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_11 = {stageClearVec_reqQueue_dataIn_hi_11, stageClearVec_reqQueue_dataIn_lo_11};
  assign stageClearVec_reqQueue_dataOut_11_ffoByOther = _stageClearVec_reqQueue_fifo_11_data_out[0];
  assign stageClearVec_reqQueue_dataOut_11_groupCounter = _stageClearVec_reqQueue_fifo_11_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_11_mask = _stageClearVec_reqQueue_fifo_11_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_11_bitMask = _stageClearVec_reqQueue_fifo_11_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_11_data = _stageClearVec_reqQueue_fifo_11_data_out[74:43];
  assign stageClearVec_reqQueue_11_deq_bits_data = stageClearVec_reqQueue_dataOut_11_data;
  assign stageClearVec_reqQueue_11_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_11_bitMask;
  assign stageClearVec_reqQueue_11_deq_bits_mask = stageClearVec_reqQueue_dataOut_11_mask;
  assign stageClearVec_reqQueue_11_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_11_groupCounter;
  assign stageClearVec_reqQueue_11_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_11_ffoByOther;
  assign stageClearVec_reqQueue_11_enq_ready = ~_stageClearVec_reqQueue_fifo_11_full;
  wire        stageClearVec_reqQueue_11_deq_ready;
  wire        stageClearVec_WaitReadQueue_11_deq_valid;
  assign stageClearVec_WaitReadQueue_11_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_11_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_11_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_11_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_11_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_11_groupCounter;
  wire [5:0]  out_11_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_11_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_11_ffoByOther;
  wire        out_11_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_11_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_11 = {stageClearVec_WaitReadQueue_11_enq_bits_groupCounter, stageClearVec_WaitReadQueue_11_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_11 = {stageClearVec_WaitReadQueue_11_enq_bits_data, stageClearVec_WaitReadQueue_11_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_11 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_11, stageClearVec_WaitReadQueue_11_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_11 = {stageClearVec_WaitReadQueue_dataIn_hi_11, stageClearVec_WaitReadQueue_dataIn_lo_11};
  assign stageClearVec_WaitReadQueue_dataOut_11_ffoByOther = _stageClearVec_WaitReadQueue_fifo_11_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_11_groupCounter = _stageClearVec_WaitReadQueue_fifo_11_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_11_mask = _stageClearVec_WaitReadQueue_fifo_11_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_11_bitMask = _stageClearVec_WaitReadQueue_fifo_11_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_11_data = _stageClearVec_WaitReadQueue_fifo_11_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_11_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_11_data;
  wire [31:0] stageClearVec_WaitReadQueue_11_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_11_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_11_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_11_mask;
  assign stageClearVec_WaitReadQueue_11_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_11_groupCounter;
  assign stageClearVec_WaitReadQueue_11_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_11_ffoByOther;
  wire        stageClearVec_WaitReadQueue_11_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_11_full;
  wire        stageClearVec_WaitReadQueue_11_enq_valid;
  wire        stageClearVec_WaitReadQueue_11_deq_ready;
  wire        stageClearVec_readReady_11 = ~needWAR | readChannel_11_ready_0;
  assign stageClearVec_WaitReadQueue_11_enq_valid = stageClearVec_reqQueue_11_deq_valid & stageClearVec_readReady_11;
  assign stageClearVec_reqQueue_11_deq_ready = stageClearVec_WaitReadQueue_11_enq_ready & stageClearVec_readReady_11;
  wire        readChannel_11_valid_0 = stageClearVec_reqQueue_11_deq_valid & needWAR & stageClearVec_WaitReadQueue_11_enq_ready;
  wire [4:0]  readChannel_11_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_11_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_11_bits_offset_0 = stageClearVec_reqQueue_11_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_11 = ~needWAR | readResult_11_valid;
  wire [31:0] stageClearVec_WARData_11 = stageClearVec_WaitReadQueue_11_deq_bits_data & stageClearVec_WaitReadQueue_11_deq_bits_bitMask | readResult_11_bits & ~stageClearVec_WaitReadQueue_11_deq_bits_bitMask;
  wire        out_11_valid_0 = stageClearVec_WaitReadQueue_11_deq_valid & stageClearVec_readResultValid_11;
  assign stageClearVec_WaitReadQueue_11_deq_ready = out_11_ready_0 & stageClearVec_readResultValid_11;
  wire [31:0] out_11_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_11 : stageClearVec_WaitReadQueue_11_deq_bits_data;
  wire [3:0]  out_11_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_11_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_11;
  wire        _stageClearVec_T_33 = in_11_ready_0 & in_11_valid_0;
  wire [2:0]  stageClearVec_counterChange_11 = _stageClearVec_T_33 ? 3'h1 : 3'h7;
  wire        stageClearVec_11 = stageClearVec_counter_11 == 3'h0;
  wire        in_12_ready_0 = stageClearVec_reqQueue_12_enq_ready;
  wire        stageClearVec_reqQueue_12_deq_valid;
  assign stageClearVec_reqQueue_12_deq_valid = ~_stageClearVec_reqQueue_fifo_12_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_12_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_12_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_12_enq_bits_data = stageClearVec_reqQueue_12_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_12_mask;
  wire [31:0] stageClearVec_WaitReadQueue_12_enq_bits_bitMask = stageClearVec_reqQueue_12_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_12_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_12_enq_bits_mask = stageClearVec_reqQueue_12_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_12_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_12_enq_bits_groupCounter = stageClearVec_reqQueue_12_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_12_enq_bits_ffoByOther = stageClearVec_reqQueue_12_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_12 = {stageClearVec_reqQueue_12_enq_bits_groupCounter, stageClearVec_reqQueue_12_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_12 = {stageClearVec_reqQueue_12_enq_bits_data, stageClearVec_reqQueue_12_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_12 = {stageClearVec_reqQueue_dataIn_hi_hi_12, stageClearVec_reqQueue_12_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_12 = {stageClearVec_reqQueue_dataIn_hi_12, stageClearVec_reqQueue_dataIn_lo_12};
  assign stageClearVec_reqQueue_dataOut_12_ffoByOther = _stageClearVec_reqQueue_fifo_12_data_out[0];
  assign stageClearVec_reqQueue_dataOut_12_groupCounter = _stageClearVec_reqQueue_fifo_12_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_12_mask = _stageClearVec_reqQueue_fifo_12_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_12_bitMask = _stageClearVec_reqQueue_fifo_12_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_12_data = _stageClearVec_reqQueue_fifo_12_data_out[74:43];
  assign stageClearVec_reqQueue_12_deq_bits_data = stageClearVec_reqQueue_dataOut_12_data;
  assign stageClearVec_reqQueue_12_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_12_bitMask;
  assign stageClearVec_reqQueue_12_deq_bits_mask = stageClearVec_reqQueue_dataOut_12_mask;
  assign stageClearVec_reqQueue_12_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_12_groupCounter;
  assign stageClearVec_reqQueue_12_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_12_ffoByOther;
  assign stageClearVec_reqQueue_12_enq_ready = ~_stageClearVec_reqQueue_fifo_12_full;
  wire        stageClearVec_reqQueue_12_deq_ready;
  wire        stageClearVec_WaitReadQueue_12_deq_valid;
  assign stageClearVec_WaitReadQueue_12_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_12_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_12_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_12_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_12_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_12_groupCounter;
  wire [5:0]  out_12_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_12_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_12_ffoByOther;
  wire        out_12_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_12_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_12 = {stageClearVec_WaitReadQueue_12_enq_bits_groupCounter, stageClearVec_WaitReadQueue_12_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_12 = {stageClearVec_WaitReadQueue_12_enq_bits_data, stageClearVec_WaitReadQueue_12_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_12 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_12, stageClearVec_WaitReadQueue_12_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_12 = {stageClearVec_WaitReadQueue_dataIn_hi_12, stageClearVec_WaitReadQueue_dataIn_lo_12};
  assign stageClearVec_WaitReadQueue_dataOut_12_ffoByOther = _stageClearVec_WaitReadQueue_fifo_12_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_12_groupCounter = _stageClearVec_WaitReadQueue_fifo_12_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_12_mask = _stageClearVec_WaitReadQueue_fifo_12_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_12_bitMask = _stageClearVec_WaitReadQueue_fifo_12_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_12_data = _stageClearVec_WaitReadQueue_fifo_12_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_12_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_12_data;
  wire [31:0] stageClearVec_WaitReadQueue_12_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_12_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_12_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_12_mask;
  assign stageClearVec_WaitReadQueue_12_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_12_groupCounter;
  assign stageClearVec_WaitReadQueue_12_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_12_ffoByOther;
  wire        stageClearVec_WaitReadQueue_12_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_12_full;
  wire        stageClearVec_WaitReadQueue_12_enq_valid;
  wire        stageClearVec_WaitReadQueue_12_deq_ready;
  wire        stageClearVec_readReady_12 = ~needWAR | readChannel_12_ready_0;
  assign stageClearVec_WaitReadQueue_12_enq_valid = stageClearVec_reqQueue_12_deq_valid & stageClearVec_readReady_12;
  assign stageClearVec_reqQueue_12_deq_ready = stageClearVec_WaitReadQueue_12_enq_ready & stageClearVec_readReady_12;
  wire        readChannel_12_valid_0 = stageClearVec_reqQueue_12_deq_valid & needWAR & stageClearVec_WaitReadQueue_12_enq_ready;
  wire [4:0]  readChannel_12_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_12_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_12_bits_offset_0 = stageClearVec_reqQueue_12_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_12 = ~needWAR | readResult_12_valid;
  wire [31:0] stageClearVec_WARData_12 = stageClearVec_WaitReadQueue_12_deq_bits_data & stageClearVec_WaitReadQueue_12_deq_bits_bitMask | readResult_12_bits & ~stageClearVec_WaitReadQueue_12_deq_bits_bitMask;
  wire        out_12_valid_0 = stageClearVec_WaitReadQueue_12_deq_valid & stageClearVec_readResultValid_12;
  assign stageClearVec_WaitReadQueue_12_deq_ready = out_12_ready_0 & stageClearVec_readResultValid_12;
  wire [31:0] out_12_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_12 : stageClearVec_WaitReadQueue_12_deq_bits_data;
  wire [3:0]  out_12_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_12_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_12;
  wire        _stageClearVec_T_36 = in_12_ready_0 & in_12_valid_0;
  wire [2:0]  stageClearVec_counterChange_12 = _stageClearVec_T_36 ? 3'h1 : 3'h7;
  wire        stageClearVec_12 = stageClearVec_counter_12 == 3'h0;
  wire        in_13_ready_0 = stageClearVec_reqQueue_13_enq_ready;
  wire        stageClearVec_reqQueue_13_deq_valid;
  assign stageClearVec_reqQueue_13_deq_valid = ~_stageClearVec_reqQueue_fifo_13_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_13_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_13_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_13_enq_bits_data = stageClearVec_reqQueue_13_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_13_mask;
  wire [31:0] stageClearVec_WaitReadQueue_13_enq_bits_bitMask = stageClearVec_reqQueue_13_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_13_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_13_enq_bits_mask = stageClearVec_reqQueue_13_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_13_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_13_enq_bits_groupCounter = stageClearVec_reqQueue_13_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_13_enq_bits_ffoByOther = stageClearVec_reqQueue_13_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_13 = {stageClearVec_reqQueue_13_enq_bits_groupCounter, stageClearVec_reqQueue_13_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_13 = {stageClearVec_reqQueue_13_enq_bits_data, stageClearVec_reqQueue_13_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_13 = {stageClearVec_reqQueue_dataIn_hi_hi_13, stageClearVec_reqQueue_13_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_13 = {stageClearVec_reqQueue_dataIn_hi_13, stageClearVec_reqQueue_dataIn_lo_13};
  assign stageClearVec_reqQueue_dataOut_13_ffoByOther = _stageClearVec_reqQueue_fifo_13_data_out[0];
  assign stageClearVec_reqQueue_dataOut_13_groupCounter = _stageClearVec_reqQueue_fifo_13_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_13_mask = _stageClearVec_reqQueue_fifo_13_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_13_bitMask = _stageClearVec_reqQueue_fifo_13_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_13_data = _stageClearVec_reqQueue_fifo_13_data_out[74:43];
  assign stageClearVec_reqQueue_13_deq_bits_data = stageClearVec_reqQueue_dataOut_13_data;
  assign stageClearVec_reqQueue_13_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_13_bitMask;
  assign stageClearVec_reqQueue_13_deq_bits_mask = stageClearVec_reqQueue_dataOut_13_mask;
  assign stageClearVec_reqQueue_13_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_13_groupCounter;
  assign stageClearVec_reqQueue_13_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_13_ffoByOther;
  assign stageClearVec_reqQueue_13_enq_ready = ~_stageClearVec_reqQueue_fifo_13_full;
  wire        stageClearVec_reqQueue_13_deq_ready;
  wire        stageClearVec_WaitReadQueue_13_deq_valid;
  assign stageClearVec_WaitReadQueue_13_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_13_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_13_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_13_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_13_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_13_groupCounter;
  wire [5:0]  out_13_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_13_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_13_ffoByOther;
  wire        out_13_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_13_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_13 = {stageClearVec_WaitReadQueue_13_enq_bits_groupCounter, stageClearVec_WaitReadQueue_13_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_13 = {stageClearVec_WaitReadQueue_13_enq_bits_data, stageClearVec_WaitReadQueue_13_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_13 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_13, stageClearVec_WaitReadQueue_13_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_13 = {stageClearVec_WaitReadQueue_dataIn_hi_13, stageClearVec_WaitReadQueue_dataIn_lo_13};
  assign stageClearVec_WaitReadQueue_dataOut_13_ffoByOther = _stageClearVec_WaitReadQueue_fifo_13_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_13_groupCounter = _stageClearVec_WaitReadQueue_fifo_13_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_13_mask = _stageClearVec_WaitReadQueue_fifo_13_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_13_bitMask = _stageClearVec_WaitReadQueue_fifo_13_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_13_data = _stageClearVec_WaitReadQueue_fifo_13_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_13_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_13_data;
  wire [31:0] stageClearVec_WaitReadQueue_13_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_13_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_13_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_13_mask;
  assign stageClearVec_WaitReadQueue_13_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_13_groupCounter;
  assign stageClearVec_WaitReadQueue_13_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_13_ffoByOther;
  wire        stageClearVec_WaitReadQueue_13_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_13_full;
  wire        stageClearVec_WaitReadQueue_13_enq_valid;
  wire        stageClearVec_WaitReadQueue_13_deq_ready;
  wire        stageClearVec_readReady_13 = ~needWAR | readChannel_13_ready_0;
  assign stageClearVec_WaitReadQueue_13_enq_valid = stageClearVec_reqQueue_13_deq_valid & stageClearVec_readReady_13;
  assign stageClearVec_reqQueue_13_deq_ready = stageClearVec_WaitReadQueue_13_enq_ready & stageClearVec_readReady_13;
  wire        readChannel_13_valid_0 = stageClearVec_reqQueue_13_deq_valid & needWAR & stageClearVec_WaitReadQueue_13_enq_ready;
  wire [4:0]  readChannel_13_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_13_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_13_bits_offset_0 = stageClearVec_reqQueue_13_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_13 = ~needWAR | readResult_13_valid;
  wire [31:0] stageClearVec_WARData_13 = stageClearVec_WaitReadQueue_13_deq_bits_data & stageClearVec_WaitReadQueue_13_deq_bits_bitMask | readResult_13_bits & ~stageClearVec_WaitReadQueue_13_deq_bits_bitMask;
  wire        out_13_valid_0 = stageClearVec_WaitReadQueue_13_deq_valid & stageClearVec_readResultValid_13;
  assign stageClearVec_WaitReadQueue_13_deq_ready = out_13_ready_0 & stageClearVec_readResultValid_13;
  wire [31:0] out_13_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_13 : stageClearVec_WaitReadQueue_13_deq_bits_data;
  wire [3:0]  out_13_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_13_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_13;
  wire        _stageClearVec_T_39 = in_13_ready_0 & in_13_valid_0;
  wire [2:0]  stageClearVec_counterChange_13 = _stageClearVec_T_39 ? 3'h1 : 3'h7;
  wire        stageClearVec_13 = stageClearVec_counter_13 == 3'h0;
  wire        in_14_ready_0 = stageClearVec_reqQueue_14_enq_ready;
  wire        stageClearVec_reqQueue_14_deq_valid;
  assign stageClearVec_reqQueue_14_deq_valid = ~_stageClearVec_reqQueue_fifo_14_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_14_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_14_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_14_enq_bits_data = stageClearVec_reqQueue_14_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_14_mask;
  wire [31:0] stageClearVec_WaitReadQueue_14_enq_bits_bitMask = stageClearVec_reqQueue_14_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_14_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_14_enq_bits_mask = stageClearVec_reqQueue_14_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_14_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_14_enq_bits_groupCounter = stageClearVec_reqQueue_14_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_14_enq_bits_ffoByOther = stageClearVec_reqQueue_14_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_14 = {stageClearVec_reqQueue_14_enq_bits_groupCounter, stageClearVec_reqQueue_14_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_14 = {stageClearVec_reqQueue_14_enq_bits_data, stageClearVec_reqQueue_14_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_14 = {stageClearVec_reqQueue_dataIn_hi_hi_14, stageClearVec_reqQueue_14_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_14 = {stageClearVec_reqQueue_dataIn_hi_14, stageClearVec_reqQueue_dataIn_lo_14};
  assign stageClearVec_reqQueue_dataOut_14_ffoByOther = _stageClearVec_reqQueue_fifo_14_data_out[0];
  assign stageClearVec_reqQueue_dataOut_14_groupCounter = _stageClearVec_reqQueue_fifo_14_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_14_mask = _stageClearVec_reqQueue_fifo_14_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_14_bitMask = _stageClearVec_reqQueue_fifo_14_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_14_data = _stageClearVec_reqQueue_fifo_14_data_out[74:43];
  assign stageClearVec_reqQueue_14_deq_bits_data = stageClearVec_reqQueue_dataOut_14_data;
  assign stageClearVec_reqQueue_14_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_14_bitMask;
  assign stageClearVec_reqQueue_14_deq_bits_mask = stageClearVec_reqQueue_dataOut_14_mask;
  assign stageClearVec_reqQueue_14_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_14_groupCounter;
  assign stageClearVec_reqQueue_14_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_14_ffoByOther;
  assign stageClearVec_reqQueue_14_enq_ready = ~_stageClearVec_reqQueue_fifo_14_full;
  wire        stageClearVec_reqQueue_14_deq_ready;
  wire        stageClearVec_WaitReadQueue_14_deq_valid;
  assign stageClearVec_WaitReadQueue_14_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_14_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_14_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_14_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_14_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_14_groupCounter;
  wire [5:0]  out_14_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_14_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_14_ffoByOther;
  wire        out_14_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_14_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_14 = {stageClearVec_WaitReadQueue_14_enq_bits_groupCounter, stageClearVec_WaitReadQueue_14_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_14 = {stageClearVec_WaitReadQueue_14_enq_bits_data, stageClearVec_WaitReadQueue_14_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_14 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_14, stageClearVec_WaitReadQueue_14_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_14 = {stageClearVec_WaitReadQueue_dataIn_hi_14, stageClearVec_WaitReadQueue_dataIn_lo_14};
  assign stageClearVec_WaitReadQueue_dataOut_14_ffoByOther = _stageClearVec_WaitReadQueue_fifo_14_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_14_groupCounter = _stageClearVec_WaitReadQueue_fifo_14_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_14_mask = _stageClearVec_WaitReadQueue_fifo_14_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_14_bitMask = _stageClearVec_WaitReadQueue_fifo_14_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_14_data = _stageClearVec_WaitReadQueue_fifo_14_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_14_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_14_data;
  wire [31:0] stageClearVec_WaitReadQueue_14_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_14_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_14_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_14_mask;
  assign stageClearVec_WaitReadQueue_14_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_14_groupCounter;
  assign stageClearVec_WaitReadQueue_14_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_14_ffoByOther;
  wire        stageClearVec_WaitReadQueue_14_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_14_full;
  wire        stageClearVec_WaitReadQueue_14_enq_valid;
  wire        stageClearVec_WaitReadQueue_14_deq_ready;
  wire        stageClearVec_readReady_14 = ~needWAR | readChannel_14_ready_0;
  assign stageClearVec_WaitReadQueue_14_enq_valid = stageClearVec_reqQueue_14_deq_valid & stageClearVec_readReady_14;
  assign stageClearVec_reqQueue_14_deq_ready = stageClearVec_WaitReadQueue_14_enq_ready & stageClearVec_readReady_14;
  wire        readChannel_14_valid_0 = stageClearVec_reqQueue_14_deq_valid & needWAR & stageClearVec_WaitReadQueue_14_enq_ready;
  wire [4:0]  readChannel_14_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_14_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_14_bits_offset_0 = stageClearVec_reqQueue_14_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_14 = ~needWAR | readResult_14_valid;
  wire [31:0] stageClearVec_WARData_14 = stageClearVec_WaitReadQueue_14_deq_bits_data & stageClearVec_WaitReadQueue_14_deq_bits_bitMask | readResult_14_bits & ~stageClearVec_WaitReadQueue_14_deq_bits_bitMask;
  wire        out_14_valid_0 = stageClearVec_WaitReadQueue_14_deq_valid & stageClearVec_readResultValid_14;
  assign stageClearVec_WaitReadQueue_14_deq_ready = out_14_ready_0 & stageClearVec_readResultValid_14;
  wire [31:0] out_14_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_14 : stageClearVec_WaitReadQueue_14_deq_bits_data;
  wire [3:0]  out_14_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_14_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_14;
  wire        _stageClearVec_T_42 = in_14_ready_0 & in_14_valid_0;
  wire [2:0]  stageClearVec_counterChange_14 = _stageClearVec_T_42 ? 3'h1 : 3'h7;
  wire        stageClearVec_14 = stageClearVec_counter_14 == 3'h0;
  wire        in_15_ready_0 = stageClearVec_reqQueue_15_enq_ready;
  wire        stageClearVec_reqQueue_15_deq_valid;
  assign stageClearVec_reqQueue_15_deq_valid = ~_stageClearVec_reqQueue_fifo_15_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_15_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_15_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_15_enq_bits_data = stageClearVec_reqQueue_15_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_15_mask;
  wire [31:0] stageClearVec_WaitReadQueue_15_enq_bits_bitMask = stageClearVec_reqQueue_15_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_15_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_15_enq_bits_mask = stageClearVec_reqQueue_15_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_15_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_15_enq_bits_groupCounter = stageClearVec_reqQueue_15_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_15_enq_bits_ffoByOther = stageClearVec_reqQueue_15_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_15 = {stageClearVec_reqQueue_15_enq_bits_groupCounter, stageClearVec_reqQueue_15_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_15 = {stageClearVec_reqQueue_15_enq_bits_data, stageClearVec_reqQueue_15_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_15 = {stageClearVec_reqQueue_dataIn_hi_hi_15, stageClearVec_reqQueue_15_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_15 = {stageClearVec_reqQueue_dataIn_hi_15, stageClearVec_reqQueue_dataIn_lo_15};
  assign stageClearVec_reqQueue_dataOut_15_ffoByOther = _stageClearVec_reqQueue_fifo_15_data_out[0];
  assign stageClearVec_reqQueue_dataOut_15_groupCounter = _stageClearVec_reqQueue_fifo_15_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_15_mask = _stageClearVec_reqQueue_fifo_15_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_15_bitMask = _stageClearVec_reqQueue_fifo_15_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_15_data = _stageClearVec_reqQueue_fifo_15_data_out[74:43];
  assign stageClearVec_reqQueue_15_deq_bits_data = stageClearVec_reqQueue_dataOut_15_data;
  assign stageClearVec_reqQueue_15_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_15_bitMask;
  assign stageClearVec_reqQueue_15_deq_bits_mask = stageClearVec_reqQueue_dataOut_15_mask;
  assign stageClearVec_reqQueue_15_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_15_groupCounter;
  assign stageClearVec_reqQueue_15_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_15_ffoByOther;
  assign stageClearVec_reqQueue_15_enq_ready = ~_stageClearVec_reqQueue_fifo_15_full;
  wire        stageClearVec_reqQueue_15_deq_ready;
  wire        stageClearVec_WaitReadQueue_15_deq_valid;
  assign stageClearVec_WaitReadQueue_15_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_15_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_15_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_15_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_15_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_15_groupCounter;
  wire [5:0]  out_15_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_15_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_15_ffoByOther;
  wire        out_15_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_15_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_15 = {stageClearVec_WaitReadQueue_15_enq_bits_groupCounter, stageClearVec_WaitReadQueue_15_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_15 = {stageClearVec_WaitReadQueue_15_enq_bits_data, stageClearVec_WaitReadQueue_15_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_15 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_15, stageClearVec_WaitReadQueue_15_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_15 = {stageClearVec_WaitReadQueue_dataIn_hi_15, stageClearVec_WaitReadQueue_dataIn_lo_15};
  assign stageClearVec_WaitReadQueue_dataOut_15_ffoByOther = _stageClearVec_WaitReadQueue_fifo_15_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_15_groupCounter = _stageClearVec_WaitReadQueue_fifo_15_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_15_mask = _stageClearVec_WaitReadQueue_fifo_15_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_15_bitMask = _stageClearVec_WaitReadQueue_fifo_15_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_15_data = _stageClearVec_WaitReadQueue_fifo_15_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_15_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_15_data;
  wire [31:0] stageClearVec_WaitReadQueue_15_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_15_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_15_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_15_mask;
  assign stageClearVec_WaitReadQueue_15_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_15_groupCounter;
  assign stageClearVec_WaitReadQueue_15_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_15_ffoByOther;
  wire        stageClearVec_WaitReadQueue_15_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_15_full;
  wire        stageClearVec_WaitReadQueue_15_enq_valid;
  wire        stageClearVec_WaitReadQueue_15_deq_ready;
  wire        stageClearVec_readReady_15 = ~needWAR | readChannel_15_ready_0;
  assign stageClearVec_WaitReadQueue_15_enq_valid = stageClearVec_reqQueue_15_deq_valid & stageClearVec_readReady_15;
  assign stageClearVec_reqQueue_15_deq_ready = stageClearVec_WaitReadQueue_15_enq_ready & stageClearVec_readReady_15;
  wire        readChannel_15_valid_0 = stageClearVec_reqQueue_15_deq_valid & needWAR & stageClearVec_WaitReadQueue_15_enq_ready;
  wire [4:0]  readChannel_15_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_15_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_15_bits_offset_0 = stageClearVec_reqQueue_15_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_15 = ~needWAR | readResult_15_valid;
  wire [31:0] stageClearVec_WARData_15 = stageClearVec_WaitReadQueue_15_deq_bits_data & stageClearVec_WaitReadQueue_15_deq_bits_bitMask | readResult_15_bits & ~stageClearVec_WaitReadQueue_15_deq_bits_bitMask;
  wire        out_15_valid_0 = stageClearVec_WaitReadQueue_15_deq_valid & stageClearVec_readResultValid_15;
  assign stageClearVec_WaitReadQueue_15_deq_ready = out_15_ready_0 & stageClearVec_readResultValid_15;
  wire [31:0] out_15_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_15 : stageClearVec_WaitReadQueue_15_deq_bits_data;
  wire [3:0]  out_15_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_15_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_15;
  wire        _stageClearVec_T_45 = in_15_ready_0 & in_15_valid_0;
  wire [2:0]  stageClearVec_counterChange_15 = _stageClearVec_T_45 ? 3'h1 : 3'h7;
  wire        stageClearVec_15 = stageClearVec_counter_15 == 3'h0;
  wire        in_16_ready_0 = stageClearVec_reqQueue_16_enq_ready;
  wire        stageClearVec_reqQueue_16_deq_valid;
  assign stageClearVec_reqQueue_16_deq_valid = ~_stageClearVec_reqQueue_fifo_16_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_16_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_16_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_16_enq_bits_data = stageClearVec_reqQueue_16_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_16_mask;
  wire [31:0] stageClearVec_WaitReadQueue_16_enq_bits_bitMask = stageClearVec_reqQueue_16_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_16_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_16_enq_bits_mask = stageClearVec_reqQueue_16_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_16_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_16_enq_bits_groupCounter = stageClearVec_reqQueue_16_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_16_enq_bits_ffoByOther = stageClearVec_reqQueue_16_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_16 = {stageClearVec_reqQueue_16_enq_bits_groupCounter, stageClearVec_reqQueue_16_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_16 = {stageClearVec_reqQueue_16_enq_bits_data, stageClearVec_reqQueue_16_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_16 = {stageClearVec_reqQueue_dataIn_hi_hi_16, stageClearVec_reqQueue_16_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_16 = {stageClearVec_reqQueue_dataIn_hi_16, stageClearVec_reqQueue_dataIn_lo_16};
  assign stageClearVec_reqQueue_dataOut_16_ffoByOther = _stageClearVec_reqQueue_fifo_16_data_out[0];
  assign stageClearVec_reqQueue_dataOut_16_groupCounter = _stageClearVec_reqQueue_fifo_16_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_16_mask = _stageClearVec_reqQueue_fifo_16_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_16_bitMask = _stageClearVec_reqQueue_fifo_16_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_16_data = _stageClearVec_reqQueue_fifo_16_data_out[74:43];
  assign stageClearVec_reqQueue_16_deq_bits_data = stageClearVec_reqQueue_dataOut_16_data;
  assign stageClearVec_reqQueue_16_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_16_bitMask;
  assign stageClearVec_reqQueue_16_deq_bits_mask = stageClearVec_reqQueue_dataOut_16_mask;
  assign stageClearVec_reqQueue_16_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_16_groupCounter;
  assign stageClearVec_reqQueue_16_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_16_ffoByOther;
  assign stageClearVec_reqQueue_16_enq_ready = ~_stageClearVec_reqQueue_fifo_16_full;
  wire        stageClearVec_reqQueue_16_deq_ready;
  wire        stageClearVec_WaitReadQueue_16_deq_valid;
  assign stageClearVec_WaitReadQueue_16_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_16_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_16_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_16_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_16_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_16_groupCounter;
  wire [5:0]  out_16_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_16_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_16_ffoByOther;
  wire        out_16_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_16_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_16 = {stageClearVec_WaitReadQueue_16_enq_bits_groupCounter, stageClearVec_WaitReadQueue_16_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_16 = {stageClearVec_WaitReadQueue_16_enq_bits_data, stageClearVec_WaitReadQueue_16_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_16 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_16, stageClearVec_WaitReadQueue_16_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_16 = {stageClearVec_WaitReadQueue_dataIn_hi_16, stageClearVec_WaitReadQueue_dataIn_lo_16};
  assign stageClearVec_WaitReadQueue_dataOut_16_ffoByOther = _stageClearVec_WaitReadQueue_fifo_16_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_16_groupCounter = _stageClearVec_WaitReadQueue_fifo_16_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_16_mask = _stageClearVec_WaitReadQueue_fifo_16_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_16_bitMask = _stageClearVec_WaitReadQueue_fifo_16_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_16_data = _stageClearVec_WaitReadQueue_fifo_16_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_16_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_16_data;
  wire [31:0] stageClearVec_WaitReadQueue_16_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_16_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_16_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_16_mask;
  assign stageClearVec_WaitReadQueue_16_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_16_groupCounter;
  assign stageClearVec_WaitReadQueue_16_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_16_ffoByOther;
  wire        stageClearVec_WaitReadQueue_16_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_16_full;
  wire        stageClearVec_WaitReadQueue_16_enq_valid;
  wire        stageClearVec_WaitReadQueue_16_deq_ready;
  wire        stageClearVec_readReady_16 = ~needWAR | readChannel_16_ready_0;
  assign stageClearVec_WaitReadQueue_16_enq_valid = stageClearVec_reqQueue_16_deq_valid & stageClearVec_readReady_16;
  assign stageClearVec_reqQueue_16_deq_ready = stageClearVec_WaitReadQueue_16_enq_ready & stageClearVec_readReady_16;
  wire        readChannel_16_valid_0 = stageClearVec_reqQueue_16_deq_valid & needWAR & stageClearVec_WaitReadQueue_16_enq_ready;
  wire [4:0]  readChannel_16_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_16_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_16_bits_offset_0 = stageClearVec_reqQueue_16_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_16 = ~needWAR | readResult_16_valid;
  wire [31:0] stageClearVec_WARData_16 = stageClearVec_WaitReadQueue_16_deq_bits_data & stageClearVec_WaitReadQueue_16_deq_bits_bitMask | readResult_16_bits & ~stageClearVec_WaitReadQueue_16_deq_bits_bitMask;
  wire        out_16_valid_0 = stageClearVec_WaitReadQueue_16_deq_valid & stageClearVec_readResultValid_16;
  assign stageClearVec_WaitReadQueue_16_deq_ready = out_16_ready_0 & stageClearVec_readResultValid_16;
  wire [31:0] out_16_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_16 : stageClearVec_WaitReadQueue_16_deq_bits_data;
  wire [3:0]  out_16_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_16_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_16;
  wire        _stageClearVec_T_48 = in_16_ready_0 & in_16_valid_0;
  wire [2:0]  stageClearVec_counterChange_16 = _stageClearVec_T_48 ? 3'h1 : 3'h7;
  wire        stageClearVec_16 = stageClearVec_counter_16 == 3'h0;
  wire        in_17_ready_0 = stageClearVec_reqQueue_17_enq_ready;
  wire        stageClearVec_reqQueue_17_deq_valid;
  assign stageClearVec_reqQueue_17_deq_valid = ~_stageClearVec_reqQueue_fifo_17_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_17_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_17_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_17_enq_bits_data = stageClearVec_reqQueue_17_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_17_mask;
  wire [31:0] stageClearVec_WaitReadQueue_17_enq_bits_bitMask = stageClearVec_reqQueue_17_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_17_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_17_enq_bits_mask = stageClearVec_reqQueue_17_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_17_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_17_enq_bits_groupCounter = stageClearVec_reqQueue_17_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_17_enq_bits_ffoByOther = stageClearVec_reqQueue_17_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_17 = {stageClearVec_reqQueue_17_enq_bits_groupCounter, stageClearVec_reqQueue_17_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_17 = {stageClearVec_reqQueue_17_enq_bits_data, stageClearVec_reqQueue_17_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_17 = {stageClearVec_reqQueue_dataIn_hi_hi_17, stageClearVec_reqQueue_17_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_17 = {stageClearVec_reqQueue_dataIn_hi_17, stageClearVec_reqQueue_dataIn_lo_17};
  assign stageClearVec_reqQueue_dataOut_17_ffoByOther = _stageClearVec_reqQueue_fifo_17_data_out[0];
  assign stageClearVec_reqQueue_dataOut_17_groupCounter = _stageClearVec_reqQueue_fifo_17_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_17_mask = _stageClearVec_reqQueue_fifo_17_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_17_bitMask = _stageClearVec_reqQueue_fifo_17_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_17_data = _stageClearVec_reqQueue_fifo_17_data_out[74:43];
  assign stageClearVec_reqQueue_17_deq_bits_data = stageClearVec_reqQueue_dataOut_17_data;
  assign stageClearVec_reqQueue_17_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_17_bitMask;
  assign stageClearVec_reqQueue_17_deq_bits_mask = stageClearVec_reqQueue_dataOut_17_mask;
  assign stageClearVec_reqQueue_17_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_17_groupCounter;
  assign stageClearVec_reqQueue_17_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_17_ffoByOther;
  assign stageClearVec_reqQueue_17_enq_ready = ~_stageClearVec_reqQueue_fifo_17_full;
  wire        stageClearVec_reqQueue_17_deq_ready;
  wire        stageClearVec_WaitReadQueue_17_deq_valid;
  assign stageClearVec_WaitReadQueue_17_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_17_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_17_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_17_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_17_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_17_groupCounter;
  wire [5:0]  out_17_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_17_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_17_ffoByOther;
  wire        out_17_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_17_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_17 = {stageClearVec_WaitReadQueue_17_enq_bits_groupCounter, stageClearVec_WaitReadQueue_17_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_17 = {stageClearVec_WaitReadQueue_17_enq_bits_data, stageClearVec_WaitReadQueue_17_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_17 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_17, stageClearVec_WaitReadQueue_17_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_17 = {stageClearVec_WaitReadQueue_dataIn_hi_17, stageClearVec_WaitReadQueue_dataIn_lo_17};
  assign stageClearVec_WaitReadQueue_dataOut_17_ffoByOther = _stageClearVec_WaitReadQueue_fifo_17_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_17_groupCounter = _stageClearVec_WaitReadQueue_fifo_17_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_17_mask = _stageClearVec_WaitReadQueue_fifo_17_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_17_bitMask = _stageClearVec_WaitReadQueue_fifo_17_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_17_data = _stageClearVec_WaitReadQueue_fifo_17_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_17_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_17_data;
  wire [31:0] stageClearVec_WaitReadQueue_17_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_17_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_17_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_17_mask;
  assign stageClearVec_WaitReadQueue_17_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_17_groupCounter;
  assign stageClearVec_WaitReadQueue_17_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_17_ffoByOther;
  wire        stageClearVec_WaitReadQueue_17_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_17_full;
  wire        stageClearVec_WaitReadQueue_17_enq_valid;
  wire        stageClearVec_WaitReadQueue_17_deq_ready;
  wire        stageClearVec_readReady_17 = ~needWAR | readChannel_17_ready_0;
  assign stageClearVec_WaitReadQueue_17_enq_valid = stageClearVec_reqQueue_17_deq_valid & stageClearVec_readReady_17;
  assign stageClearVec_reqQueue_17_deq_ready = stageClearVec_WaitReadQueue_17_enq_ready & stageClearVec_readReady_17;
  wire        readChannel_17_valid_0 = stageClearVec_reqQueue_17_deq_valid & needWAR & stageClearVec_WaitReadQueue_17_enq_ready;
  wire [4:0]  readChannel_17_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_17_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_17_bits_offset_0 = stageClearVec_reqQueue_17_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_17 = ~needWAR | readResult_17_valid;
  wire [31:0] stageClearVec_WARData_17 = stageClearVec_WaitReadQueue_17_deq_bits_data & stageClearVec_WaitReadQueue_17_deq_bits_bitMask | readResult_17_bits & ~stageClearVec_WaitReadQueue_17_deq_bits_bitMask;
  wire        out_17_valid_0 = stageClearVec_WaitReadQueue_17_deq_valid & stageClearVec_readResultValid_17;
  assign stageClearVec_WaitReadQueue_17_deq_ready = out_17_ready_0 & stageClearVec_readResultValid_17;
  wire [31:0] out_17_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_17 : stageClearVec_WaitReadQueue_17_deq_bits_data;
  wire [3:0]  out_17_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_17_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_17;
  wire        _stageClearVec_T_51 = in_17_ready_0 & in_17_valid_0;
  wire [2:0]  stageClearVec_counterChange_17 = _stageClearVec_T_51 ? 3'h1 : 3'h7;
  wire        stageClearVec_17 = stageClearVec_counter_17 == 3'h0;
  wire        in_18_ready_0 = stageClearVec_reqQueue_18_enq_ready;
  wire        stageClearVec_reqQueue_18_deq_valid;
  assign stageClearVec_reqQueue_18_deq_valid = ~_stageClearVec_reqQueue_fifo_18_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_18_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_18_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_18_enq_bits_data = stageClearVec_reqQueue_18_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_18_mask;
  wire [31:0] stageClearVec_WaitReadQueue_18_enq_bits_bitMask = stageClearVec_reqQueue_18_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_18_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_18_enq_bits_mask = stageClearVec_reqQueue_18_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_18_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_18_enq_bits_groupCounter = stageClearVec_reqQueue_18_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_18_enq_bits_ffoByOther = stageClearVec_reqQueue_18_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_18 = {stageClearVec_reqQueue_18_enq_bits_groupCounter, stageClearVec_reqQueue_18_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_18 = {stageClearVec_reqQueue_18_enq_bits_data, stageClearVec_reqQueue_18_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_18 = {stageClearVec_reqQueue_dataIn_hi_hi_18, stageClearVec_reqQueue_18_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_18 = {stageClearVec_reqQueue_dataIn_hi_18, stageClearVec_reqQueue_dataIn_lo_18};
  assign stageClearVec_reqQueue_dataOut_18_ffoByOther = _stageClearVec_reqQueue_fifo_18_data_out[0];
  assign stageClearVec_reqQueue_dataOut_18_groupCounter = _stageClearVec_reqQueue_fifo_18_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_18_mask = _stageClearVec_reqQueue_fifo_18_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_18_bitMask = _stageClearVec_reqQueue_fifo_18_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_18_data = _stageClearVec_reqQueue_fifo_18_data_out[74:43];
  assign stageClearVec_reqQueue_18_deq_bits_data = stageClearVec_reqQueue_dataOut_18_data;
  assign stageClearVec_reqQueue_18_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_18_bitMask;
  assign stageClearVec_reqQueue_18_deq_bits_mask = stageClearVec_reqQueue_dataOut_18_mask;
  assign stageClearVec_reqQueue_18_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_18_groupCounter;
  assign stageClearVec_reqQueue_18_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_18_ffoByOther;
  assign stageClearVec_reqQueue_18_enq_ready = ~_stageClearVec_reqQueue_fifo_18_full;
  wire        stageClearVec_reqQueue_18_deq_ready;
  wire        stageClearVec_WaitReadQueue_18_deq_valid;
  assign stageClearVec_WaitReadQueue_18_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_18_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_18_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_18_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_18_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_18_groupCounter;
  wire [5:0]  out_18_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_18_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_18_ffoByOther;
  wire        out_18_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_18_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_18 = {stageClearVec_WaitReadQueue_18_enq_bits_groupCounter, stageClearVec_WaitReadQueue_18_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_18 = {stageClearVec_WaitReadQueue_18_enq_bits_data, stageClearVec_WaitReadQueue_18_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_18 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_18, stageClearVec_WaitReadQueue_18_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_18 = {stageClearVec_WaitReadQueue_dataIn_hi_18, stageClearVec_WaitReadQueue_dataIn_lo_18};
  assign stageClearVec_WaitReadQueue_dataOut_18_ffoByOther = _stageClearVec_WaitReadQueue_fifo_18_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_18_groupCounter = _stageClearVec_WaitReadQueue_fifo_18_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_18_mask = _stageClearVec_WaitReadQueue_fifo_18_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_18_bitMask = _stageClearVec_WaitReadQueue_fifo_18_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_18_data = _stageClearVec_WaitReadQueue_fifo_18_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_18_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_18_data;
  wire [31:0] stageClearVec_WaitReadQueue_18_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_18_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_18_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_18_mask;
  assign stageClearVec_WaitReadQueue_18_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_18_groupCounter;
  assign stageClearVec_WaitReadQueue_18_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_18_ffoByOther;
  wire        stageClearVec_WaitReadQueue_18_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_18_full;
  wire        stageClearVec_WaitReadQueue_18_enq_valid;
  wire        stageClearVec_WaitReadQueue_18_deq_ready;
  wire        stageClearVec_readReady_18 = ~needWAR | readChannel_18_ready_0;
  assign stageClearVec_WaitReadQueue_18_enq_valid = stageClearVec_reqQueue_18_deq_valid & stageClearVec_readReady_18;
  assign stageClearVec_reqQueue_18_deq_ready = stageClearVec_WaitReadQueue_18_enq_ready & stageClearVec_readReady_18;
  wire        readChannel_18_valid_0 = stageClearVec_reqQueue_18_deq_valid & needWAR & stageClearVec_WaitReadQueue_18_enq_ready;
  wire [4:0]  readChannel_18_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_18_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_18_bits_offset_0 = stageClearVec_reqQueue_18_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_18 = ~needWAR | readResult_18_valid;
  wire [31:0] stageClearVec_WARData_18 = stageClearVec_WaitReadQueue_18_deq_bits_data & stageClearVec_WaitReadQueue_18_deq_bits_bitMask | readResult_18_bits & ~stageClearVec_WaitReadQueue_18_deq_bits_bitMask;
  wire        out_18_valid_0 = stageClearVec_WaitReadQueue_18_deq_valid & stageClearVec_readResultValid_18;
  assign stageClearVec_WaitReadQueue_18_deq_ready = out_18_ready_0 & stageClearVec_readResultValid_18;
  wire [31:0] out_18_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_18 : stageClearVec_WaitReadQueue_18_deq_bits_data;
  wire [3:0]  out_18_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_18_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_18;
  wire        _stageClearVec_T_54 = in_18_ready_0 & in_18_valid_0;
  wire [2:0]  stageClearVec_counterChange_18 = _stageClearVec_T_54 ? 3'h1 : 3'h7;
  wire        stageClearVec_18 = stageClearVec_counter_18 == 3'h0;
  wire        in_19_ready_0 = stageClearVec_reqQueue_19_enq_ready;
  wire        stageClearVec_reqQueue_19_deq_valid;
  assign stageClearVec_reqQueue_19_deq_valid = ~_stageClearVec_reqQueue_fifo_19_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_19_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_19_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_19_enq_bits_data = stageClearVec_reqQueue_19_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_19_mask;
  wire [31:0] stageClearVec_WaitReadQueue_19_enq_bits_bitMask = stageClearVec_reqQueue_19_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_19_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_19_enq_bits_mask = stageClearVec_reqQueue_19_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_19_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_19_enq_bits_groupCounter = stageClearVec_reqQueue_19_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_19_enq_bits_ffoByOther = stageClearVec_reqQueue_19_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_19 = {stageClearVec_reqQueue_19_enq_bits_groupCounter, stageClearVec_reqQueue_19_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_19 = {stageClearVec_reqQueue_19_enq_bits_data, stageClearVec_reqQueue_19_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_19 = {stageClearVec_reqQueue_dataIn_hi_hi_19, stageClearVec_reqQueue_19_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_19 = {stageClearVec_reqQueue_dataIn_hi_19, stageClearVec_reqQueue_dataIn_lo_19};
  assign stageClearVec_reqQueue_dataOut_19_ffoByOther = _stageClearVec_reqQueue_fifo_19_data_out[0];
  assign stageClearVec_reqQueue_dataOut_19_groupCounter = _stageClearVec_reqQueue_fifo_19_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_19_mask = _stageClearVec_reqQueue_fifo_19_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_19_bitMask = _stageClearVec_reqQueue_fifo_19_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_19_data = _stageClearVec_reqQueue_fifo_19_data_out[74:43];
  assign stageClearVec_reqQueue_19_deq_bits_data = stageClearVec_reqQueue_dataOut_19_data;
  assign stageClearVec_reqQueue_19_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_19_bitMask;
  assign stageClearVec_reqQueue_19_deq_bits_mask = stageClearVec_reqQueue_dataOut_19_mask;
  assign stageClearVec_reqQueue_19_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_19_groupCounter;
  assign stageClearVec_reqQueue_19_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_19_ffoByOther;
  assign stageClearVec_reqQueue_19_enq_ready = ~_stageClearVec_reqQueue_fifo_19_full;
  wire        stageClearVec_reqQueue_19_deq_ready;
  wire        stageClearVec_WaitReadQueue_19_deq_valid;
  assign stageClearVec_WaitReadQueue_19_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_19_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_19_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_19_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_19_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_19_groupCounter;
  wire [5:0]  out_19_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_19_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_19_ffoByOther;
  wire        out_19_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_19_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_19 = {stageClearVec_WaitReadQueue_19_enq_bits_groupCounter, stageClearVec_WaitReadQueue_19_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_19 = {stageClearVec_WaitReadQueue_19_enq_bits_data, stageClearVec_WaitReadQueue_19_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_19 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_19, stageClearVec_WaitReadQueue_19_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_19 = {stageClearVec_WaitReadQueue_dataIn_hi_19, stageClearVec_WaitReadQueue_dataIn_lo_19};
  assign stageClearVec_WaitReadQueue_dataOut_19_ffoByOther = _stageClearVec_WaitReadQueue_fifo_19_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_19_groupCounter = _stageClearVec_WaitReadQueue_fifo_19_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_19_mask = _stageClearVec_WaitReadQueue_fifo_19_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_19_bitMask = _stageClearVec_WaitReadQueue_fifo_19_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_19_data = _stageClearVec_WaitReadQueue_fifo_19_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_19_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_19_data;
  wire [31:0] stageClearVec_WaitReadQueue_19_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_19_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_19_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_19_mask;
  assign stageClearVec_WaitReadQueue_19_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_19_groupCounter;
  assign stageClearVec_WaitReadQueue_19_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_19_ffoByOther;
  wire        stageClearVec_WaitReadQueue_19_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_19_full;
  wire        stageClearVec_WaitReadQueue_19_enq_valid;
  wire        stageClearVec_WaitReadQueue_19_deq_ready;
  wire        stageClearVec_readReady_19 = ~needWAR | readChannel_19_ready_0;
  assign stageClearVec_WaitReadQueue_19_enq_valid = stageClearVec_reqQueue_19_deq_valid & stageClearVec_readReady_19;
  assign stageClearVec_reqQueue_19_deq_ready = stageClearVec_WaitReadQueue_19_enq_ready & stageClearVec_readReady_19;
  wire        readChannel_19_valid_0 = stageClearVec_reqQueue_19_deq_valid & needWAR & stageClearVec_WaitReadQueue_19_enq_ready;
  wire [4:0]  readChannel_19_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_19_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_19_bits_offset_0 = stageClearVec_reqQueue_19_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_19 = ~needWAR | readResult_19_valid;
  wire [31:0] stageClearVec_WARData_19 = stageClearVec_WaitReadQueue_19_deq_bits_data & stageClearVec_WaitReadQueue_19_deq_bits_bitMask | readResult_19_bits & ~stageClearVec_WaitReadQueue_19_deq_bits_bitMask;
  wire        out_19_valid_0 = stageClearVec_WaitReadQueue_19_deq_valid & stageClearVec_readResultValid_19;
  assign stageClearVec_WaitReadQueue_19_deq_ready = out_19_ready_0 & stageClearVec_readResultValid_19;
  wire [31:0] out_19_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_19 : stageClearVec_WaitReadQueue_19_deq_bits_data;
  wire [3:0]  out_19_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_19_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_19;
  wire        _stageClearVec_T_57 = in_19_ready_0 & in_19_valid_0;
  wire [2:0]  stageClearVec_counterChange_19 = _stageClearVec_T_57 ? 3'h1 : 3'h7;
  wire        stageClearVec_19 = stageClearVec_counter_19 == 3'h0;
  wire        in_20_ready_0 = stageClearVec_reqQueue_20_enq_ready;
  wire        stageClearVec_reqQueue_20_deq_valid;
  assign stageClearVec_reqQueue_20_deq_valid = ~_stageClearVec_reqQueue_fifo_20_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_20_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_20_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_20_enq_bits_data = stageClearVec_reqQueue_20_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_20_mask;
  wire [31:0] stageClearVec_WaitReadQueue_20_enq_bits_bitMask = stageClearVec_reqQueue_20_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_20_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_20_enq_bits_mask = stageClearVec_reqQueue_20_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_20_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_20_enq_bits_groupCounter = stageClearVec_reqQueue_20_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_20_enq_bits_ffoByOther = stageClearVec_reqQueue_20_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_20 = {stageClearVec_reqQueue_20_enq_bits_groupCounter, stageClearVec_reqQueue_20_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_20 = {stageClearVec_reqQueue_20_enq_bits_data, stageClearVec_reqQueue_20_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_20 = {stageClearVec_reqQueue_dataIn_hi_hi_20, stageClearVec_reqQueue_20_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_20 = {stageClearVec_reqQueue_dataIn_hi_20, stageClearVec_reqQueue_dataIn_lo_20};
  assign stageClearVec_reqQueue_dataOut_20_ffoByOther = _stageClearVec_reqQueue_fifo_20_data_out[0];
  assign stageClearVec_reqQueue_dataOut_20_groupCounter = _stageClearVec_reqQueue_fifo_20_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_20_mask = _stageClearVec_reqQueue_fifo_20_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_20_bitMask = _stageClearVec_reqQueue_fifo_20_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_20_data = _stageClearVec_reqQueue_fifo_20_data_out[74:43];
  assign stageClearVec_reqQueue_20_deq_bits_data = stageClearVec_reqQueue_dataOut_20_data;
  assign stageClearVec_reqQueue_20_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_20_bitMask;
  assign stageClearVec_reqQueue_20_deq_bits_mask = stageClearVec_reqQueue_dataOut_20_mask;
  assign stageClearVec_reqQueue_20_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_20_groupCounter;
  assign stageClearVec_reqQueue_20_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_20_ffoByOther;
  assign stageClearVec_reqQueue_20_enq_ready = ~_stageClearVec_reqQueue_fifo_20_full;
  wire        stageClearVec_reqQueue_20_deq_ready;
  wire        stageClearVec_WaitReadQueue_20_deq_valid;
  assign stageClearVec_WaitReadQueue_20_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_20_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_20_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_20_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_20_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_20_groupCounter;
  wire [5:0]  out_20_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_20_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_20_ffoByOther;
  wire        out_20_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_20_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_20 = {stageClearVec_WaitReadQueue_20_enq_bits_groupCounter, stageClearVec_WaitReadQueue_20_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_20 = {stageClearVec_WaitReadQueue_20_enq_bits_data, stageClearVec_WaitReadQueue_20_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_20 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_20, stageClearVec_WaitReadQueue_20_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_20 = {stageClearVec_WaitReadQueue_dataIn_hi_20, stageClearVec_WaitReadQueue_dataIn_lo_20};
  assign stageClearVec_WaitReadQueue_dataOut_20_ffoByOther = _stageClearVec_WaitReadQueue_fifo_20_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_20_groupCounter = _stageClearVec_WaitReadQueue_fifo_20_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_20_mask = _stageClearVec_WaitReadQueue_fifo_20_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_20_bitMask = _stageClearVec_WaitReadQueue_fifo_20_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_20_data = _stageClearVec_WaitReadQueue_fifo_20_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_20_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_20_data;
  wire [31:0] stageClearVec_WaitReadQueue_20_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_20_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_20_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_20_mask;
  assign stageClearVec_WaitReadQueue_20_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_20_groupCounter;
  assign stageClearVec_WaitReadQueue_20_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_20_ffoByOther;
  wire        stageClearVec_WaitReadQueue_20_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_20_full;
  wire        stageClearVec_WaitReadQueue_20_enq_valid;
  wire        stageClearVec_WaitReadQueue_20_deq_ready;
  wire        stageClearVec_readReady_20 = ~needWAR | readChannel_20_ready_0;
  assign stageClearVec_WaitReadQueue_20_enq_valid = stageClearVec_reqQueue_20_deq_valid & stageClearVec_readReady_20;
  assign stageClearVec_reqQueue_20_deq_ready = stageClearVec_WaitReadQueue_20_enq_ready & stageClearVec_readReady_20;
  wire        readChannel_20_valid_0 = stageClearVec_reqQueue_20_deq_valid & needWAR & stageClearVec_WaitReadQueue_20_enq_ready;
  wire [4:0]  readChannel_20_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_20_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_20_bits_offset_0 = stageClearVec_reqQueue_20_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_20 = ~needWAR | readResult_20_valid;
  wire [31:0] stageClearVec_WARData_20 = stageClearVec_WaitReadQueue_20_deq_bits_data & stageClearVec_WaitReadQueue_20_deq_bits_bitMask | readResult_20_bits & ~stageClearVec_WaitReadQueue_20_deq_bits_bitMask;
  wire        out_20_valid_0 = stageClearVec_WaitReadQueue_20_deq_valid & stageClearVec_readResultValid_20;
  assign stageClearVec_WaitReadQueue_20_deq_ready = out_20_ready_0 & stageClearVec_readResultValid_20;
  wire [31:0] out_20_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_20 : stageClearVec_WaitReadQueue_20_deq_bits_data;
  wire [3:0]  out_20_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_20_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_20;
  wire        _stageClearVec_T_60 = in_20_ready_0 & in_20_valid_0;
  wire [2:0]  stageClearVec_counterChange_20 = _stageClearVec_T_60 ? 3'h1 : 3'h7;
  wire        stageClearVec_20 = stageClearVec_counter_20 == 3'h0;
  wire        in_21_ready_0 = stageClearVec_reqQueue_21_enq_ready;
  wire        stageClearVec_reqQueue_21_deq_valid;
  assign stageClearVec_reqQueue_21_deq_valid = ~_stageClearVec_reqQueue_fifo_21_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_21_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_21_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_21_enq_bits_data = stageClearVec_reqQueue_21_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_21_mask;
  wire [31:0] stageClearVec_WaitReadQueue_21_enq_bits_bitMask = stageClearVec_reqQueue_21_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_21_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_21_enq_bits_mask = stageClearVec_reqQueue_21_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_21_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_21_enq_bits_groupCounter = stageClearVec_reqQueue_21_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_21_enq_bits_ffoByOther = stageClearVec_reqQueue_21_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_21 = {stageClearVec_reqQueue_21_enq_bits_groupCounter, stageClearVec_reqQueue_21_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_21 = {stageClearVec_reqQueue_21_enq_bits_data, stageClearVec_reqQueue_21_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_21 = {stageClearVec_reqQueue_dataIn_hi_hi_21, stageClearVec_reqQueue_21_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_21 = {stageClearVec_reqQueue_dataIn_hi_21, stageClearVec_reqQueue_dataIn_lo_21};
  assign stageClearVec_reqQueue_dataOut_21_ffoByOther = _stageClearVec_reqQueue_fifo_21_data_out[0];
  assign stageClearVec_reqQueue_dataOut_21_groupCounter = _stageClearVec_reqQueue_fifo_21_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_21_mask = _stageClearVec_reqQueue_fifo_21_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_21_bitMask = _stageClearVec_reqQueue_fifo_21_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_21_data = _stageClearVec_reqQueue_fifo_21_data_out[74:43];
  assign stageClearVec_reqQueue_21_deq_bits_data = stageClearVec_reqQueue_dataOut_21_data;
  assign stageClearVec_reqQueue_21_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_21_bitMask;
  assign stageClearVec_reqQueue_21_deq_bits_mask = stageClearVec_reqQueue_dataOut_21_mask;
  assign stageClearVec_reqQueue_21_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_21_groupCounter;
  assign stageClearVec_reqQueue_21_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_21_ffoByOther;
  assign stageClearVec_reqQueue_21_enq_ready = ~_stageClearVec_reqQueue_fifo_21_full;
  wire        stageClearVec_reqQueue_21_deq_ready;
  wire        stageClearVec_WaitReadQueue_21_deq_valid;
  assign stageClearVec_WaitReadQueue_21_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_21_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_21_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_21_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_21_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_21_groupCounter;
  wire [5:0]  out_21_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_21_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_21_ffoByOther;
  wire        out_21_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_21_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_21 = {stageClearVec_WaitReadQueue_21_enq_bits_groupCounter, stageClearVec_WaitReadQueue_21_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_21 = {stageClearVec_WaitReadQueue_21_enq_bits_data, stageClearVec_WaitReadQueue_21_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_21 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_21, stageClearVec_WaitReadQueue_21_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_21 = {stageClearVec_WaitReadQueue_dataIn_hi_21, stageClearVec_WaitReadQueue_dataIn_lo_21};
  assign stageClearVec_WaitReadQueue_dataOut_21_ffoByOther = _stageClearVec_WaitReadQueue_fifo_21_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_21_groupCounter = _stageClearVec_WaitReadQueue_fifo_21_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_21_mask = _stageClearVec_WaitReadQueue_fifo_21_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_21_bitMask = _stageClearVec_WaitReadQueue_fifo_21_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_21_data = _stageClearVec_WaitReadQueue_fifo_21_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_21_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_21_data;
  wire [31:0] stageClearVec_WaitReadQueue_21_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_21_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_21_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_21_mask;
  assign stageClearVec_WaitReadQueue_21_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_21_groupCounter;
  assign stageClearVec_WaitReadQueue_21_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_21_ffoByOther;
  wire        stageClearVec_WaitReadQueue_21_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_21_full;
  wire        stageClearVec_WaitReadQueue_21_enq_valid;
  wire        stageClearVec_WaitReadQueue_21_deq_ready;
  wire        stageClearVec_readReady_21 = ~needWAR | readChannel_21_ready_0;
  assign stageClearVec_WaitReadQueue_21_enq_valid = stageClearVec_reqQueue_21_deq_valid & stageClearVec_readReady_21;
  assign stageClearVec_reqQueue_21_deq_ready = stageClearVec_WaitReadQueue_21_enq_ready & stageClearVec_readReady_21;
  wire        readChannel_21_valid_0 = stageClearVec_reqQueue_21_deq_valid & needWAR & stageClearVec_WaitReadQueue_21_enq_ready;
  wire [4:0]  readChannel_21_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_21_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_21_bits_offset_0 = stageClearVec_reqQueue_21_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_21 = ~needWAR | readResult_21_valid;
  wire [31:0] stageClearVec_WARData_21 = stageClearVec_WaitReadQueue_21_deq_bits_data & stageClearVec_WaitReadQueue_21_deq_bits_bitMask | readResult_21_bits & ~stageClearVec_WaitReadQueue_21_deq_bits_bitMask;
  wire        out_21_valid_0 = stageClearVec_WaitReadQueue_21_deq_valid & stageClearVec_readResultValid_21;
  assign stageClearVec_WaitReadQueue_21_deq_ready = out_21_ready_0 & stageClearVec_readResultValid_21;
  wire [31:0] out_21_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_21 : stageClearVec_WaitReadQueue_21_deq_bits_data;
  wire [3:0]  out_21_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_21_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_21;
  wire        _stageClearVec_T_63 = in_21_ready_0 & in_21_valid_0;
  wire [2:0]  stageClearVec_counterChange_21 = _stageClearVec_T_63 ? 3'h1 : 3'h7;
  wire        stageClearVec_21 = stageClearVec_counter_21 == 3'h0;
  wire        in_22_ready_0 = stageClearVec_reqQueue_22_enq_ready;
  wire        stageClearVec_reqQueue_22_deq_valid;
  assign stageClearVec_reqQueue_22_deq_valid = ~_stageClearVec_reqQueue_fifo_22_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_22_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_22_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_22_enq_bits_data = stageClearVec_reqQueue_22_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_22_mask;
  wire [31:0] stageClearVec_WaitReadQueue_22_enq_bits_bitMask = stageClearVec_reqQueue_22_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_22_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_22_enq_bits_mask = stageClearVec_reqQueue_22_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_22_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_22_enq_bits_groupCounter = stageClearVec_reqQueue_22_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_22_enq_bits_ffoByOther = stageClearVec_reqQueue_22_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_22 = {stageClearVec_reqQueue_22_enq_bits_groupCounter, stageClearVec_reqQueue_22_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_22 = {stageClearVec_reqQueue_22_enq_bits_data, stageClearVec_reqQueue_22_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_22 = {stageClearVec_reqQueue_dataIn_hi_hi_22, stageClearVec_reqQueue_22_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_22 = {stageClearVec_reqQueue_dataIn_hi_22, stageClearVec_reqQueue_dataIn_lo_22};
  assign stageClearVec_reqQueue_dataOut_22_ffoByOther = _stageClearVec_reqQueue_fifo_22_data_out[0];
  assign stageClearVec_reqQueue_dataOut_22_groupCounter = _stageClearVec_reqQueue_fifo_22_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_22_mask = _stageClearVec_reqQueue_fifo_22_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_22_bitMask = _stageClearVec_reqQueue_fifo_22_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_22_data = _stageClearVec_reqQueue_fifo_22_data_out[74:43];
  assign stageClearVec_reqQueue_22_deq_bits_data = stageClearVec_reqQueue_dataOut_22_data;
  assign stageClearVec_reqQueue_22_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_22_bitMask;
  assign stageClearVec_reqQueue_22_deq_bits_mask = stageClearVec_reqQueue_dataOut_22_mask;
  assign stageClearVec_reqQueue_22_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_22_groupCounter;
  assign stageClearVec_reqQueue_22_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_22_ffoByOther;
  assign stageClearVec_reqQueue_22_enq_ready = ~_stageClearVec_reqQueue_fifo_22_full;
  wire        stageClearVec_reqQueue_22_deq_ready;
  wire        stageClearVec_WaitReadQueue_22_deq_valid;
  assign stageClearVec_WaitReadQueue_22_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_22_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_22_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_22_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_22_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_22_groupCounter;
  wire [5:0]  out_22_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_22_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_22_ffoByOther;
  wire        out_22_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_22_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_22 = {stageClearVec_WaitReadQueue_22_enq_bits_groupCounter, stageClearVec_WaitReadQueue_22_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_22 = {stageClearVec_WaitReadQueue_22_enq_bits_data, stageClearVec_WaitReadQueue_22_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_22 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_22, stageClearVec_WaitReadQueue_22_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_22 = {stageClearVec_WaitReadQueue_dataIn_hi_22, stageClearVec_WaitReadQueue_dataIn_lo_22};
  assign stageClearVec_WaitReadQueue_dataOut_22_ffoByOther = _stageClearVec_WaitReadQueue_fifo_22_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_22_groupCounter = _stageClearVec_WaitReadQueue_fifo_22_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_22_mask = _stageClearVec_WaitReadQueue_fifo_22_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_22_bitMask = _stageClearVec_WaitReadQueue_fifo_22_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_22_data = _stageClearVec_WaitReadQueue_fifo_22_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_22_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_22_data;
  wire [31:0] stageClearVec_WaitReadQueue_22_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_22_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_22_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_22_mask;
  assign stageClearVec_WaitReadQueue_22_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_22_groupCounter;
  assign stageClearVec_WaitReadQueue_22_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_22_ffoByOther;
  wire        stageClearVec_WaitReadQueue_22_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_22_full;
  wire        stageClearVec_WaitReadQueue_22_enq_valid;
  wire        stageClearVec_WaitReadQueue_22_deq_ready;
  wire        stageClearVec_readReady_22 = ~needWAR | readChannel_22_ready_0;
  assign stageClearVec_WaitReadQueue_22_enq_valid = stageClearVec_reqQueue_22_deq_valid & stageClearVec_readReady_22;
  assign stageClearVec_reqQueue_22_deq_ready = stageClearVec_WaitReadQueue_22_enq_ready & stageClearVec_readReady_22;
  wire        readChannel_22_valid_0 = stageClearVec_reqQueue_22_deq_valid & needWAR & stageClearVec_WaitReadQueue_22_enq_ready;
  wire [4:0]  readChannel_22_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_22_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_22_bits_offset_0 = stageClearVec_reqQueue_22_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_22 = ~needWAR | readResult_22_valid;
  wire [31:0] stageClearVec_WARData_22 = stageClearVec_WaitReadQueue_22_deq_bits_data & stageClearVec_WaitReadQueue_22_deq_bits_bitMask | readResult_22_bits & ~stageClearVec_WaitReadQueue_22_deq_bits_bitMask;
  wire        out_22_valid_0 = stageClearVec_WaitReadQueue_22_deq_valid & stageClearVec_readResultValid_22;
  assign stageClearVec_WaitReadQueue_22_deq_ready = out_22_ready_0 & stageClearVec_readResultValid_22;
  wire [31:0] out_22_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_22 : stageClearVec_WaitReadQueue_22_deq_bits_data;
  wire [3:0]  out_22_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_22_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_22;
  wire        _stageClearVec_T_66 = in_22_ready_0 & in_22_valid_0;
  wire [2:0]  stageClearVec_counterChange_22 = _stageClearVec_T_66 ? 3'h1 : 3'h7;
  wire        stageClearVec_22 = stageClearVec_counter_22 == 3'h0;
  wire        in_23_ready_0 = stageClearVec_reqQueue_23_enq_ready;
  wire        stageClearVec_reqQueue_23_deq_valid;
  assign stageClearVec_reqQueue_23_deq_valid = ~_stageClearVec_reqQueue_fifo_23_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_23_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_23_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_23_enq_bits_data = stageClearVec_reqQueue_23_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_23_mask;
  wire [31:0] stageClearVec_WaitReadQueue_23_enq_bits_bitMask = stageClearVec_reqQueue_23_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_23_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_23_enq_bits_mask = stageClearVec_reqQueue_23_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_23_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_23_enq_bits_groupCounter = stageClearVec_reqQueue_23_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_23_enq_bits_ffoByOther = stageClearVec_reqQueue_23_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_23 = {stageClearVec_reqQueue_23_enq_bits_groupCounter, stageClearVec_reqQueue_23_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_23 = {stageClearVec_reqQueue_23_enq_bits_data, stageClearVec_reqQueue_23_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_23 = {stageClearVec_reqQueue_dataIn_hi_hi_23, stageClearVec_reqQueue_23_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_23 = {stageClearVec_reqQueue_dataIn_hi_23, stageClearVec_reqQueue_dataIn_lo_23};
  assign stageClearVec_reqQueue_dataOut_23_ffoByOther = _stageClearVec_reqQueue_fifo_23_data_out[0];
  assign stageClearVec_reqQueue_dataOut_23_groupCounter = _stageClearVec_reqQueue_fifo_23_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_23_mask = _stageClearVec_reqQueue_fifo_23_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_23_bitMask = _stageClearVec_reqQueue_fifo_23_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_23_data = _stageClearVec_reqQueue_fifo_23_data_out[74:43];
  assign stageClearVec_reqQueue_23_deq_bits_data = stageClearVec_reqQueue_dataOut_23_data;
  assign stageClearVec_reqQueue_23_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_23_bitMask;
  assign stageClearVec_reqQueue_23_deq_bits_mask = stageClearVec_reqQueue_dataOut_23_mask;
  assign stageClearVec_reqQueue_23_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_23_groupCounter;
  assign stageClearVec_reqQueue_23_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_23_ffoByOther;
  assign stageClearVec_reqQueue_23_enq_ready = ~_stageClearVec_reqQueue_fifo_23_full;
  wire        stageClearVec_reqQueue_23_deq_ready;
  wire        stageClearVec_WaitReadQueue_23_deq_valid;
  assign stageClearVec_WaitReadQueue_23_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_23_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_23_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_23_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_23_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_23_groupCounter;
  wire [5:0]  out_23_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_23_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_23_ffoByOther;
  wire        out_23_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_23_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_23 = {stageClearVec_WaitReadQueue_23_enq_bits_groupCounter, stageClearVec_WaitReadQueue_23_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_23 = {stageClearVec_WaitReadQueue_23_enq_bits_data, stageClearVec_WaitReadQueue_23_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_23 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_23, stageClearVec_WaitReadQueue_23_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_23 = {stageClearVec_WaitReadQueue_dataIn_hi_23, stageClearVec_WaitReadQueue_dataIn_lo_23};
  assign stageClearVec_WaitReadQueue_dataOut_23_ffoByOther = _stageClearVec_WaitReadQueue_fifo_23_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_23_groupCounter = _stageClearVec_WaitReadQueue_fifo_23_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_23_mask = _stageClearVec_WaitReadQueue_fifo_23_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_23_bitMask = _stageClearVec_WaitReadQueue_fifo_23_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_23_data = _stageClearVec_WaitReadQueue_fifo_23_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_23_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_23_data;
  wire [31:0] stageClearVec_WaitReadQueue_23_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_23_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_23_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_23_mask;
  assign stageClearVec_WaitReadQueue_23_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_23_groupCounter;
  assign stageClearVec_WaitReadQueue_23_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_23_ffoByOther;
  wire        stageClearVec_WaitReadQueue_23_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_23_full;
  wire        stageClearVec_WaitReadQueue_23_enq_valid;
  wire        stageClearVec_WaitReadQueue_23_deq_ready;
  wire        stageClearVec_readReady_23 = ~needWAR | readChannel_23_ready_0;
  assign stageClearVec_WaitReadQueue_23_enq_valid = stageClearVec_reqQueue_23_deq_valid & stageClearVec_readReady_23;
  assign stageClearVec_reqQueue_23_deq_ready = stageClearVec_WaitReadQueue_23_enq_ready & stageClearVec_readReady_23;
  wire        readChannel_23_valid_0 = stageClearVec_reqQueue_23_deq_valid & needWAR & stageClearVec_WaitReadQueue_23_enq_ready;
  wire [4:0]  readChannel_23_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_23_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_23_bits_offset_0 = stageClearVec_reqQueue_23_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_23 = ~needWAR | readResult_23_valid;
  wire [31:0] stageClearVec_WARData_23 = stageClearVec_WaitReadQueue_23_deq_bits_data & stageClearVec_WaitReadQueue_23_deq_bits_bitMask | readResult_23_bits & ~stageClearVec_WaitReadQueue_23_deq_bits_bitMask;
  wire        out_23_valid_0 = stageClearVec_WaitReadQueue_23_deq_valid & stageClearVec_readResultValid_23;
  assign stageClearVec_WaitReadQueue_23_deq_ready = out_23_ready_0 & stageClearVec_readResultValid_23;
  wire [31:0] out_23_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_23 : stageClearVec_WaitReadQueue_23_deq_bits_data;
  wire [3:0]  out_23_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_23_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_23;
  wire        _stageClearVec_T_69 = in_23_ready_0 & in_23_valid_0;
  wire [2:0]  stageClearVec_counterChange_23 = _stageClearVec_T_69 ? 3'h1 : 3'h7;
  wire        stageClearVec_23 = stageClearVec_counter_23 == 3'h0;
  wire        in_24_ready_0 = stageClearVec_reqQueue_24_enq_ready;
  wire        stageClearVec_reqQueue_24_deq_valid;
  assign stageClearVec_reqQueue_24_deq_valid = ~_stageClearVec_reqQueue_fifo_24_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_24_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_24_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_24_enq_bits_data = stageClearVec_reqQueue_24_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_24_mask;
  wire [31:0] stageClearVec_WaitReadQueue_24_enq_bits_bitMask = stageClearVec_reqQueue_24_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_24_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_24_enq_bits_mask = stageClearVec_reqQueue_24_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_24_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_24_enq_bits_groupCounter = stageClearVec_reqQueue_24_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_24_enq_bits_ffoByOther = stageClearVec_reqQueue_24_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_24 = {stageClearVec_reqQueue_24_enq_bits_groupCounter, stageClearVec_reqQueue_24_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_24 = {stageClearVec_reqQueue_24_enq_bits_data, stageClearVec_reqQueue_24_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_24 = {stageClearVec_reqQueue_dataIn_hi_hi_24, stageClearVec_reqQueue_24_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_24 = {stageClearVec_reqQueue_dataIn_hi_24, stageClearVec_reqQueue_dataIn_lo_24};
  assign stageClearVec_reqQueue_dataOut_24_ffoByOther = _stageClearVec_reqQueue_fifo_24_data_out[0];
  assign stageClearVec_reqQueue_dataOut_24_groupCounter = _stageClearVec_reqQueue_fifo_24_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_24_mask = _stageClearVec_reqQueue_fifo_24_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_24_bitMask = _stageClearVec_reqQueue_fifo_24_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_24_data = _stageClearVec_reqQueue_fifo_24_data_out[74:43];
  assign stageClearVec_reqQueue_24_deq_bits_data = stageClearVec_reqQueue_dataOut_24_data;
  assign stageClearVec_reqQueue_24_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_24_bitMask;
  assign stageClearVec_reqQueue_24_deq_bits_mask = stageClearVec_reqQueue_dataOut_24_mask;
  assign stageClearVec_reqQueue_24_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_24_groupCounter;
  assign stageClearVec_reqQueue_24_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_24_ffoByOther;
  assign stageClearVec_reqQueue_24_enq_ready = ~_stageClearVec_reqQueue_fifo_24_full;
  wire        stageClearVec_reqQueue_24_deq_ready;
  wire        stageClearVec_WaitReadQueue_24_deq_valid;
  assign stageClearVec_WaitReadQueue_24_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_24_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_24_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_24_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_24_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_24_groupCounter;
  wire [5:0]  out_24_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_24_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_24_ffoByOther;
  wire        out_24_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_24_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_24 = {stageClearVec_WaitReadQueue_24_enq_bits_groupCounter, stageClearVec_WaitReadQueue_24_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_24 = {stageClearVec_WaitReadQueue_24_enq_bits_data, stageClearVec_WaitReadQueue_24_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_24 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_24, stageClearVec_WaitReadQueue_24_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_24 = {stageClearVec_WaitReadQueue_dataIn_hi_24, stageClearVec_WaitReadQueue_dataIn_lo_24};
  assign stageClearVec_WaitReadQueue_dataOut_24_ffoByOther = _stageClearVec_WaitReadQueue_fifo_24_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_24_groupCounter = _stageClearVec_WaitReadQueue_fifo_24_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_24_mask = _stageClearVec_WaitReadQueue_fifo_24_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_24_bitMask = _stageClearVec_WaitReadQueue_fifo_24_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_24_data = _stageClearVec_WaitReadQueue_fifo_24_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_24_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_24_data;
  wire [31:0] stageClearVec_WaitReadQueue_24_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_24_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_24_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_24_mask;
  assign stageClearVec_WaitReadQueue_24_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_24_groupCounter;
  assign stageClearVec_WaitReadQueue_24_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_24_ffoByOther;
  wire        stageClearVec_WaitReadQueue_24_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_24_full;
  wire        stageClearVec_WaitReadQueue_24_enq_valid;
  wire        stageClearVec_WaitReadQueue_24_deq_ready;
  wire        stageClearVec_readReady_24 = ~needWAR | readChannel_24_ready_0;
  assign stageClearVec_WaitReadQueue_24_enq_valid = stageClearVec_reqQueue_24_deq_valid & stageClearVec_readReady_24;
  assign stageClearVec_reqQueue_24_deq_ready = stageClearVec_WaitReadQueue_24_enq_ready & stageClearVec_readReady_24;
  wire        readChannel_24_valid_0 = stageClearVec_reqQueue_24_deq_valid & needWAR & stageClearVec_WaitReadQueue_24_enq_ready;
  wire [4:0]  readChannel_24_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_24_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_24_bits_offset_0 = stageClearVec_reqQueue_24_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_24 = ~needWAR | readResult_24_valid;
  wire [31:0] stageClearVec_WARData_24 = stageClearVec_WaitReadQueue_24_deq_bits_data & stageClearVec_WaitReadQueue_24_deq_bits_bitMask | readResult_24_bits & ~stageClearVec_WaitReadQueue_24_deq_bits_bitMask;
  wire        out_24_valid_0 = stageClearVec_WaitReadQueue_24_deq_valid & stageClearVec_readResultValid_24;
  assign stageClearVec_WaitReadQueue_24_deq_ready = out_24_ready_0 & stageClearVec_readResultValid_24;
  wire [31:0] out_24_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_24 : stageClearVec_WaitReadQueue_24_deq_bits_data;
  wire [3:0]  out_24_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_24_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_24;
  wire        _stageClearVec_T_72 = in_24_ready_0 & in_24_valid_0;
  wire [2:0]  stageClearVec_counterChange_24 = _stageClearVec_T_72 ? 3'h1 : 3'h7;
  wire        stageClearVec_24 = stageClearVec_counter_24 == 3'h0;
  wire        in_25_ready_0 = stageClearVec_reqQueue_25_enq_ready;
  wire        stageClearVec_reqQueue_25_deq_valid;
  assign stageClearVec_reqQueue_25_deq_valid = ~_stageClearVec_reqQueue_fifo_25_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_25_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_25_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_25_enq_bits_data = stageClearVec_reqQueue_25_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_25_mask;
  wire [31:0] stageClearVec_WaitReadQueue_25_enq_bits_bitMask = stageClearVec_reqQueue_25_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_25_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_25_enq_bits_mask = stageClearVec_reqQueue_25_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_25_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_25_enq_bits_groupCounter = stageClearVec_reqQueue_25_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_25_enq_bits_ffoByOther = stageClearVec_reqQueue_25_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_25 = {stageClearVec_reqQueue_25_enq_bits_groupCounter, stageClearVec_reqQueue_25_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_25 = {stageClearVec_reqQueue_25_enq_bits_data, stageClearVec_reqQueue_25_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_25 = {stageClearVec_reqQueue_dataIn_hi_hi_25, stageClearVec_reqQueue_25_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_25 = {stageClearVec_reqQueue_dataIn_hi_25, stageClearVec_reqQueue_dataIn_lo_25};
  assign stageClearVec_reqQueue_dataOut_25_ffoByOther = _stageClearVec_reqQueue_fifo_25_data_out[0];
  assign stageClearVec_reqQueue_dataOut_25_groupCounter = _stageClearVec_reqQueue_fifo_25_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_25_mask = _stageClearVec_reqQueue_fifo_25_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_25_bitMask = _stageClearVec_reqQueue_fifo_25_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_25_data = _stageClearVec_reqQueue_fifo_25_data_out[74:43];
  assign stageClearVec_reqQueue_25_deq_bits_data = stageClearVec_reqQueue_dataOut_25_data;
  assign stageClearVec_reqQueue_25_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_25_bitMask;
  assign stageClearVec_reqQueue_25_deq_bits_mask = stageClearVec_reqQueue_dataOut_25_mask;
  assign stageClearVec_reqQueue_25_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_25_groupCounter;
  assign stageClearVec_reqQueue_25_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_25_ffoByOther;
  assign stageClearVec_reqQueue_25_enq_ready = ~_stageClearVec_reqQueue_fifo_25_full;
  wire        stageClearVec_reqQueue_25_deq_ready;
  wire        stageClearVec_WaitReadQueue_25_deq_valid;
  assign stageClearVec_WaitReadQueue_25_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_25_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_25_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_25_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_25_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_25_groupCounter;
  wire [5:0]  out_25_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_25_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_25_ffoByOther;
  wire        out_25_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_25_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_25 = {stageClearVec_WaitReadQueue_25_enq_bits_groupCounter, stageClearVec_WaitReadQueue_25_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_25 = {stageClearVec_WaitReadQueue_25_enq_bits_data, stageClearVec_WaitReadQueue_25_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_25 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_25, stageClearVec_WaitReadQueue_25_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_25 = {stageClearVec_WaitReadQueue_dataIn_hi_25, stageClearVec_WaitReadQueue_dataIn_lo_25};
  assign stageClearVec_WaitReadQueue_dataOut_25_ffoByOther = _stageClearVec_WaitReadQueue_fifo_25_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_25_groupCounter = _stageClearVec_WaitReadQueue_fifo_25_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_25_mask = _stageClearVec_WaitReadQueue_fifo_25_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_25_bitMask = _stageClearVec_WaitReadQueue_fifo_25_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_25_data = _stageClearVec_WaitReadQueue_fifo_25_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_25_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_25_data;
  wire [31:0] stageClearVec_WaitReadQueue_25_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_25_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_25_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_25_mask;
  assign stageClearVec_WaitReadQueue_25_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_25_groupCounter;
  assign stageClearVec_WaitReadQueue_25_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_25_ffoByOther;
  wire        stageClearVec_WaitReadQueue_25_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_25_full;
  wire        stageClearVec_WaitReadQueue_25_enq_valid;
  wire        stageClearVec_WaitReadQueue_25_deq_ready;
  wire        stageClearVec_readReady_25 = ~needWAR | readChannel_25_ready_0;
  assign stageClearVec_WaitReadQueue_25_enq_valid = stageClearVec_reqQueue_25_deq_valid & stageClearVec_readReady_25;
  assign stageClearVec_reqQueue_25_deq_ready = stageClearVec_WaitReadQueue_25_enq_ready & stageClearVec_readReady_25;
  wire        readChannel_25_valid_0 = stageClearVec_reqQueue_25_deq_valid & needWAR & stageClearVec_WaitReadQueue_25_enq_ready;
  wire [4:0]  readChannel_25_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_25_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_25_bits_offset_0 = stageClearVec_reqQueue_25_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_25 = ~needWAR | readResult_25_valid;
  wire [31:0] stageClearVec_WARData_25 = stageClearVec_WaitReadQueue_25_deq_bits_data & stageClearVec_WaitReadQueue_25_deq_bits_bitMask | readResult_25_bits & ~stageClearVec_WaitReadQueue_25_deq_bits_bitMask;
  wire        out_25_valid_0 = stageClearVec_WaitReadQueue_25_deq_valid & stageClearVec_readResultValid_25;
  assign stageClearVec_WaitReadQueue_25_deq_ready = out_25_ready_0 & stageClearVec_readResultValid_25;
  wire [31:0] out_25_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_25 : stageClearVec_WaitReadQueue_25_deq_bits_data;
  wire [3:0]  out_25_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_25_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_25;
  wire        _stageClearVec_T_75 = in_25_ready_0 & in_25_valid_0;
  wire [2:0]  stageClearVec_counterChange_25 = _stageClearVec_T_75 ? 3'h1 : 3'h7;
  wire        stageClearVec_25 = stageClearVec_counter_25 == 3'h0;
  wire        in_26_ready_0 = stageClearVec_reqQueue_26_enq_ready;
  wire        stageClearVec_reqQueue_26_deq_valid;
  assign stageClearVec_reqQueue_26_deq_valid = ~_stageClearVec_reqQueue_fifo_26_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_26_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_26_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_26_enq_bits_data = stageClearVec_reqQueue_26_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_26_mask;
  wire [31:0] stageClearVec_WaitReadQueue_26_enq_bits_bitMask = stageClearVec_reqQueue_26_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_26_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_26_enq_bits_mask = stageClearVec_reqQueue_26_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_26_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_26_enq_bits_groupCounter = stageClearVec_reqQueue_26_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_26_enq_bits_ffoByOther = stageClearVec_reqQueue_26_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_26 = {stageClearVec_reqQueue_26_enq_bits_groupCounter, stageClearVec_reqQueue_26_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_26 = {stageClearVec_reqQueue_26_enq_bits_data, stageClearVec_reqQueue_26_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_26 = {stageClearVec_reqQueue_dataIn_hi_hi_26, stageClearVec_reqQueue_26_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_26 = {stageClearVec_reqQueue_dataIn_hi_26, stageClearVec_reqQueue_dataIn_lo_26};
  assign stageClearVec_reqQueue_dataOut_26_ffoByOther = _stageClearVec_reqQueue_fifo_26_data_out[0];
  assign stageClearVec_reqQueue_dataOut_26_groupCounter = _stageClearVec_reqQueue_fifo_26_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_26_mask = _stageClearVec_reqQueue_fifo_26_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_26_bitMask = _stageClearVec_reqQueue_fifo_26_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_26_data = _stageClearVec_reqQueue_fifo_26_data_out[74:43];
  assign stageClearVec_reqQueue_26_deq_bits_data = stageClearVec_reqQueue_dataOut_26_data;
  assign stageClearVec_reqQueue_26_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_26_bitMask;
  assign stageClearVec_reqQueue_26_deq_bits_mask = stageClearVec_reqQueue_dataOut_26_mask;
  assign stageClearVec_reqQueue_26_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_26_groupCounter;
  assign stageClearVec_reqQueue_26_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_26_ffoByOther;
  assign stageClearVec_reqQueue_26_enq_ready = ~_stageClearVec_reqQueue_fifo_26_full;
  wire        stageClearVec_reqQueue_26_deq_ready;
  wire        stageClearVec_WaitReadQueue_26_deq_valid;
  assign stageClearVec_WaitReadQueue_26_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_26_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_26_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_26_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_26_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_26_groupCounter;
  wire [5:0]  out_26_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_26_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_26_ffoByOther;
  wire        out_26_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_26_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_26 = {stageClearVec_WaitReadQueue_26_enq_bits_groupCounter, stageClearVec_WaitReadQueue_26_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_26 = {stageClearVec_WaitReadQueue_26_enq_bits_data, stageClearVec_WaitReadQueue_26_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_26 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_26, stageClearVec_WaitReadQueue_26_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_26 = {stageClearVec_WaitReadQueue_dataIn_hi_26, stageClearVec_WaitReadQueue_dataIn_lo_26};
  assign stageClearVec_WaitReadQueue_dataOut_26_ffoByOther = _stageClearVec_WaitReadQueue_fifo_26_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_26_groupCounter = _stageClearVec_WaitReadQueue_fifo_26_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_26_mask = _stageClearVec_WaitReadQueue_fifo_26_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_26_bitMask = _stageClearVec_WaitReadQueue_fifo_26_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_26_data = _stageClearVec_WaitReadQueue_fifo_26_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_26_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_26_data;
  wire [31:0] stageClearVec_WaitReadQueue_26_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_26_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_26_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_26_mask;
  assign stageClearVec_WaitReadQueue_26_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_26_groupCounter;
  assign stageClearVec_WaitReadQueue_26_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_26_ffoByOther;
  wire        stageClearVec_WaitReadQueue_26_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_26_full;
  wire        stageClearVec_WaitReadQueue_26_enq_valid;
  wire        stageClearVec_WaitReadQueue_26_deq_ready;
  wire        stageClearVec_readReady_26 = ~needWAR | readChannel_26_ready_0;
  assign stageClearVec_WaitReadQueue_26_enq_valid = stageClearVec_reqQueue_26_deq_valid & stageClearVec_readReady_26;
  assign stageClearVec_reqQueue_26_deq_ready = stageClearVec_WaitReadQueue_26_enq_ready & stageClearVec_readReady_26;
  wire        readChannel_26_valid_0 = stageClearVec_reqQueue_26_deq_valid & needWAR & stageClearVec_WaitReadQueue_26_enq_ready;
  wire [4:0]  readChannel_26_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_26_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_26_bits_offset_0 = stageClearVec_reqQueue_26_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_26 = ~needWAR | readResult_26_valid;
  wire [31:0] stageClearVec_WARData_26 = stageClearVec_WaitReadQueue_26_deq_bits_data & stageClearVec_WaitReadQueue_26_deq_bits_bitMask | readResult_26_bits & ~stageClearVec_WaitReadQueue_26_deq_bits_bitMask;
  wire        out_26_valid_0 = stageClearVec_WaitReadQueue_26_deq_valid & stageClearVec_readResultValid_26;
  assign stageClearVec_WaitReadQueue_26_deq_ready = out_26_ready_0 & stageClearVec_readResultValid_26;
  wire [31:0] out_26_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_26 : stageClearVec_WaitReadQueue_26_deq_bits_data;
  wire [3:0]  out_26_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_26_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_26;
  wire        _stageClearVec_T_78 = in_26_ready_0 & in_26_valid_0;
  wire [2:0]  stageClearVec_counterChange_26 = _stageClearVec_T_78 ? 3'h1 : 3'h7;
  wire        stageClearVec_26 = stageClearVec_counter_26 == 3'h0;
  wire        in_27_ready_0 = stageClearVec_reqQueue_27_enq_ready;
  wire        stageClearVec_reqQueue_27_deq_valid;
  assign stageClearVec_reqQueue_27_deq_valid = ~_stageClearVec_reqQueue_fifo_27_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_27_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_27_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_27_enq_bits_data = stageClearVec_reqQueue_27_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_27_mask;
  wire [31:0] stageClearVec_WaitReadQueue_27_enq_bits_bitMask = stageClearVec_reqQueue_27_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_27_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_27_enq_bits_mask = stageClearVec_reqQueue_27_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_27_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_27_enq_bits_groupCounter = stageClearVec_reqQueue_27_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_27_enq_bits_ffoByOther = stageClearVec_reqQueue_27_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_27 = {stageClearVec_reqQueue_27_enq_bits_groupCounter, stageClearVec_reqQueue_27_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_27 = {stageClearVec_reqQueue_27_enq_bits_data, stageClearVec_reqQueue_27_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_27 = {stageClearVec_reqQueue_dataIn_hi_hi_27, stageClearVec_reqQueue_27_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_27 = {stageClearVec_reqQueue_dataIn_hi_27, stageClearVec_reqQueue_dataIn_lo_27};
  assign stageClearVec_reqQueue_dataOut_27_ffoByOther = _stageClearVec_reqQueue_fifo_27_data_out[0];
  assign stageClearVec_reqQueue_dataOut_27_groupCounter = _stageClearVec_reqQueue_fifo_27_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_27_mask = _stageClearVec_reqQueue_fifo_27_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_27_bitMask = _stageClearVec_reqQueue_fifo_27_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_27_data = _stageClearVec_reqQueue_fifo_27_data_out[74:43];
  assign stageClearVec_reqQueue_27_deq_bits_data = stageClearVec_reqQueue_dataOut_27_data;
  assign stageClearVec_reqQueue_27_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_27_bitMask;
  assign stageClearVec_reqQueue_27_deq_bits_mask = stageClearVec_reqQueue_dataOut_27_mask;
  assign stageClearVec_reqQueue_27_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_27_groupCounter;
  assign stageClearVec_reqQueue_27_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_27_ffoByOther;
  assign stageClearVec_reqQueue_27_enq_ready = ~_stageClearVec_reqQueue_fifo_27_full;
  wire        stageClearVec_reqQueue_27_deq_ready;
  wire        stageClearVec_WaitReadQueue_27_deq_valid;
  assign stageClearVec_WaitReadQueue_27_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_27_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_27_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_27_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_27_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_27_groupCounter;
  wire [5:0]  out_27_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_27_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_27_ffoByOther;
  wire        out_27_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_27_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_27 = {stageClearVec_WaitReadQueue_27_enq_bits_groupCounter, stageClearVec_WaitReadQueue_27_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_27 = {stageClearVec_WaitReadQueue_27_enq_bits_data, stageClearVec_WaitReadQueue_27_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_27 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_27, stageClearVec_WaitReadQueue_27_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_27 = {stageClearVec_WaitReadQueue_dataIn_hi_27, stageClearVec_WaitReadQueue_dataIn_lo_27};
  assign stageClearVec_WaitReadQueue_dataOut_27_ffoByOther = _stageClearVec_WaitReadQueue_fifo_27_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_27_groupCounter = _stageClearVec_WaitReadQueue_fifo_27_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_27_mask = _stageClearVec_WaitReadQueue_fifo_27_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_27_bitMask = _stageClearVec_WaitReadQueue_fifo_27_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_27_data = _stageClearVec_WaitReadQueue_fifo_27_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_27_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_27_data;
  wire [31:0] stageClearVec_WaitReadQueue_27_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_27_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_27_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_27_mask;
  assign stageClearVec_WaitReadQueue_27_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_27_groupCounter;
  assign stageClearVec_WaitReadQueue_27_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_27_ffoByOther;
  wire        stageClearVec_WaitReadQueue_27_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_27_full;
  wire        stageClearVec_WaitReadQueue_27_enq_valid;
  wire        stageClearVec_WaitReadQueue_27_deq_ready;
  wire        stageClearVec_readReady_27 = ~needWAR | readChannel_27_ready_0;
  assign stageClearVec_WaitReadQueue_27_enq_valid = stageClearVec_reqQueue_27_deq_valid & stageClearVec_readReady_27;
  assign stageClearVec_reqQueue_27_deq_ready = stageClearVec_WaitReadQueue_27_enq_ready & stageClearVec_readReady_27;
  wire        readChannel_27_valid_0 = stageClearVec_reqQueue_27_deq_valid & needWAR & stageClearVec_WaitReadQueue_27_enq_ready;
  wire [4:0]  readChannel_27_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_27_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_27_bits_offset_0 = stageClearVec_reqQueue_27_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_27 = ~needWAR | readResult_27_valid;
  wire [31:0] stageClearVec_WARData_27 = stageClearVec_WaitReadQueue_27_deq_bits_data & stageClearVec_WaitReadQueue_27_deq_bits_bitMask | readResult_27_bits & ~stageClearVec_WaitReadQueue_27_deq_bits_bitMask;
  wire        out_27_valid_0 = stageClearVec_WaitReadQueue_27_deq_valid & stageClearVec_readResultValid_27;
  assign stageClearVec_WaitReadQueue_27_deq_ready = out_27_ready_0 & stageClearVec_readResultValid_27;
  wire [31:0] out_27_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_27 : stageClearVec_WaitReadQueue_27_deq_bits_data;
  wire [3:0]  out_27_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_27_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_27;
  wire        _stageClearVec_T_81 = in_27_ready_0 & in_27_valid_0;
  wire [2:0]  stageClearVec_counterChange_27 = _stageClearVec_T_81 ? 3'h1 : 3'h7;
  wire        stageClearVec_27 = stageClearVec_counter_27 == 3'h0;
  wire        in_28_ready_0 = stageClearVec_reqQueue_28_enq_ready;
  wire        stageClearVec_reqQueue_28_deq_valid;
  assign stageClearVec_reqQueue_28_deq_valid = ~_stageClearVec_reqQueue_fifo_28_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_28_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_28_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_28_enq_bits_data = stageClearVec_reqQueue_28_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_28_mask;
  wire [31:0] stageClearVec_WaitReadQueue_28_enq_bits_bitMask = stageClearVec_reqQueue_28_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_28_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_28_enq_bits_mask = stageClearVec_reqQueue_28_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_28_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_28_enq_bits_groupCounter = stageClearVec_reqQueue_28_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_28_enq_bits_ffoByOther = stageClearVec_reqQueue_28_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_28 = {stageClearVec_reqQueue_28_enq_bits_groupCounter, stageClearVec_reqQueue_28_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_28 = {stageClearVec_reqQueue_28_enq_bits_data, stageClearVec_reqQueue_28_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_28 = {stageClearVec_reqQueue_dataIn_hi_hi_28, stageClearVec_reqQueue_28_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_28 = {stageClearVec_reqQueue_dataIn_hi_28, stageClearVec_reqQueue_dataIn_lo_28};
  assign stageClearVec_reqQueue_dataOut_28_ffoByOther = _stageClearVec_reqQueue_fifo_28_data_out[0];
  assign stageClearVec_reqQueue_dataOut_28_groupCounter = _stageClearVec_reqQueue_fifo_28_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_28_mask = _stageClearVec_reqQueue_fifo_28_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_28_bitMask = _stageClearVec_reqQueue_fifo_28_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_28_data = _stageClearVec_reqQueue_fifo_28_data_out[74:43];
  assign stageClearVec_reqQueue_28_deq_bits_data = stageClearVec_reqQueue_dataOut_28_data;
  assign stageClearVec_reqQueue_28_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_28_bitMask;
  assign stageClearVec_reqQueue_28_deq_bits_mask = stageClearVec_reqQueue_dataOut_28_mask;
  assign stageClearVec_reqQueue_28_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_28_groupCounter;
  assign stageClearVec_reqQueue_28_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_28_ffoByOther;
  assign stageClearVec_reqQueue_28_enq_ready = ~_stageClearVec_reqQueue_fifo_28_full;
  wire        stageClearVec_reqQueue_28_deq_ready;
  wire        stageClearVec_WaitReadQueue_28_deq_valid;
  assign stageClearVec_WaitReadQueue_28_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_28_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_28_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_28_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_28_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_28_groupCounter;
  wire [5:0]  out_28_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_28_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_28_ffoByOther;
  wire        out_28_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_28_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_28 = {stageClearVec_WaitReadQueue_28_enq_bits_groupCounter, stageClearVec_WaitReadQueue_28_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_28 = {stageClearVec_WaitReadQueue_28_enq_bits_data, stageClearVec_WaitReadQueue_28_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_28 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_28, stageClearVec_WaitReadQueue_28_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_28 = {stageClearVec_WaitReadQueue_dataIn_hi_28, stageClearVec_WaitReadQueue_dataIn_lo_28};
  assign stageClearVec_WaitReadQueue_dataOut_28_ffoByOther = _stageClearVec_WaitReadQueue_fifo_28_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_28_groupCounter = _stageClearVec_WaitReadQueue_fifo_28_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_28_mask = _stageClearVec_WaitReadQueue_fifo_28_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_28_bitMask = _stageClearVec_WaitReadQueue_fifo_28_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_28_data = _stageClearVec_WaitReadQueue_fifo_28_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_28_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_28_data;
  wire [31:0] stageClearVec_WaitReadQueue_28_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_28_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_28_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_28_mask;
  assign stageClearVec_WaitReadQueue_28_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_28_groupCounter;
  assign stageClearVec_WaitReadQueue_28_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_28_ffoByOther;
  wire        stageClearVec_WaitReadQueue_28_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_28_full;
  wire        stageClearVec_WaitReadQueue_28_enq_valid;
  wire        stageClearVec_WaitReadQueue_28_deq_ready;
  wire        stageClearVec_readReady_28 = ~needWAR | readChannel_28_ready_0;
  assign stageClearVec_WaitReadQueue_28_enq_valid = stageClearVec_reqQueue_28_deq_valid & stageClearVec_readReady_28;
  assign stageClearVec_reqQueue_28_deq_ready = stageClearVec_WaitReadQueue_28_enq_ready & stageClearVec_readReady_28;
  wire        readChannel_28_valid_0 = stageClearVec_reqQueue_28_deq_valid & needWAR & stageClearVec_WaitReadQueue_28_enq_ready;
  wire [4:0]  readChannel_28_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_28_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_28_bits_offset_0 = stageClearVec_reqQueue_28_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_28 = ~needWAR | readResult_28_valid;
  wire [31:0] stageClearVec_WARData_28 = stageClearVec_WaitReadQueue_28_deq_bits_data & stageClearVec_WaitReadQueue_28_deq_bits_bitMask | readResult_28_bits & ~stageClearVec_WaitReadQueue_28_deq_bits_bitMask;
  wire        out_28_valid_0 = stageClearVec_WaitReadQueue_28_deq_valid & stageClearVec_readResultValid_28;
  assign stageClearVec_WaitReadQueue_28_deq_ready = out_28_ready_0 & stageClearVec_readResultValid_28;
  wire [31:0] out_28_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_28 : stageClearVec_WaitReadQueue_28_deq_bits_data;
  wire [3:0]  out_28_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_28_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_28;
  wire        _stageClearVec_T_84 = in_28_ready_0 & in_28_valid_0;
  wire [2:0]  stageClearVec_counterChange_28 = _stageClearVec_T_84 ? 3'h1 : 3'h7;
  wire        stageClearVec_28 = stageClearVec_counter_28 == 3'h0;
  wire        in_29_ready_0 = stageClearVec_reqQueue_29_enq_ready;
  wire        stageClearVec_reqQueue_29_deq_valid;
  assign stageClearVec_reqQueue_29_deq_valid = ~_stageClearVec_reqQueue_fifo_29_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_29_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_29_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_29_enq_bits_data = stageClearVec_reqQueue_29_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_29_mask;
  wire [31:0] stageClearVec_WaitReadQueue_29_enq_bits_bitMask = stageClearVec_reqQueue_29_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_29_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_29_enq_bits_mask = stageClearVec_reqQueue_29_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_29_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_29_enq_bits_groupCounter = stageClearVec_reqQueue_29_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_29_enq_bits_ffoByOther = stageClearVec_reqQueue_29_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_29 = {stageClearVec_reqQueue_29_enq_bits_groupCounter, stageClearVec_reqQueue_29_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_29 = {stageClearVec_reqQueue_29_enq_bits_data, stageClearVec_reqQueue_29_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_29 = {stageClearVec_reqQueue_dataIn_hi_hi_29, stageClearVec_reqQueue_29_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_29 = {stageClearVec_reqQueue_dataIn_hi_29, stageClearVec_reqQueue_dataIn_lo_29};
  assign stageClearVec_reqQueue_dataOut_29_ffoByOther = _stageClearVec_reqQueue_fifo_29_data_out[0];
  assign stageClearVec_reqQueue_dataOut_29_groupCounter = _stageClearVec_reqQueue_fifo_29_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_29_mask = _stageClearVec_reqQueue_fifo_29_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_29_bitMask = _stageClearVec_reqQueue_fifo_29_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_29_data = _stageClearVec_reqQueue_fifo_29_data_out[74:43];
  assign stageClearVec_reqQueue_29_deq_bits_data = stageClearVec_reqQueue_dataOut_29_data;
  assign stageClearVec_reqQueue_29_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_29_bitMask;
  assign stageClearVec_reqQueue_29_deq_bits_mask = stageClearVec_reqQueue_dataOut_29_mask;
  assign stageClearVec_reqQueue_29_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_29_groupCounter;
  assign stageClearVec_reqQueue_29_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_29_ffoByOther;
  assign stageClearVec_reqQueue_29_enq_ready = ~_stageClearVec_reqQueue_fifo_29_full;
  wire        stageClearVec_reqQueue_29_deq_ready;
  wire        stageClearVec_WaitReadQueue_29_deq_valid;
  assign stageClearVec_WaitReadQueue_29_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_29_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_29_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_29_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_29_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_29_groupCounter;
  wire [5:0]  out_29_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_29_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_29_ffoByOther;
  wire        out_29_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_29_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_29 = {stageClearVec_WaitReadQueue_29_enq_bits_groupCounter, stageClearVec_WaitReadQueue_29_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_29 = {stageClearVec_WaitReadQueue_29_enq_bits_data, stageClearVec_WaitReadQueue_29_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_29 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_29, stageClearVec_WaitReadQueue_29_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_29 = {stageClearVec_WaitReadQueue_dataIn_hi_29, stageClearVec_WaitReadQueue_dataIn_lo_29};
  assign stageClearVec_WaitReadQueue_dataOut_29_ffoByOther = _stageClearVec_WaitReadQueue_fifo_29_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_29_groupCounter = _stageClearVec_WaitReadQueue_fifo_29_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_29_mask = _stageClearVec_WaitReadQueue_fifo_29_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_29_bitMask = _stageClearVec_WaitReadQueue_fifo_29_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_29_data = _stageClearVec_WaitReadQueue_fifo_29_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_29_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_29_data;
  wire [31:0] stageClearVec_WaitReadQueue_29_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_29_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_29_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_29_mask;
  assign stageClearVec_WaitReadQueue_29_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_29_groupCounter;
  assign stageClearVec_WaitReadQueue_29_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_29_ffoByOther;
  wire        stageClearVec_WaitReadQueue_29_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_29_full;
  wire        stageClearVec_WaitReadQueue_29_enq_valid;
  wire        stageClearVec_WaitReadQueue_29_deq_ready;
  wire        stageClearVec_readReady_29 = ~needWAR | readChannel_29_ready_0;
  assign stageClearVec_WaitReadQueue_29_enq_valid = stageClearVec_reqQueue_29_deq_valid & stageClearVec_readReady_29;
  assign stageClearVec_reqQueue_29_deq_ready = stageClearVec_WaitReadQueue_29_enq_ready & stageClearVec_readReady_29;
  wire        readChannel_29_valid_0 = stageClearVec_reqQueue_29_deq_valid & needWAR & stageClearVec_WaitReadQueue_29_enq_ready;
  wire [4:0]  readChannel_29_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_29_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_29_bits_offset_0 = stageClearVec_reqQueue_29_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_29 = ~needWAR | readResult_29_valid;
  wire [31:0] stageClearVec_WARData_29 = stageClearVec_WaitReadQueue_29_deq_bits_data & stageClearVec_WaitReadQueue_29_deq_bits_bitMask | readResult_29_bits & ~stageClearVec_WaitReadQueue_29_deq_bits_bitMask;
  wire        out_29_valid_0 = stageClearVec_WaitReadQueue_29_deq_valid & stageClearVec_readResultValid_29;
  assign stageClearVec_WaitReadQueue_29_deq_ready = out_29_ready_0 & stageClearVec_readResultValid_29;
  wire [31:0] out_29_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_29 : stageClearVec_WaitReadQueue_29_deq_bits_data;
  wire [3:0]  out_29_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_29_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_29;
  wire        _stageClearVec_T_87 = in_29_ready_0 & in_29_valid_0;
  wire [2:0]  stageClearVec_counterChange_29 = _stageClearVec_T_87 ? 3'h1 : 3'h7;
  wire        stageClearVec_29 = stageClearVec_counter_29 == 3'h0;
  wire        in_30_ready_0 = stageClearVec_reqQueue_30_enq_ready;
  wire        stageClearVec_reqQueue_30_deq_valid;
  assign stageClearVec_reqQueue_30_deq_valid = ~_stageClearVec_reqQueue_fifo_30_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_30_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_30_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_30_enq_bits_data = stageClearVec_reqQueue_30_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_30_mask;
  wire [31:0] stageClearVec_WaitReadQueue_30_enq_bits_bitMask = stageClearVec_reqQueue_30_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_30_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_30_enq_bits_mask = stageClearVec_reqQueue_30_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_30_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_30_enq_bits_groupCounter = stageClearVec_reqQueue_30_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_30_enq_bits_ffoByOther = stageClearVec_reqQueue_30_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_30 = {stageClearVec_reqQueue_30_enq_bits_groupCounter, stageClearVec_reqQueue_30_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_30 = {stageClearVec_reqQueue_30_enq_bits_data, stageClearVec_reqQueue_30_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_30 = {stageClearVec_reqQueue_dataIn_hi_hi_30, stageClearVec_reqQueue_30_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_30 = {stageClearVec_reqQueue_dataIn_hi_30, stageClearVec_reqQueue_dataIn_lo_30};
  assign stageClearVec_reqQueue_dataOut_30_ffoByOther = _stageClearVec_reqQueue_fifo_30_data_out[0];
  assign stageClearVec_reqQueue_dataOut_30_groupCounter = _stageClearVec_reqQueue_fifo_30_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_30_mask = _stageClearVec_reqQueue_fifo_30_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_30_bitMask = _stageClearVec_reqQueue_fifo_30_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_30_data = _stageClearVec_reqQueue_fifo_30_data_out[74:43];
  assign stageClearVec_reqQueue_30_deq_bits_data = stageClearVec_reqQueue_dataOut_30_data;
  assign stageClearVec_reqQueue_30_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_30_bitMask;
  assign stageClearVec_reqQueue_30_deq_bits_mask = stageClearVec_reqQueue_dataOut_30_mask;
  assign stageClearVec_reqQueue_30_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_30_groupCounter;
  assign stageClearVec_reqQueue_30_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_30_ffoByOther;
  assign stageClearVec_reqQueue_30_enq_ready = ~_stageClearVec_reqQueue_fifo_30_full;
  wire        stageClearVec_reqQueue_30_deq_ready;
  wire        stageClearVec_WaitReadQueue_30_deq_valid;
  assign stageClearVec_WaitReadQueue_30_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_30_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_30_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_30_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_30_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_30_groupCounter;
  wire [5:0]  out_30_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_30_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_30_ffoByOther;
  wire        out_30_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_30_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_30 = {stageClearVec_WaitReadQueue_30_enq_bits_groupCounter, stageClearVec_WaitReadQueue_30_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_30 = {stageClearVec_WaitReadQueue_30_enq_bits_data, stageClearVec_WaitReadQueue_30_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_30 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_30, stageClearVec_WaitReadQueue_30_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_30 = {stageClearVec_WaitReadQueue_dataIn_hi_30, stageClearVec_WaitReadQueue_dataIn_lo_30};
  assign stageClearVec_WaitReadQueue_dataOut_30_ffoByOther = _stageClearVec_WaitReadQueue_fifo_30_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_30_groupCounter = _stageClearVec_WaitReadQueue_fifo_30_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_30_mask = _stageClearVec_WaitReadQueue_fifo_30_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_30_bitMask = _stageClearVec_WaitReadQueue_fifo_30_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_30_data = _stageClearVec_WaitReadQueue_fifo_30_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_30_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_30_data;
  wire [31:0] stageClearVec_WaitReadQueue_30_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_30_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_30_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_30_mask;
  assign stageClearVec_WaitReadQueue_30_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_30_groupCounter;
  assign stageClearVec_WaitReadQueue_30_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_30_ffoByOther;
  wire        stageClearVec_WaitReadQueue_30_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_30_full;
  wire        stageClearVec_WaitReadQueue_30_enq_valid;
  wire        stageClearVec_WaitReadQueue_30_deq_ready;
  wire        stageClearVec_readReady_30 = ~needWAR | readChannel_30_ready_0;
  assign stageClearVec_WaitReadQueue_30_enq_valid = stageClearVec_reqQueue_30_deq_valid & stageClearVec_readReady_30;
  assign stageClearVec_reqQueue_30_deq_ready = stageClearVec_WaitReadQueue_30_enq_ready & stageClearVec_readReady_30;
  wire        readChannel_30_valid_0 = stageClearVec_reqQueue_30_deq_valid & needWAR & stageClearVec_WaitReadQueue_30_enq_ready;
  wire [4:0]  readChannel_30_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_30_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_30_bits_offset_0 = stageClearVec_reqQueue_30_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_30 = ~needWAR | readResult_30_valid;
  wire [31:0] stageClearVec_WARData_30 = stageClearVec_WaitReadQueue_30_deq_bits_data & stageClearVec_WaitReadQueue_30_deq_bits_bitMask | readResult_30_bits & ~stageClearVec_WaitReadQueue_30_deq_bits_bitMask;
  wire        out_30_valid_0 = stageClearVec_WaitReadQueue_30_deq_valid & stageClearVec_readResultValid_30;
  assign stageClearVec_WaitReadQueue_30_deq_ready = out_30_ready_0 & stageClearVec_readResultValid_30;
  wire [31:0] out_30_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_30 : stageClearVec_WaitReadQueue_30_deq_bits_data;
  wire [3:0]  out_30_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_30_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_30;
  wire        _stageClearVec_T_90 = in_30_ready_0 & in_30_valid_0;
  wire [2:0]  stageClearVec_counterChange_30 = _stageClearVec_T_90 ? 3'h1 : 3'h7;
  wire        stageClearVec_30 = stageClearVec_counter_30 == 3'h0;
  wire        in_31_ready_0 = stageClearVec_reqQueue_31_enq_ready;
  wire        stageClearVec_reqQueue_31_deq_valid;
  assign stageClearVec_reqQueue_31_deq_valid = ~_stageClearVec_reqQueue_fifo_31_empty;
  wire [31:0] stageClearVec_reqQueue_dataOut_31_data;
  wire [31:0] stageClearVec_reqQueue_dataOut_31_bitMask;
  wire [31:0] stageClearVec_WaitReadQueue_31_enq_bits_data = stageClearVec_reqQueue_31_deq_bits_data;
  wire [3:0]  stageClearVec_reqQueue_dataOut_31_mask;
  wire [31:0] stageClearVec_WaitReadQueue_31_enq_bits_bitMask = stageClearVec_reqQueue_31_deq_bits_bitMask;
  wire [5:0]  stageClearVec_reqQueue_dataOut_31_groupCounter;
  wire [3:0]  stageClearVec_WaitReadQueue_31_enq_bits_mask = stageClearVec_reqQueue_31_deq_bits_mask;
  wire        stageClearVec_reqQueue_dataOut_31_ffoByOther;
  wire [5:0]  stageClearVec_WaitReadQueue_31_enq_bits_groupCounter = stageClearVec_reqQueue_31_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_31_enq_bits_ffoByOther = stageClearVec_reqQueue_31_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_reqQueue_dataIn_lo_31 = {stageClearVec_reqQueue_31_enq_bits_groupCounter, stageClearVec_reqQueue_31_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_reqQueue_dataIn_hi_hi_31 = {stageClearVec_reqQueue_31_enq_bits_data, stageClearVec_reqQueue_31_enq_bits_bitMask};
  wire [67:0] stageClearVec_reqQueue_dataIn_hi_31 = {stageClearVec_reqQueue_dataIn_hi_hi_31, stageClearVec_reqQueue_31_enq_bits_mask};
  wire [74:0] stageClearVec_reqQueue_dataIn_31 = {stageClearVec_reqQueue_dataIn_hi_31, stageClearVec_reqQueue_dataIn_lo_31};
  assign stageClearVec_reqQueue_dataOut_31_ffoByOther = _stageClearVec_reqQueue_fifo_31_data_out[0];
  assign stageClearVec_reqQueue_dataOut_31_groupCounter = _stageClearVec_reqQueue_fifo_31_data_out[6:1];
  assign stageClearVec_reqQueue_dataOut_31_mask = _stageClearVec_reqQueue_fifo_31_data_out[10:7];
  assign stageClearVec_reqQueue_dataOut_31_bitMask = _stageClearVec_reqQueue_fifo_31_data_out[42:11];
  assign stageClearVec_reqQueue_dataOut_31_data = _stageClearVec_reqQueue_fifo_31_data_out[74:43];
  assign stageClearVec_reqQueue_31_deq_bits_data = stageClearVec_reqQueue_dataOut_31_data;
  assign stageClearVec_reqQueue_31_deq_bits_bitMask = stageClearVec_reqQueue_dataOut_31_bitMask;
  assign stageClearVec_reqQueue_31_deq_bits_mask = stageClearVec_reqQueue_dataOut_31_mask;
  assign stageClearVec_reqQueue_31_deq_bits_groupCounter = stageClearVec_reqQueue_dataOut_31_groupCounter;
  assign stageClearVec_reqQueue_31_deq_bits_ffoByOther = stageClearVec_reqQueue_dataOut_31_ffoByOther;
  assign stageClearVec_reqQueue_31_enq_ready = ~_stageClearVec_reqQueue_fifo_31_full;
  wire        stageClearVec_reqQueue_31_deq_ready;
  wire        stageClearVec_WaitReadQueue_31_deq_valid;
  assign stageClearVec_WaitReadQueue_31_deq_valid = ~_stageClearVec_WaitReadQueue_fifo_31_empty;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_31_data;
  wire [31:0] stageClearVec_WaitReadQueue_dataOut_31_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_dataOut_31_mask;
  wire [5:0]  stageClearVec_WaitReadQueue_dataOut_31_groupCounter;
  wire [5:0]  out_31_bits_writeData_groupCounter_0 = stageClearVec_WaitReadQueue_31_deq_bits_groupCounter;
  wire        stageClearVec_WaitReadQueue_dataOut_31_ffoByOther;
  wire        out_31_bits_ffoByOther_0 = stageClearVec_WaitReadQueue_31_deq_bits_ffoByOther;
  wire [6:0]  stageClearVec_WaitReadQueue_dataIn_lo_31 = {stageClearVec_WaitReadQueue_31_enq_bits_groupCounter, stageClearVec_WaitReadQueue_31_enq_bits_ffoByOther};
  wire [63:0] stageClearVec_WaitReadQueue_dataIn_hi_hi_31 = {stageClearVec_WaitReadQueue_31_enq_bits_data, stageClearVec_WaitReadQueue_31_enq_bits_bitMask};
  wire [67:0] stageClearVec_WaitReadQueue_dataIn_hi_31 = {stageClearVec_WaitReadQueue_dataIn_hi_hi_31, stageClearVec_WaitReadQueue_31_enq_bits_mask};
  wire [74:0] stageClearVec_WaitReadQueue_dataIn_31 = {stageClearVec_WaitReadQueue_dataIn_hi_31, stageClearVec_WaitReadQueue_dataIn_lo_31};
  assign stageClearVec_WaitReadQueue_dataOut_31_ffoByOther = _stageClearVec_WaitReadQueue_fifo_31_data_out[0];
  assign stageClearVec_WaitReadQueue_dataOut_31_groupCounter = _stageClearVec_WaitReadQueue_fifo_31_data_out[6:1];
  assign stageClearVec_WaitReadQueue_dataOut_31_mask = _stageClearVec_WaitReadQueue_fifo_31_data_out[10:7];
  assign stageClearVec_WaitReadQueue_dataOut_31_bitMask = _stageClearVec_WaitReadQueue_fifo_31_data_out[42:11];
  assign stageClearVec_WaitReadQueue_dataOut_31_data = _stageClearVec_WaitReadQueue_fifo_31_data_out[74:43];
  wire [31:0] stageClearVec_WaitReadQueue_31_deq_bits_data = stageClearVec_WaitReadQueue_dataOut_31_data;
  wire [31:0] stageClearVec_WaitReadQueue_31_deq_bits_bitMask = stageClearVec_WaitReadQueue_dataOut_31_bitMask;
  wire [3:0]  stageClearVec_WaitReadQueue_31_deq_bits_mask = stageClearVec_WaitReadQueue_dataOut_31_mask;
  assign stageClearVec_WaitReadQueue_31_deq_bits_groupCounter = stageClearVec_WaitReadQueue_dataOut_31_groupCounter;
  assign stageClearVec_WaitReadQueue_31_deq_bits_ffoByOther = stageClearVec_WaitReadQueue_dataOut_31_ffoByOther;
  wire        stageClearVec_WaitReadQueue_31_enq_ready = ~_stageClearVec_WaitReadQueue_fifo_31_full;
  wire        stageClearVec_WaitReadQueue_31_enq_valid;
  wire        stageClearVec_WaitReadQueue_31_deq_ready;
  wire        stageClearVec_readReady_31 = ~needWAR | readChannel_31_ready_0;
  assign stageClearVec_WaitReadQueue_31_enq_valid = stageClearVec_reqQueue_31_deq_valid & stageClearVec_readReady_31;
  assign stageClearVec_reqQueue_31_deq_ready = stageClearVec_WaitReadQueue_31_enq_ready & stageClearVec_readReady_31;
  wire        readChannel_31_valid_0 = stageClearVec_reqQueue_31_deq_valid & needWAR & stageClearVec_WaitReadQueue_31_enq_ready;
  wire [4:0]  readChannel_31_bits_vs_0 = vd + {1'h0, stageClearVec_reqQueue_31_deq_bits_groupCounter[5:2]};
  wire [1:0]  readChannel_31_bits_offset_0 = stageClearVec_reqQueue_31_deq_bits_groupCounter[1:0];
  wire        stageClearVec_readResultValid_31 = ~needWAR | readResult_31_valid;
  wire [31:0] stageClearVec_WARData_31 = stageClearVec_WaitReadQueue_31_deq_bits_data & stageClearVec_WaitReadQueue_31_deq_bits_bitMask | readResult_31_bits & ~stageClearVec_WaitReadQueue_31_deq_bits_bitMask;
  wire        out_31_valid_0 = stageClearVec_WaitReadQueue_31_deq_valid & stageClearVec_readResultValid_31;
  assign stageClearVec_WaitReadQueue_31_deq_ready = out_31_ready_0 & stageClearVec_readResultValid_31;
  wire [31:0] out_31_bits_writeData_data_0 = needWAR ? stageClearVec_WARData_31 : stageClearVec_WaitReadQueue_31_deq_bits_data;
  wire [3:0]  out_31_bits_writeData_mask_0 = needWAR ? 4'hF : stageClearVec_WaitReadQueue_31_deq_bits_mask;
  reg  [2:0]  stageClearVec_counter_31;
  wire        _stageClearVec_T_93 = in_31_ready_0 & in_31_valid_0;
  wire [2:0]  stageClearVec_counterChange_31 = _stageClearVec_T_93 ? 3'h1 : 3'h7;
  wire        stageClearVec_31 = stageClearVec_counter_31 == 3'h0;
  always @(posedge clock) begin
    if (reset) begin
      stageClearVec_counter <= 3'h0;
      stageClearVec_counter_1 <= 3'h0;
      stageClearVec_counter_2 <= 3'h0;
      stageClearVec_counter_3 <= 3'h0;
      stageClearVec_counter_4 <= 3'h0;
      stageClearVec_counter_5 <= 3'h0;
      stageClearVec_counter_6 <= 3'h0;
      stageClearVec_counter_7 <= 3'h0;
      stageClearVec_counter_8 <= 3'h0;
      stageClearVec_counter_9 <= 3'h0;
      stageClearVec_counter_10 <= 3'h0;
      stageClearVec_counter_11 <= 3'h0;
      stageClearVec_counter_12 <= 3'h0;
      stageClearVec_counter_13 <= 3'h0;
      stageClearVec_counter_14 <= 3'h0;
      stageClearVec_counter_15 <= 3'h0;
      stageClearVec_counter_16 <= 3'h0;
      stageClearVec_counter_17 <= 3'h0;
      stageClearVec_counter_18 <= 3'h0;
      stageClearVec_counter_19 <= 3'h0;
      stageClearVec_counter_20 <= 3'h0;
      stageClearVec_counter_21 <= 3'h0;
      stageClearVec_counter_22 <= 3'h0;
      stageClearVec_counter_23 <= 3'h0;
      stageClearVec_counter_24 <= 3'h0;
      stageClearVec_counter_25 <= 3'h0;
      stageClearVec_counter_26 <= 3'h0;
      stageClearVec_counter_27 <= 3'h0;
      stageClearVec_counter_28 <= 3'h0;
      stageClearVec_counter_29 <= 3'h0;
      stageClearVec_counter_30 <= 3'h0;
      stageClearVec_counter_31 <= 3'h0;
    end
    else begin
      if (_stageClearVec_T ^ out_0_ready_0 & out_0_valid_0)
        stageClearVec_counter <= stageClearVec_counter + stageClearVec_counterChange;
      if (_stageClearVec_T_3 ^ out_1_ready_0 & out_1_valid_0)
        stageClearVec_counter_1 <= stageClearVec_counter_1 + stageClearVec_counterChange_1;
      if (_stageClearVec_T_6 ^ out_2_ready_0 & out_2_valid_0)
        stageClearVec_counter_2 <= stageClearVec_counter_2 + stageClearVec_counterChange_2;
      if (_stageClearVec_T_9 ^ out_3_ready_0 & out_3_valid_0)
        stageClearVec_counter_3 <= stageClearVec_counter_3 + stageClearVec_counterChange_3;
      if (_stageClearVec_T_12 ^ out_4_ready_0 & out_4_valid_0)
        stageClearVec_counter_4 <= stageClearVec_counter_4 + stageClearVec_counterChange_4;
      if (_stageClearVec_T_15 ^ out_5_ready_0 & out_5_valid_0)
        stageClearVec_counter_5 <= stageClearVec_counter_5 + stageClearVec_counterChange_5;
      if (_stageClearVec_T_18 ^ out_6_ready_0 & out_6_valid_0)
        stageClearVec_counter_6 <= stageClearVec_counter_6 + stageClearVec_counterChange_6;
      if (_stageClearVec_T_21 ^ out_7_ready_0 & out_7_valid_0)
        stageClearVec_counter_7 <= stageClearVec_counter_7 + stageClearVec_counterChange_7;
      if (_stageClearVec_T_24 ^ out_8_ready_0 & out_8_valid_0)
        stageClearVec_counter_8 <= stageClearVec_counter_8 + stageClearVec_counterChange_8;
      if (_stageClearVec_T_27 ^ out_9_ready_0 & out_9_valid_0)
        stageClearVec_counter_9 <= stageClearVec_counter_9 + stageClearVec_counterChange_9;
      if (_stageClearVec_T_30 ^ out_10_ready_0 & out_10_valid_0)
        stageClearVec_counter_10 <= stageClearVec_counter_10 + stageClearVec_counterChange_10;
      if (_stageClearVec_T_33 ^ out_11_ready_0 & out_11_valid_0)
        stageClearVec_counter_11 <= stageClearVec_counter_11 + stageClearVec_counterChange_11;
      if (_stageClearVec_T_36 ^ out_12_ready_0 & out_12_valid_0)
        stageClearVec_counter_12 <= stageClearVec_counter_12 + stageClearVec_counterChange_12;
      if (_stageClearVec_T_39 ^ out_13_ready_0 & out_13_valid_0)
        stageClearVec_counter_13 <= stageClearVec_counter_13 + stageClearVec_counterChange_13;
      if (_stageClearVec_T_42 ^ out_14_ready_0 & out_14_valid_0)
        stageClearVec_counter_14 <= stageClearVec_counter_14 + stageClearVec_counterChange_14;
      if (_stageClearVec_T_45 ^ out_15_ready_0 & out_15_valid_0)
        stageClearVec_counter_15 <= stageClearVec_counter_15 + stageClearVec_counterChange_15;
      if (_stageClearVec_T_48 ^ out_16_ready_0 & out_16_valid_0)
        stageClearVec_counter_16 <= stageClearVec_counter_16 + stageClearVec_counterChange_16;
      if (_stageClearVec_T_51 ^ out_17_ready_0 & out_17_valid_0)
        stageClearVec_counter_17 <= stageClearVec_counter_17 + stageClearVec_counterChange_17;
      if (_stageClearVec_T_54 ^ out_18_ready_0 & out_18_valid_0)
        stageClearVec_counter_18 <= stageClearVec_counter_18 + stageClearVec_counterChange_18;
      if (_stageClearVec_T_57 ^ out_19_ready_0 & out_19_valid_0)
        stageClearVec_counter_19 <= stageClearVec_counter_19 + stageClearVec_counterChange_19;
      if (_stageClearVec_T_60 ^ out_20_ready_0 & out_20_valid_0)
        stageClearVec_counter_20 <= stageClearVec_counter_20 + stageClearVec_counterChange_20;
      if (_stageClearVec_T_63 ^ out_21_ready_0 & out_21_valid_0)
        stageClearVec_counter_21 <= stageClearVec_counter_21 + stageClearVec_counterChange_21;
      if (_stageClearVec_T_66 ^ out_22_ready_0 & out_22_valid_0)
        stageClearVec_counter_22 <= stageClearVec_counter_22 + stageClearVec_counterChange_22;
      if (_stageClearVec_T_69 ^ out_23_ready_0 & out_23_valid_0)
        stageClearVec_counter_23 <= stageClearVec_counter_23 + stageClearVec_counterChange_23;
      if (_stageClearVec_T_72 ^ out_24_ready_0 & out_24_valid_0)
        stageClearVec_counter_24 <= stageClearVec_counter_24 + stageClearVec_counterChange_24;
      if (_stageClearVec_T_75 ^ out_25_ready_0 & out_25_valid_0)
        stageClearVec_counter_25 <= stageClearVec_counter_25 + stageClearVec_counterChange_25;
      if (_stageClearVec_T_78 ^ out_26_ready_0 & out_26_valid_0)
        stageClearVec_counter_26 <= stageClearVec_counter_26 + stageClearVec_counterChange_26;
      if (_stageClearVec_T_81 ^ out_27_ready_0 & out_27_valid_0)
        stageClearVec_counter_27 <= stageClearVec_counter_27 + stageClearVec_counterChange_27;
      if (_stageClearVec_T_84 ^ out_28_ready_0 & out_28_valid_0)
        stageClearVec_counter_28 <= stageClearVec_counter_28 + stageClearVec_counterChange_28;
      if (_stageClearVec_T_87 ^ out_29_ready_0 & out_29_valid_0)
        stageClearVec_counter_29 <= stageClearVec_counter_29 + stageClearVec_counterChange_29;
      if (_stageClearVec_T_90 ^ out_30_ready_0 & out_30_valid_0)
        stageClearVec_counter_30 <= stageClearVec_counter_30 + stageClearVec_counterChange_30;
      if (_stageClearVec_T_93 ^ out_31_ready_0 & out_31_valid_0)
        stageClearVec_counter_31 <= stageClearVec_counter_31 + stageClearVec_counterChange_31;
    end
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:2];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [1:0] i = 2'h0; i < 2'h3; i += 2'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        stageClearVec_counter = _RANDOM[2'h0][2:0];
        stageClearVec_counter_1 = _RANDOM[2'h0][5:3];
        stageClearVec_counter_2 = _RANDOM[2'h0][8:6];
        stageClearVec_counter_3 = _RANDOM[2'h0][11:9];
        stageClearVec_counter_4 = _RANDOM[2'h0][14:12];
        stageClearVec_counter_5 = _RANDOM[2'h0][17:15];
        stageClearVec_counter_6 = _RANDOM[2'h0][20:18];
        stageClearVec_counter_7 = _RANDOM[2'h0][23:21];
        stageClearVec_counter_8 = _RANDOM[2'h0][26:24];
        stageClearVec_counter_9 = _RANDOM[2'h0][29:27];
        stageClearVec_counter_10 = {_RANDOM[2'h0][31:30], _RANDOM[2'h1][0]};
        stageClearVec_counter_11 = _RANDOM[2'h1][3:1];
        stageClearVec_counter_12 = _RANDOM[2'h1][6:4];
        stageClearVec_counter_13 = _RANDOM[2'h1][9:7];
        stageClearVec_counter_14 = _RANDOM[2'h1][12:10];
        stageClearVec_counter_15 = _RANDOM[2'h1][15:13];
        stageClearVec_counter_16 = _RANDOM[2'h1][18:16];
        stageClearVec_counter_17 = _RANDOM[2'h1][21:19];
        stageClearVec_counter_18 = _RANDOM[2'h1][24:22];
        stageClearVec_counter_19 = _RANDOM[2'h1][27:25];
        stageClearVec_counter_20 = _RANDOM[2'h1][30:28];
        stageClearVec_counter_21 = {_RANDOM[2'h1][31], _RANDOM[2'h2][1:0]};
        stageClearVec_counter_22 = _RANDOM[2'h2][4:2];
        stageClearVec_counter_23 = _RANDOM[2'h2][7:5];
        stageClearVec_counter_24 = _RANDOM[2'h2][10:8];
        stageClearVec_counter_25 = _RANDOM[2'h2][13:11];
        stageClearVec_counter_26 = _RANDOM[2'h2][16:14];
        stageClearVec_counter_27 = _RANDOM[2'h2][19:17];
        stageClearVec_counter_28 = _RANDOM[2'h2][22:20];
        stageClearVec_counter_29 = _RANDOM[2'h2][25:23];
        stageClearVec_counter_30 = _RANDOM[2'h2][28:26];
        stageClearVec_counter_31 = _RANDOM[2'h2][31:29];
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  wire        stageClearVec_reqQueue_empty;
  assign stageClearVec_reqQueue_empty = _stageClearVec_reqQueue_fifo_empty;
  wire        stageClearVec_reqQueue_full;
  assign stageClearVec_reqQueue_full = _stageClearVec_reqQueue_fifo_full;
  wire        stageClearVec_WaitReadQueue_empty;
  assign stageClearVec_WaitReadQueue_empty = _stageClearVec_WaitReadQueue_fifo_empty;
  wire        stageClearVec_WaitReadQueue_full;
  assign stageClearVec_WaitReadQueue_full = _stageClearVec_WaitReadQueue_fifo_full;
  wire        stageClearVec_reqQueue_1_empty;
  assign stageClearVec_reqQueue_1_empty = _stageClearVec_reqQueue_fifo_1_empty;
  wire        stageClearVec_reqQueue_1_full;
  assign stageClearVec_reqQueue_1_full = _stageClearVec_reqQueue_fifo_1_full;
  wire        stageClearVec_WaitReadQueue_1_empty;
  assign stageClearVec_WaitReadQueue_1_empty = _stageClearVec_WaitReadQueue_fifo_1_empty;
  wire        stageClearVec_WaitReadQueue_1_full;
  assign stageClearVec_WaitReadQueue_1_full = _stageClearVec_WaitReadQueue_fifo_1_full;
  wire        stageClearVec_reqQueue_2_empty;
  assign stageClearVec_reqQueue_2_empty = _stageClearVec_reqQueue_fifo_2_empty;
  wire        stageClearVec_reqQueue_2_full;
  assign stageClearVec_reqQueue_2_full = _stageClearVec_reqQueue_fifo_2_full;
  wire        stageClearVec_WaitReadQueue_2_empty;
  assign stageClearVec_WaitReadQueue_2_empty = _stageClearVec_WaitReadQueue_fifo_2_empty;
  wire        stageClearVec_WaitReadQueue_2_full;
  assign stageClearVec_WaitReadQueue_2_full = _stageClearVec_WaitReadQueue_fifo_2_full;
  wire        stageClearVec_reqQueue_3_empty;
  assign stageClearVec_reqQueue_3_empty = _stageClearVec_reqQueue_fifo_3_empty;
  wire        stageClearVec_reqQueue_3_full;
  assign stageClearVec_reqQueue_3_full = _stageClearVec_reqQueue_fifo_3_full;
  wire        stageClearVec_WaitReadQueue_3_empty;
  assign stageClearVec_WaitReadQueue_3_empty = _stageClearVec_WaitReadQueue_fifo_3_empty;
  wire        stageClearVec_WaitReadQueue_3_full;
  assign stageClearVec_WaitReadQueue_3_full = _stageClearVec_WaitReadQueue_fifo_3_full;
  wire        stageClearVec_reqQueue_4_empty;
  assign stageClearVec_reqQueue_4_empty = _stageClearVec_reqQueue_fifo_4_empty;
  wire        stageClearVec_reqQueue_4_full;
  assign stageClearVec_reqQueue_4_full = _stageClearVec_reqQueue_fifo_4_full;
  wire        stageClearVec_WaitReadQueue_4_empty;
  assign stageClearVec_WaitReadQueue_4_empty = _stageClearVec_WaitReadQueue_fifo_4_empty;
  wire        stageClearVec_WaitReadQueue_4_full;
  assign stageClearVec_WaitReadQueue_4_full = _stageClearVec_WaitReadQueue_fifo_4_full;
  wire        stageClearVec_reqQueue_5_empty;
  assign stageClearVec_reqQueue_5_empty = _stageClearVec_reqQueue_fifo_5_empty;
  wire        stageClearVec_reqQueue_5_full;
  assign stageClearVec_reqQueue_5_full = _stageClearVec_reqQueue_fifo_5_full;
  wire        stageClearVec_WaitReadQueue_5_empty;
  assign stageClearVec_WaitReadQueue_5_empty = _stageClearVec_WaitReadQueue_fifo_5_empty;
  wire        stageClearVec_WaitReadQueue_5_full;
  assign stageClearVec_WaitReadQueue_5_full = _stageClearVec_WaitReadQueue_fifo_5_full;
  wire        stageClearVec_reqQueue_6_empty;
  assign stageClearVec_reqQueue_6_empty = _stageClearVec_reqQueue_fifo_6_empty;
  wire        stageClearVec_reqQueue_6_full;
  assign stageClearVec_reqQueue_6_full = _stageClearVec_reqQueue_fifo_6_full;
  wire        stageClearVec_WaitReadQueue_6_empty;
  assign stageClearVec_WaitReadQueue_6_empty = _stageClearVec_WaitReadQueue_fifo_6_empty;
  wire        stageClearVec_WaitReadQueue_6_full;
  assign stageClearVec_WaitReadQueue_6_full = _stageClearVec_WaitReadQueue_fifo_6_full;
  wire        stageClearVec_reqQueue_7_empty;
  assign stageClearVec_reqQueue_7_empty = _stageClearVec_reqQueue_fifo_7_empty;
  wire        stageClearVec_reqQueue_7_full;
  assign stageClearVec_reqQueue_7_full = _stageClearVec_reqQueue_fifo_7_full;
  wire        stageClearVec_WaitReadQueue_7_empty;
  assign stageClearVec_WaitReadQueue_7_empty = _stageClearVec_WaitReadQueue_fifo_7_empty;
  wire        stageClearVec_WaitReadQueue_7_full;
  assign stageClearVec_WaitReadQueue_7_full = _stageClearVec_WaitReadQueue_fifo_7_full;
  wire        stageClearVec_reqQueue_8_empty;
  assign stageClearVec_reqQueue_8_empty = _stageClearVec_reqQueue_fifo_8_empty;
  wire        stageClearVec_reqQueue_8_full;
  assign stageClearVec_reqQueue_8_full = _stageClearVec_reqQueue_fifo_8_full;
  wire        stageClearVec_WaitReadQueue_8_empty;
  assign stageClearVec_WaitReadQueue_8_empty = _stageClearVec_WaitReadQueue_fifo_8_empty;
  wire        stageClearVec_WaitReadQueue_8_full;
  assign stageClearVec_WaitReadQueue_8_full = _stageClearVec_WaitReadQueue_fifo_8_full;
  wire        stageClearVec_reqQueue_9_empty;
  assign stageClearVec_reqQueue_9_empty = _stageClearVec_reqQueue_fifo_9_empty;
  wire        stageClearVec_reqQueue_9_full;
  assign stageClearVec_reqQueue_9_full = _stageClearVec_reqQueue_fifo_9_full;
  wire        stageClearVec_WaitReadQueue_9_empty;
  assign stageClearVec_WaitReadQueue_9_empty = _stageClearVec_WaitReadQueue_fifo_9_empty;
  wire        stageClearVec_WaitReadQueue_9_full;
  assign stageClearVec_WaitReadQueue_9_full = _stageClearVec_WaitReadQueue_fifo_9_full;
  wire        stageClearVec_reqQueue_10_empty;
  assign stageClearVec_reqQueue_10_empty = _stageClearVec_reqQueue_fifo_10_empty;
  wire        stageClearVec_reqQueue_10_full;
  assign stageClearVec_reqQueue_10_full = _stageClearVec_reqQueue_fifo_10_full;
  wire        stageClearVec_WaitReadQueue_10_empty;
  assign stageClearVec_WaitReadQueue_10_empty = _stageClearVec_WaitReadQueue_fifo_10_empty;
  wire        stageClearVec_WaitReadQueue_10_full;
  assign stageClearVec_WaitReadQueue_10_full = _stageClearVec_WaitReadQueue_fifo_10_full;
  wire        stageClearVec_reqQueue_11_empty;
  assign stageClearVec_reqQueue_11_empty = _stageClearVec_reqQueue_fifo_11_empty;
  wire        stageClearVec_reqQueue_11_full;
  assign stageClearVec_reqQueue_11_full = _stageClearVec_reqQueue_fifo_11_full;
  wire        stageClearVec_WaitReadQueue_11_empty;
  assign stageClearVec_WaitReadQueue_11_empty = _stageClearVec_WaitReadQueue_fifo_11_empty;
  wire        stageClearVec_WaitReadQueue_11_full;
  assign stageClearVec_WaitReadQueue_11_full = _stageClearVec_WaitReadQueue_fifo_11_full;
  wire        stageClearVec_reqQueue_12_empty;
  assign stageClearVec_reqQueue_12_empty = _stageClearVec_reqQueue_fifo_12_empty;
  wire        stageClearVec_reqQueue_12_full;
  assign stageClearVec_reqQueue_12_full = _stageClearVec_reqQueue_fifo_12_full;
  wire        stageClearVec_WaitReadQueue_12_empty;
  assign stageClearVec_WaitReadQueue_12_empty = _stageClearVec_WaitReadQueue_fifo_12_empty;
  wire        stageClearVec_WaitReadQueue_12_full;
  assign stageClearVec_WaitReadQueue_12_full = _stageClearVec_WaitReadQueue_fifo_12_full;
  wire        stageClearVec_reqQueue_13_empty;
  assign stageClearVec_reqQueue_13_empty = _stageClearVec_reqQueue_fifo_13_empty;
  wire        stageClearVec_reqQueue_13_full;
  assign stageClearVec_reqQueue_13_full = _stageClearVec_reqQueue_fifo_13_full;
  wire        stageClearVec_WaitReadQueue_13_empty;
  assign stageClearVec_WaitReadQueue_13_empty = _stageClearVec_WaitReadQueue_fifo_13_empty;
  wire        stageClearVec_WaitReadQueue_13_full;
  assign stageClearVec_WaitReadQueue_13_full = _stageClearVec_WaitReadQueue_fifo_13_full;
  wire        stageClearVec_reqQueue_14_empty;
  assign stageClearVec_reqQueue_14_empty = _stageClearVec_reqQueue_fifo_14_empty;
  wire        stageClearVec_reqQueue_14_full;
  assign stageClearVec_reqQueue_14_full = _stageClearVec_reqQueue_fifo_14_full;
  wire        stageClearVec_WaitReadQueue_14_empty;
  assign stageClearVec_WaitReadQueue_14_empty = _stageClearVec_WaitReadQueue_fifo_14_empty;
  wire        stageClearVec_WaitReadQueue_14_full;
  assign stageClearVec_WaitReadQueue_14_full = _stageClearVec_WaitReadQueue_fifo_14_full;
  wire        stageClearVec_reqQueue_15_empty;
  assign stageClearVec_reqQueue_15_empty = _stageClearVec_reqQueue_fifo_15_empty;
  wire        stageClearVec_reqQueue_15_full;
  assign stageClearVec_reqQueue_15_full = _stageClearVec_reqQueue_fifo_15_full;
  wire        stageClearVec_WaitReadQueue_15_empty;
  assign stageClearVec_WaitReadQueue_15_empty = _stageClearVec_WaitReadQueue_fifo_15_empty;
  wire        stageClearVec_WaitReadQueue_15_full;
  assign stageClearVec_WaitReadQueue_15_full = _stageClearVec_WaitReadQueue_fifo_15_full;
  wire        stageClearVec_reqQueue_16_empty;
  assign stageClearVec_reqQueue_16_empty = _stageClearVec_reqQueue_fifo_16_empty;
  wire        stageClearVec_reqQueue_16_full;
  assign stageClearVec_reqQueue_16_full = _stageClearVec_reqQueue_fifo_16_full;
  wire        stageClearVec_WaitReadQueue_16_empty;
  assign stageClearVec_WaitReadQueue_16_empty = _stageClearVec_WaitReadQueue_fifo_16_empty;
  wire        stageClearVec_WaitReadQueue_16_full;
  assign stageClearVec_WaitReadQueue_16_full = _stageClearVec_WaitReadQueue_fifo_16_full;
  wire        stageClearVec_reqQueue_17_empty;
  assign stageClearVec_reqQueue_17_empty = _stageClearVec_reqQueue_fifo_17_empty;
  wire        stageClearVec_reqQueue_17_full;
  assign stageClearVec_reqQueue_17_full = _stageClearVec_reqQueue_fifo_17_full;
  wire        stageClearVec_WaitReadQueue_17_empty;
  assign stageClearVec_WaitReadQueue_17_empty = _stageClearVec_WaitReadQueue_fifo_17_empty;
  wire        stageClearVec_WaitReadQueue_17_full;
  assign stageClearVec_WaitReadQueue_17_full = _stageClearVec_WaitReadQueue_fifo_17_full;
  wire        stageClearVec_reqQueue_18_empty;
  assign stageClearVec_reqQueue_18_empty = _stageClearVec_reqQueue_fifo_18_empty;
  wire        stageClearVec_reqQueue_18_full;
  assign stageClearVec_reqQueue_18_full = _stageClearVec_reqQueue_fifo_18_full;
  wire        stageClearVec_WaitReadQueue_18_empty;
  assign stageClearVec_WaitReadQueue_18_empty = _stageClearVec_WaitReadQueue_fifo_18_empty;
  wire        stageClearVec_WaitReadQueue_18_full;
  assign stageClearVec_WaitReadQueue_18_full = _stageClearVec_WaitReadQueue_fifo_18_full;
  wire        stageClearVec_reqQueue_19_empty;
  assign stageClearVec_reqQueue_19_empty = _stageClearVec_reqQueue_fifo_19_empty;
  wire        stageClearVec_reqQueue_19_full;
  assign stageClearVec_reqQueue_19_full = _stageClearVec_reqQueue_fifo_19_full;
  wire        stageClearVec_WaitReadQueue_19_empty;
  assign stageClearVec_WaitReadQueue_19_empty = _stageClearVec_WaitReadQueue_fifo_19_empty;
  wire        stageClearVec_WaitReadQueue_19_full;
  assign stageClearVec_WaitReadQueue_19_full = _stageClearVec_WaitReadQueue_fifo_19_full;
  wire        stageClearVec_reqQueue_20_empty;
  assign stageClearVec_reqQueue_20_empty = _stageClearVec_reqQueue_fifo_20_empty;
  wire        stageClearVec_reqQueue_20_full;
  assign stageClearVec_reqQueue_20_full = _stageClearVec_reqQueue_fifo_20_full;
  wire        stageClearVec_WaitReadQueue_20_empty;
  assign stageClearVec_WaitReadQueue_20_empty = _stageClearVec_WaitReadQueue_fifo_20_empty;
  wire        stageClearVec_WaitReadQueue_20_full;
  assign stageClearVec_WaitReadQueue_20_full = _stageClearVec_WaitReadQueue_fifo_20_full;
  wire        stageClearVec_reqQueue_21_empty;
  assign stageClearVec_reqQueue_21_empty = _stageClearVec_reqQueue_fifo_21_empty;
  wire        stageClearVec_reqQueue_21_full;
  assign stageClearVec_reqQueue_21_full = _stageClearVec_reqQueue_fifo_21_full;
  wire        stageClearVec_WaitReadQueue_21_empty;
  assign stageClearVec_WaitReadQueue_21_empty = _stageClearVec_WaitReadQueue_fifo_21_empty;
  wire        stageClearVec_WaitReadQueue_21_full;
  assign stageClearVec_WaitReadQueue_21_full = _stageClearVec_WaitReadQueue_fifo_21_full;
  wire        stageClearVec_reqQueue_22_empty;
  assign stageClearVec_reqQueue_22_empty = _stageClearVec_reqQueue_fifo_22_empty;
  wire        stageClearVec_reqQueue_22_full;
  assign stageClearVec_reqQueue_22_full = _stageClearVec_reqQueue_fifo_22_full;
  wire        stageClearVec_WaitReadQueue_22_empty;
  assign stageClearVec_WaitReadQueue_22_empty = _stageClearVec_WaitReadQueue_fifo_22_empty;
  wire        stageClearVec_WaitReadQueue_22_full;
  assign stageClearVec_WaitReadQueue_22_full = _stageClearVec_WaitReadQueue_fifo_22_full;
  wire        stageClearVec_reqQueue_23_empty;
  assign stageClearVec_reqQueue_23_empty = _stageClearVec_reqQueue_fifo_23_empty;
  wire        stageClearVec_reqQueue_23_full;
  assign stageClearVec_reqQueue_23_full = _stageClearVec_reqQueue_fifo_23_full;
  wire        stageClearVec_WaitReadQueue_23_empty;
  assign stageClearVec_WaitReadQueue_23_empty = _stageClearVec_WaitReadQueue_fifo_23_empty;
  wire        stageClearVec_WaitReadQueue_23_full;
  assign stageClearVec_WaitReadQueue_23_full = _stageClearVec_WaitReadQueue_fifo_23_full;
  wire        stageClearVec_reqQueue_24_empty;
  assign stageClearVec_reqQueue_24_empty = _stageClearVec_reqQueue_fifo_24_empty;
  wire        stageClearVec_reqQueue_24_full;
  assign stageClearVec_reqQueue_24_full = _stageClearVec_reqQueue_fifo_24_full;
  wire        stageClearVec_WaitReadQueue_24_empty;
  assign stageClearVec_WaitReadQueue_24_empty = _stageClearVec_WaitReadQueue_fifo_24_empty;
  wire        stageClearVec_WaitReadQueue_24_full;
  assign stageClearVec_WaitReadQueue_24_full = _stageClearVec_WaitReadQueue_fifo_24_full;
  wire        stageClearVec_reqQueue_25_empty;
  assign stageClearVec_reqQueue_25_empty = _stageClearVec_reqQueue_fifo_25_empty;
  wire        stageClearVec_reqQueue_25_full;
  assign stageClearVec_reqQueue_25_full = _stageClearVec_reqQueue_fifo_25_full;
  wire        stageClearVec_WaitReadQueue_25_empty;
  assign stageClearVec_WaitReadQueue_25_empty = _stageClearVec_WaitReadQueue_fifo_25_empty;
  wire        stageClearVec_WaitReadQueue_25_full;
  assign stageClearVec_WaitReadQueue_25_full = _stageClearVec_WaitReadQueue_fifo_25_full;
  wire        stageClearVec_reqQueue_26_empty;
  assign stageClearVec_reqQueue_26_empty = _stageClearVec_reqQueue_fifo_26_empty;
  wire        stageClearVec_reqQueue_26_full;
  assign stageClearVec_reqQueue_26_full = _stageClearVec_reqQueue_fifo_26_full;
  wire        stageClearVec_WaitReadQueue_26_empty;
  assign stageClearVec_WaitReadQueue_26_empty = _stageClearVec_WaitReadQueue_fifo_26_empty;
  wire        stageClearVec_WaitReadQueue_26_full;
  assign stageClearVec_WaitReadQueue_26_full = _stageClearVec_WaitReadQueue_fifo_26_full;
  wire        stageClearVec_reqQueue_27_empty;
  assign stageClearVec_reqQueue_27_empty = _stageClearVec_reqQueue_fifo_27_empty;
  wire        stageClearVec_reqQueue_27_full;
  assign stageClearVec_reqQueue_27_full = _stageClearVec_reqQueue_fifo_27_full;
  wire        stageClearVec_WaitReadQueue_27_empty;
  assign stageClearVec_WaitReadQueue_27_empty = _stageClearVec_WaitReadQueue_fifo_27_empty;
  wire        stageClearVec_WaitReadQueue_27_full;
  assign stageClearVec_WaitReadQueue_27_full = _stageClearVec_WaitReadQueue_fifo_27_full;
  wire        stageClearVec_reqQueue_28_empty;
  assign stageClearVec_reqQueue_28_empty = _stageClearVec_reqQueue_fifo_28_empty;
  wire        stageClearVec_reqQueue_28_full;
  assign stageClearVec_reqQueue_28_full = _stageClearVec_reqQueue_fifo_28_full;
  wire        stageClearVec_WaitReadQueue_28_empty;
  assign stageClearVec_WaitReadQueue_28_empty = _stageClearVec_WaitReadQueue_fifo_28_empty;
  wire        stageClearVec_WaitReadQueue_28_full;
  assign stageClearVec_WaitReadQueue_28_full = _stageClearVec_WaitReadQueue_fifo_28_full;
  wire        stageClearVec_reqQueue_29_empty;
  assign stageClearVec_reqQueue_29_empty = _stageClearVec_reqQueue_fifo_29_empty;
  wire        stageClearVec_reqQueue_29_full;
  assign stageClearVec_reqQueue_29_full = _stageClearVec_reqQueue_fifo_29_full;
  wire        stageClearVec_WaitReadQueue_29_empty;
  assign stageClearVec_WaitReadQueue_29_empty = _stageClearVec_WaitReadQueue_fifo_29_empty;
  wire        stageClearVec_WaitReadQueue_29_full;
  assign stageClearVec_WaitReadQueue_29_full = _stageClearVec_WaitReadQueue_fifo_29_full;
  wire        stageClearVec_reqQueue_30_empty;
  assign stageClearVec_reqQueue_30_empty = _stageClearVec_reqQueue_fifo_30_empty;
  wire        stageClearVec_reqQueue_30_full;
  assign stageClearVec_reqQueue_30_full = _stageClearVec_reqQueue_fifo_30_full;
  wire        stageClearVec_WaitReadQueue_30_empty;
  assign stageClearVec_WaitReadQueue_30_empty = _stageClearVec_WaitReadQueue_fifo_30_empty;
  wire        stageClearVec_WaitReadQueue_30_full;
  assign stageClearVec_WaitReadQueue_30_full = _stageClearVec_WaitReadQueue_fifo_30_full;
  wire        stageClearVec_reqQueue_31_empty;
  assign stageClearVec_reqQueue_31_empty = _stageClearVec_reqQueue_fifo_31_empty;
  wire        stageClearVec_reqQueue_31_full;
  assign stageClearVec_reqQueue_31_full = _stageClearVec_reqQueue_fifo_31_full;
  wire        stageClearVec_WaitReadQueue_31_empty;
  assign stageClearVec_WaitReadQueue_31_empty = _stageClearVec_WaitReadQueue_fifo_31_empty;
  wire        stageClearVec_WaitReadQueue_31_full;
  assign stageClearVec_WaitReadQueue_31_full = _stageClearVec_WaitReadQueue_fifo_31_full;
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_enq_ready & stageClearVec_reqQueue_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_deq_ready & ~_stageClearVec_reqQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn),
    .empty        (_stageClearVec_reqQueue_fifo_empty),
    .almost_empty (stageClearVec_reqQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_full),
    .error        (_stageClearVec_reqQueue_fifo_error),
    .data_out     (_stageClearVec_reqQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_enq_ready & stageClearVec_WaitReadQueue_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn),
    .empty        (_stageClearVec_WaitReadQueue_fifo_empty),
    .almost_empty (stageClearVec_WaitReadQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_1_enq_ready & stageClearVec_reqQueue_1_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_1_deq_ready & ~_stageClearVec_reqQueue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_1),
    .empty        (_stageClearVec_reqQueue_fifo_1_empty),
    .almost_empty (stageClearVec_reqQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_1_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_1_full),
    .error        (_stageClearVec_reqQueue_fifo_1_error),
    .data_out     (_stageClearVec_reqQueue_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_1_enq_ready & stageClearVec_WaitReadQueue_1_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_1_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_1),
    .empty        (_stageClearVec_WaitReadQueue_fifo_1_empty),
    .almost_empty (stageClearVec_WaitReadQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_1_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_1_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_1_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_2_enq_ready & stageClearVec_reqQueue_2_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_2_deq_ready & ~_stageClearVec_reqQueue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_2),
    .empty        (_stageClearVec_reqQueue_fifo_2_empty),
    .almost_empty (stageClearVec_reqQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_2_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_2_full),
    .error        (_stageClearVec_reqQueue_fifo_2_error),
    .data_out     (_stageClearVec_reqQueue_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_2_enq_ready & stageClearVec_WaitReadQueue_2_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_2_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_2),
    .empty        (_stageClearVec_WaitReadQueue_fifo_2_empty),
    .almost_empty (stageClearVec_WaitReadQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_2_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_2_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_2_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_3_enq_ready & stageClearVec_reqQueue_3_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_3_deq_ready & ~_stageClearVec_reqQueue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_3),
    .empty        (_stageClearVec_reqQueue_fifo_3_empty),
    .almost_empty (stageClearVec_reqQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_3_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_3_full),
    .error        (_stageClearVec_reqQueue_fifo_3_error),
    .data_out     (_stageClearVec_reqQueue_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_3_enq_ready & stageClearVec_WaitReadQueue_3_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_3_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_3),
    .empty        (_stageClearVec_WaitReadQueue_fifo_3_empty),
    .almost_empty (stageClearVec_WaitReadQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_3_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_3_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_3_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_4_enq_ready & stageClearVec_reqQueue_4_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_4_deq_ready & ~_stageClearVec_reqQueue_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_4),
    .empty        (_stageClearVec_reqQueue_fifo_4_empty),
    .almost_empty (stageClearVec_reqQueue_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_4_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_4_full),
    .error        (_stageClearVec_reqQueue_fifo_4_error),
    .data_out     (_stageClearVec_reqQueue_fifo_4_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_4_enq_ready & stageClearVec_WaitReadQueue_4_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_4_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_4),
    .empty        (_stageClearVec_WaitReadQueue_fifo_4_empty),
    .almost_empty (stageClearVec_WaitReadQueue_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_4_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_4_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_4_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_4_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_5_enq_ready & stageClearVec_reqQueue_5_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_5_deq_ready & ~_stageClearVec_reqQueue_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_5),
    .empty        (_stageClearVec_reqQueue_fifo_5_empty),
    .almost_empty (stageClearVec_reqQueue_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_5_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_5_full),
    .error        (_stageClearVec_reqQueue_fifo_5_error),
    .data_out     (_stageClearVec_reqQueue_fifo_5_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_5_enq_ready & stageClearVec_WaitReadQueue_5_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_5_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_5),
    .empty        (_stageClearVec_WaitReadQueue_fifo_5_empty),
    .almost_empty (stageClearVec_WaitReadQueue_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_5_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_5_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_5_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_5_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_6_enq_ready & stageClearVec_reqQueue_6_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_6_deq_ready & ~_stageClearVec_reqQueue_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_6),
    .empty        (_stageClearVec_reqQueue_fifo_6_empty),
    .almost_empty (stageClearVec_reqQueue_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_6_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_6_full),
    .error        (_stageClearVec_reqQueue_fifo_6_error),
    .data_out     (_stageClearVec_reqQueue_fifo_6_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_6_enq_ready & stageClearVec_WaitReadQueue_6_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_6_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_6),
    .empty        (_stageClearVec_WaitReadQueue_fifo_6_empty),
    .almost_empty (stageClearVec_WaitReadQueue_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_6_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_6_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_6_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_6_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_7_enq_ready & stageClearVec_reqQueue_7_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_7_deq_ready & ~_stageClearVec_reqQueue_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_7),
    .empty        (_stageClearVec_reqQueue_fifo_7_empty),
    .almost_empty (stageClearVec_reqQueue_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_7_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_7_full),
    .error        (_stageClearVec_reqQueue_fifo_7_error),
    .data_out     (_stageClearVec_reqQueue_fifo_7_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_7_enq_ready & stageClearVec_WaitReadQueue_7_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_7_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_7),
    .empty        (_stageClearVec_WaitReadQueue_fifo_7_empty),
    .almost_empty (stageClearVec_WaitReadQueue_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_7_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_7_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_7_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_7_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_8 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_8_enq_ready & stageClearVec_reqQueue_8_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_8_deq_ready & ~_stageClearVec_reqQueue_fifo_8_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_8),
    .empty        (_stageClearVec_reqQueue_fifo_8_empty),
    .almost_empty (stageClearVec_reqQueue_8_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_8_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_8_full),
    .error        (_stageClearVec_reqQueue_fifo_8_error),
    .data_out     (_stageClearVec_reqQueue_fifo_8_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_8 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_8_enq_ready & stageClearVec_WaitReadQueue_8_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_8_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_8_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_8),
    .empty        (_stageClearVec_WaitReadQueue_fifo_8_empty),
    .almost_empty (stageClearVec_WaitReadQueue_8_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_8_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_8_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_8_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_8_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_9 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_9_enq_ready & stageClearVec_reqQueue_9_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_9_deq_ready & ~_stageClearVec_reqQueue_fifo_9_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_9),
    .empty        (_stageClearVec_reqQueue_fifo_9_empty),
    .almost_empty (stageClearVec_reqQueue_9_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_9_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_9_full),
    .error        (_stageClearVec_reqQueue_fifo_9_error),
    .data_out     (_stageClearVec_reqQueue_fifo_9_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_9 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_9_enq_ready & stageClearVec_WaitReadQueue_9_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_9_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_9_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_9),
    .empty        (_stageClearVec_WaitReadQueue_fifo_9_empty),
    .almost_empty (stageClearVec_WaitReadQueue_9_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_9_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_9_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_9_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_9_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_10 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_10_enq_ready & stageClearVec_reqQueue_10_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_10_deq_ready & ~_stageClearVec_reqQueue_fifo_10_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_10),
    .empty        (_stageClearVec_reqQueue_fifo_10_empty),
    .almost_empty (stageClearVec_reqQueue_10_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_10_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_10_full),
    .error        (_stageClearVec_reqQueue_fifo_10_error),
    .data_out     (_stageClearVec_reqQueue_fifo_10_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_10 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_10_enq_ready & stageClearVec_WaitReadQueue_10_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_10_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_10_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_10),
    .empty        (_stageClearVec_WaitReadQueue_fifo_10_empty),
    .almost_empty (stageClearVec_WaitReadQueue_10_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_10_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_10_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_10_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_10_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_11 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_11_enq_ready & stageClearVec_reqQueue_11_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_11_deq_ready & ~_stageClearVec_reqQueue_fifo_11_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_11),
    .empty        (_stageClearVec_reqQueue_fifo_11_empty),
    .almost_empty (stageClearVec_reqQueue_11_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_11_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_11_full),
    .error        (_stageClearVec_reqQueue_fifo_11_error),
    .data_out     (_stageClearVec_reqQueue_fifo_11_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_11 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_11_enq_ready & stageClearVec_WaitReadQueue_11_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_11_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_11_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_11),
    .empty        (_stageClearVec_WaitReadQueue_fifo_11_empty),
    .almost_empty (stageClearVec_WaitReadQueue_11_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_11_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_11_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_11_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_11_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_12 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_12_enq_ready & stageClearVec_reqQueue_12_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_12_deq_ready & ~_stageClearVec_reqQueue_fifo_12_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_12),
    .empty        (_stageClearVec_reqQueue_fifo_12_empty),
    .almost_empty (stageClearVec_reqQueue_12_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_12_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_12_full),
    .error        (_stageClearVec_reqQueue_fifo_12_error),
    .data_out     (_stageClearVec_reqQueue_fifo_12_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_12 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_12_enq_ready & stageClearVec_WaitReadQueue_12_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_12_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_12_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_12),
    .empty        (_stageClearVec_WaitReadQueue_fifo_12_empty),
    .almost_empty (stageClearVec_WaitReadQueue_12_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_12_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_12_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_12_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_12_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_13 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_13_enq_ready & stageClearVec_reqQueue_13_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_13_deq_ready & ~_stageClearVec_reqQueue_fifo_13_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_13),
    .empty        (_stageClearVec_reqQueue_fifo_13_empty),
    .almost_empty (stageClearVec_reqQueue_13_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_13_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_13_full),
    .error        (_stageClearVec_reqQueue_fifo_13_error),
    .data_out     (_stageClearVec_reqQueue_fifo_13_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_13 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_13_enq_ready & stageClearVec_WaitReadQueue_13_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_13_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_13_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_13),
    .empty        (_stageClearVec_WaitReadQueue_fifo_13_empty),
    .almost_empty (stageClearVec_WaitReadQueue_13_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_13_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_13_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_13_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_13_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_14 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_14_enq_ready & stageClearVec_reqQueue_14_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_14_deq_ready & ~_stageClearVec_reqQueue_fifo_14_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_14),
    .empty        (_stageClearVec_reqQueue_fifo_14_empty),
    .almost_empty (stageClearVec_reqQueue_14_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_14_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_14_full),
    .error        (_stageClearVec_reqQueue_fifo_14_error),
    .data_out     (_stageClearVec_reqQueue_fifo_14_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_14 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_14_enq_ready & stageClearVec_WaitReadQueue_14_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_14_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_14_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_14),
    .empty        (_stageClearVec_WaitReadQueue_fifo_14_empty),
    .almost_empty (stageClearVec_WaitReadQueue_14_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_14_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_14_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_14_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_14_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_15 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_15_enq_ready & stageClearVec_reqQueue_15_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_15_deq_ready & ~_stageClearVec_reqQueue_fifo_15_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_15),
    .empty        (_stageClearVec_reqQueue_fifo_15_empty),
    .almost_empty (stageClearVec_reqQueue_15_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_15_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_15_full),
    .error        (_stageClearVec_reqQueue_fifo_15_error),
    .data_out     (_stageClearVec_reqQueue_fifo_15_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_15 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_15_enq_ready & stageClearVec_WaitReadQueue_15_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_15_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_15_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_15),
    .empty        (_stageClearVec_WaitReadQueue_fifo_15_empty),
    .almost_empty (stageClearVec_WaitReadQueue_15_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_15_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_15_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_15_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_15_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_16 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_16_enq_ready & stageClearVec_reqQueue_16_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_16_deq_ready & ~_stageClearVec_reqQueue_fifo_16_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_16),
    .empty        (_stageClearVec_reqQueue_fifo_16_empty),
    .almost_empty (stageClearVec_reqQueue_16_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_16_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_16_full),
    .error        (_stageClearVec_reqQueue_fifo_16_error),
    .data_out     (_stageClearVec_reqQueue_fifo_16_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_16 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_16_enq_ready & stageClearVec_WaitReadQueue_16_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_16_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_16_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_16),
    .empty        (_stageClearVec_WaitReadQueue_fifo_16_empty),
    .almost_empty (stageClearVec_WaitReadQueue_16_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_16_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_16_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_16_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_16_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_17 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_17_enq_ready & stageClearVec_reqQueue_17_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_17_deq_ready & ~_stageClearVec_reqQueue_fifo_17_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_17),
    .empty        (_stageClearVec_reqQueue_fifo_17_empty),
    .almost_empty (stageClearVec_reqQueue_17_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_17_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_17_full),
    .error        (_stageClearVec_reqQueue_fifo_17_error),
    .data_out     (_stageClearVec_reqQueue_fifo_17_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_17 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_17_enq_ready & stageClearVec_WaitReadQueue_17_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_17_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_17_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_17),
    .empty        (_stageClearVec_WaitReadQueue_fifo_17_empty),
    .almost_empty (stageClearVec_WaitReadQueue_17_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_17_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_17_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_17_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_17_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_18 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_18_enq_ready & stageClearVec_reqQueue_18_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_18_deq_ready & ~_stageClearVec_reqQueue_fifo_18_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_18),
    .empty        (_stageClearVec_reqQueue_fifo_18_empty),
    .almost_empty (stageClearVec_reqQueue_18_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_18_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_18_full),
    .error        (_stageClearVec_reqQueue_fifo_18_error),
    .data_out     (_stageClearVec_reqQueue_fifo_18_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_18 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_18_enq_ready & stageClearVec_WaitReadQueue_18_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_18_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_18_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_18),
    .empty        (_stageClearVec_WaitReadQueue_fifo_18_empty),
    .almost_empty (stageClearVec_WaitReadQueue_18_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_18_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_18_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_18_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_18_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_19 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_19_enq_ready & stageClearVec_reqQueue_19_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_19_deq_ready & ~_stageClearVec_reqQueue_fifo_19_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_19),
    .empty        (_stageClearVec_reqQueue_fifo_19_empty),
    .almost_empty (stageClearVec_reqQueue_19_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_19_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_19_full),
    .error        (_stageClearVec_reqQueue_fifo_19_error),
    .data_out     (_stageClearVec_reqQueue_fifo_19_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_19 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_19_enq_ready & stageClearVec_WaitReadQueue_19_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_19_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_19_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_19),
    .empty        (_stageClearVec_WaitReadQueue_fifo_19_empty),
    .almost_empty (stageClearVec_WaitReadQueue_19_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_19_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_19_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_19_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_19_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_20 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_20_enq_ready & stageClearVec_reqQueue_20_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_20_deq_ready & ~_stageClearVec_reqQueue_fifo_20_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_20),
    .empty        (_stageClearVec_reqQueue_fifo_20_empty),
    .almost_empty (stageClearVec_reqQueue_20_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_20_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_20_full),
    .error        (_stageClearVec_reqQueue_fifo_20_error),
    .data_out     (_stageClearVec_reqQueue_fifo_20_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_20 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_20_enq_ready & stageClearVec_WaitReadQueue_20_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_20_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_20_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_20),
    .empty        (_stageClearVec_WaitReadQueue_fifo_20_empty),
    .almost_empty (stageClearVec_WaitReadQueue_20_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_20_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_20_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_20_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_20_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_21 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_21_enq_ready & stageClearVec_reqQueue_21_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_21_deq_ready & ~_stageClearVec_reqQueue_fifo_21_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_21),
    .empty        (_stageClearVec_reqQueue_fifo_21_empty),
    .almost_empty (stageClearVec_reqQueue_21_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_21_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_21_full),
    .error        (_stageClearVec_reqQueue_fifo_21_error),
    .data_out     (_stageClearVec_reqQueue_fifo_21_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_21 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_21_enq_ready & stageClearVec_WaitReadQueue_21_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_21_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_21_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_21),
    .empty        (_stageClearVec_WaitReadQueue_fifo_21_empty),
    .almost_empty (stageClearVec_WaitReadQueue_21_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_21_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_21_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_21_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_21_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_22 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_22_enq_ready & stageClearVec_reqQueue_22_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_22_deq_ready & ~_stageClearVec_reqQueue_fifo_22_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_22),
    .empty        (_stageClearVec_reqQueue_fifo_22_empty),
    .almost_empty (stageClearVec_reqQueue_22_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_22_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_22_full),
    .error        (_stageClearVec_reqQueue_fifo_22_error),
    .data_out     (_stageClearVec_reqQueue_fifo_22_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_22 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_22_enq_ready & stageClearVec_WaitReadQueue_22_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_22_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_22_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_22),
    .empty        (_stageClearVec_WaitReadQueue_fifo_22_empty),
    .almost_empty (stageClearVec_WaitReadQueue_22_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_22_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_22_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_22_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_22_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_23 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_23_enq_ready & stageClearVec_reqQueue_23_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_23_deq_ready & ~_stageClearVec_reqQueue_fifo_23_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_23),
    .empty        (_stageClearVec_reqQueue_fifo_23_empty),
    .almost_empty (stageClearVec_reqQueue_23_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_23_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_23_full),
    .error        (_stageClearVec_reqQueue_fifo_23_error),
    .data_out     (_stageClearVec_reqQueue_fifo_23_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_23 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_23_enq_ready & stageClearVec_WaitReadQueue_23_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_23_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_23_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_23),
    .empty        (_stageClearVec_WaitReadQueue_fifo_23_empty),
    .almost_empty (stageClearVec_WaitReadQueue_23_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_23_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_23_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_23_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_23_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_24 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_24_enq_ready & stageClearVec_reqQueue_24_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_24_deq_ready & ~_stageClearVec_reqQueue_fifo_24_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_24),
    .empty        (_stageClearVec_reqQueue_fifo_24_empty),
    .almost_empty (stageClearVec_reqQueue_24_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_24_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_24_full),
    .error        (_stageClearVec_reqQueue_fifo_24_error),
    .data_out     (_stageClearVec_reqQueue_fifo_24_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_24 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_24_enq_ready & stageClearVec_WaitReadQueue_24_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_24_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_24_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_24),
    .empty        (_stageClearVec_WaitReadQueue_fifo_24_empty),
    .almost_empty (stageClearVec_WaitReadQueue_24_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_24_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_24_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_24_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_24_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_25 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_25_enq_ready & stageClearVec_reqQueue_25_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_25_deq_ready & ~_stageClearVec_reqQueue_fifo_25_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_25),
    .empty        (_stageClearVec_reqQueue_fifo_25_empty),
    .almost_empty (stageClearVec_reqQueue_25_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_25_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_25_full),
    .error        (_stageClearVec_reqQueue_fifo_25_error),
    .data_out     (_stageClearVec_reqQueue_fifo_25_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_25 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_25_enq_ready & stageClearVec_WaitReadQueue_25_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_25_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_25_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_25),
    .empty        (_stageClearVec_WaitReadQueue_fifo_25_empty),
    .almost_empty (stageClearVec_WaitReadQueue_25_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_25_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_25_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_25_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_25_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_26 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_26_enq_ready & stageClearVec_reqQueue_26_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_26_deq_ready & ~_stageClearVec_reqQueue_fifo_26_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_26),
    .empty        (_stageClearVec_reqQueue_fifo_26_empty),
    .almost_empty (stageClearVec_reqQueue_26_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_26_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_26_full),
    .error        (_stageClearVec_reqQueue_fifo_26_error),
    .data_out     (_stageClearVec_reqQueue_fifo_26_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_26 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_26_enq_ready & stageClearVec_WaitReadQueue_26_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_26_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_26_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_26),
    .empty        (_stageClearVec_WaitReadQueue_fifo_26_empty),
    .almost_empty (stageClearVec_WaitReadQueue_26_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_26_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_26_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_26_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_26_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_27 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_27_enq_ready & stageClearVec_reqQueue_27_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_27_deq_ready & ~_stageClearVec_reqQueue_fifo_27_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_27),
    .empty        (_stageClearVec_reqQueue_fifo_27_empty),
    .almost_empty (stageClearVec_reqQueue_27_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_27_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_27_full),
    .error        (_stageClearVec_reqQueue_fifo_27_error),
    .data_out     (_stageClearVec_reqQueue_fifo_27_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_27 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_27_enq_ready & stageClearVec_WaitReadQueue_27_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_27_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_27_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_27),
    .empty        (_stageClearVec_WaitReadQueue_fifo_27_empty),
    .almost_empty (stageClearVec_WaitReadQueue_27_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_27_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_27_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_27_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_27_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_28 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_28_enq_ready & stageClearVec_reqQueue_28_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_28_deq_ready & ~_stageClearVec_reqQueue_fifo_28_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_28),
    .empty        (_stageClearVec_reqQueue_fifo_28_empty),
    .almost_empty (stageClearVec_reqQueue_28_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_28_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_28_full),
    .error        (_stageClearVec_reqQueue_fifo_28_error),
    .data_out     (_stageClearVec_reqQueue_fifo_28_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_28 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_28_enq_ready & stageClearVec_WaitReadQueue_28_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_28_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_28_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_28),
    .empty        (_stageClearVec_WaitReadQueue_fifo_28_empty),
    .almost_empty (stageClearVec_WaitReadQueue_28_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_28_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_28_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_28_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_28_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_29 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_29_enq_ready & stageClearVec_reqQueue_29_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_29_deq_ready & ~_stageClearVec_reqQueue_fifo_29_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_29),
    .empty        (_stageClearVec_reqQueue_fifo_29_empty),
    .almost_empty (stageClearVec_reqQueue_29_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_29_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_29_full),
    .error        (_stageClearVec_reqQueue_fifo_29_error),
    .data_out     (_stageClearVec_reqQueue_fifo_29_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_29 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_29_enq_ready & stageClearVec_WaitReadQueue_29_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_29_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_29_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_29),
    .empty        (_stageClearVec_WaitReadQueue_fifo_29_empty),
    .almost_empty (stageClearVec_WaitReadQueue_29_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_29_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_29_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_29_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_29_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_30 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_30_enq_ready & stageClearVec_reqQueue_30_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_30_deq_ready & ~_stageClearVec_reqQueue_fifo_30_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_30),
    .empty        (_stageClearVec_reqQueue_fifo_30_empty),
    .almost_empty (stageClearVec_reqQueue_30_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_30_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_30_full),
    .error        (_stageClearVec_reqQueue_fifo_30_error),
    .data_out     (_stageClearVec_reqQueue_fifo_30_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_30 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_30_enq_ready & stageClearVec_WaitReadQueue_30_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_30_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_30_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_30),
    .empty        (_stageClearVec_WaitReadQueue_fifo_30_empty),
    .almost_empty (stageClearVec_WaitReadQueue_30_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_30_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_30_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_30_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_30_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_reqQueue_fifo_31 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_reqQueue_31_enq_ready & stageClearVec_reqQueue_31_enq_valid)),
    .pop_req_n    (~(stageClearVec_reqQueue_31_deq_ready & ~_stageClearVec_reqQueue_fifo_31_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_reqQueue_dataIn_31),
    .empty        (_stageClearVec_reqQueue_fifo_31_empty),
    .almost_empty (stageClearVec_reqQueue_31_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_reqQueue_31_almostFull),
    .full         (_stageClearVec_reqQueue_fifo_31_full),
    .error        (_stageClearVec_reqQueue_fifo_31_error),
    .data_out     (_stageClearVec_reqQueue_fifo_31_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(75)
  ) stageClearVec_WaitReadQueue_fifo_31 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(stageClearVec_WaitReadQueue_31_enq_ready & stageClearVec_WaitReadQueue_31_enq_valid)),
    .pop_req_n    (~(stageClearVec_WaitReadQueue_31_deq_ready & ~_stageClearVec_WaitReadQueue_fifo_31_empty)),
    .diag_n       (1'h1),
    .data_in      (stageClearVec_WaitReadQueue_dataIn_31),
    .empty        (_stageClearVec_WaitReadQueue_fifo_31_empty),
    .almost_empty (stageClearVec_WaitReadQueue_31_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (stageClearVec_WaitReadQueue_31_almostFull),
    .full         (_stageClearVec_WaitReadQueue_fifo_31_full),
    .error        (_stageClearVec_WaitReadQueue_fifo_31_error),
    .data_out     (_stageClearVec_WaitReadQueue_fifo_31_data_out)
  );
  assign in_0_ready = in_0_ready_0;
  assign in_1_ready = in_1_ready_0;
  assign in_2_ready = in_2_ready_0;
  assign in_3_ready = in_3_ready_0;
  assign in_4_ready = in_4_ready_0;
  assign in_5_ready = in_5_ready_0;
  assign in_6_ready = in_6_ready_0;
  assign in_7_ready = in_7_ready_0;
  assign in_8_ready = in_8_ready_0;
  assign in_9_ready = in_9_ready_0;
  assign in_10_ready = in_10_ready_0;
  assign in_11_ready = in_11_ready_0;
  assign in_12_ready = in_12_ready_0;
  assign in_13_ready = in_13_ready_0;
  assign in_14_ready = in_14_ready_0;
  assign in_15_ready = in_15_ready_0;
  assign in_16_ready = in_16_ready_0;
  assign in_17_ready = in_17_ready_0;
  assign in_18_ready = in_18_ready_0;
  assign in_19_ready = in_19_ready_0;
  assign in_20_ready = in_20_ready_0;
  assign in_21_ready = in_21_ready_0;
  assign in_22_ready = in_22_ready_0;
  assign in_23_ready = in_23_ready_0;
  assign in_24_ready = in_24_ready_0;
  assign in_25_ready = in_25_ready_0;
  assign in_26_ready = in_26_ready_0;
  assign in_27_ready = in_27_ready_0;
  assign in_28_ready = in_28_ready_0;
  assign in_29_ready = in_29_ready_0;
  assign in_30_ready = in_30_ready_0;
  assign in_31_ready = in_31_ready_0;
  assign out_0_valid = out_0_valid_0;
  assign out_0_bits_ffoByOther = out_0_bits_ffoByOther_0;
  assign out_0_bits_writeData_data = out_0_bits_writeData_data_0;
  assign out_0_bits_writeData_mask = out_0_bits_writeData_mask_0;
  assign out_0_bits_writeData_groupCounter = out_0_bits_writeData_groupCounter_0;
  assign out_1_valid = out_1_valid_0;
  assign out_1_bits_ffoByOther = out_1_bits_ffoByOther_0;
  assign out_1_bits_writeData_data = out_1_bits_writeData_data_0;
  assign out_1_bits_writeData_mask = out_1_bits_writeData_mask_0;
  assign out_1_bits_writeData_groupCounter = out_1_bits_writeData_groupCounter_0;
  assign out_2_valid = out_2_valid_0;
  assign out_2_bits_ffoByOther = out_2_bits_ffoByOther_0;
  assign out_2_bits_writeData_data = out_2_bits_writeData_data_0;
  assign out_2_bits_writeData_mask = out_2_bits_writeData_mask_0;
  assign out_2_bits_writeData_groupCounter = out_2_bits_writeData_groupCounter_0;
  assign out_3_valid = out_3_valid_0;
  assign out_3_bits_ffoByOther = out_3_bits_ffoByOther_0;
  assign out_3_bits_writeData_data = out_3_bits_writeData_data_0;
  assign out_3_bits_writeData_mask = out_3_bits_writeData_mask_0;
  assign out_3_bits_writeData_groupCounter = out_3_bits_writeData_groupCounter_0;
  assign out_4_valid = out_4_valid_0;
  assign out_4_bits_ffoByOther = out_4_bits_ffoByOther_0;
  assign out_4_bits_writeData_data = out_4_bits_writeData_data_0;
  assign out_4_bits_writeData_mask = out_4_bits_writeData_mask_0;
  assign out_4_bits_writeData_groupCounter = out_4_bits_writeData_groupCounter_0;
  assign out_5_valid = out_5_valid_0;
  assign out_5_bits_ffoByOther = out_5_bits_ffoByOther_0;
  assign out_5_bits_writeData_data = out_5_bits_writeData_data_0;
  assign out_5_bits_writeData_mask = out_5_bits_writeData_mask_0;
  assign out_5_bits_writeData_groupCounter = out_5_bits_writeData_groupCounter_0;
  assign out_6_valid = out_6_valid_0;
  assign out_6_bits_ffoByOther = out_6_bits_ffoByOther_0;
  assign out_6_bits_writeData_data = out_6_bits_writeData_data_0;
  assign out_6_bits_writeData_mask = out_6_bits_writeData_mask_0;
  assign out_6_bits_writeData_groupCounter = out_6_bits_writeData_groupCounter_0;
  assign out_7_valid = out_7_valid_0;
  assign out_7_bits_ffoByOther = out_7_bits_ffoByOther_0;
  assign out_7_bits_writeData_data = out_7_bits_writeData_data_0;
  assign out_7_bits_writeData_mask = out_7_bits_writeData_mask_0;
  assign out_7_bits_writeData_groupCounter = out_7_bits_writeData_groupCounter_0;
  assign out_8_valid = out_8_valid_0;
  assign out_8_bits_ffoByOther = out_8_bits_ffoByOther_0;
  assign out_8_bits_writeData_data = out_8_bits_writeData_data_0;
  assign out_8_bits_writeData_mask = out_8_bits_writeData_mask_0;
  assign out_8_bits_writeData_groupCounter = out_8_bits_writeData_groupCounter_0;
  assign out_9_valid = out_9_valid_0;
  assign out_9_bits_ffoByOther = out_9_bits_ffoByOther_0;
  assign out_9_bits_writeData_data = out_9_bits_writeData_data_0;
  assign out_9_bits_writeData_mask = out_9_bits_writeData_mask_0;
  assign out_9_bits_writeData_groupCounter = out_9_bits_writeData_groupCounter_0;
  assign out_10_valid = out_10_valid_0;
  assign out_10_bits_ffoByOther = out_10_bits_ffoByOther_0;
  assign out_10_bits_writeData_data = out_10_bits_writeData_data_0;
  assign out_10_bits_writeData_mask = out_10_bits_writeData_mask_0;
  assign out_10_bits_writeData_groupCounter = out_10_bits_writeData_groupCounter_0;
  assign out_11_valid = out_11_valid_0;
  assign out_11_bits_ffoByOther = out_11_bits_ffoByOther_0;
  assign out_11_bits_writeData_data = out_11_bits_writeData_data_0;
  assign out_11_bits_writeData_mask = out_11_bits_writeData_mask_0;
  assign out_11_bits_writeData_groupCounter = out_11_bits_writeData_groupCounter_0;
  assign out_12_valid = out_12_valid_0;
  assign out_12_bits_ffoByOther = out_12_bits_ffoByOther_0;
  assign out_12_bits_writeData_data = out_12_bits_writeData_data_0;
  assign out_12_bits_writeData_mask = out_12_bits_writeData_mask_0;
  assign out_12_bits_writeData_groupCounter = out_12_bits_writeData_groupCounter_0;
  assign out_13_valid = out_13_valid_0;
  assign out_13_bits_ffoByOther = out_13_bits_ffoByOther_0;
  assign out_13_bits_writeData_data = out_13_bits_writeData_data_0;
  assign out_13_bits_writeData_mask = out_13_bits_writeData_mask_0;
  assign out_13_bits_writeData_groupCounter = out_13_bits_writeData_groupCounter_0;
  assign out_14_valid = out_14_valid_0;
  assign out_14_bits_ffoByOther = out_14_bits_ffoByOther_0;
  assign out_14_bits_writeData_data = out_14_bits_writeData_data_0;
  assign out_14_bits_writeData_mask = out_14_bits_writeData_mask_0;
  assign out_14_bits_writeData_groupCounter = out_14_bits_writeData_groupCounter_0;
  assign out_15_valid = out_15_valid_0;
  assign out_15_bits_ffoByOther = out_15_bits_ffoByOther_0;
  assign out_15_bits_writeData_data = out_15_bits_writeData_data_0;
  assign out_15_bits_writeData_mask = out_15_bits_writeData_mask_0;
  assign out_15_bits_writeData_groupCounter = out_15_bits_writeData_groupCounter_0;
  assign out_16_valid = out_16_valid_0;
  assign out_16_bits_ffoByOther = out_16_bits_ffoByOther_0;
  assign out_16_bits_writeData_data = out_16_bits_writeData_data_0;
  assign out_16_bits_writeData_mask = out_16_bits_writeData_mask_0;
  assign out_16_bits_writeData_groupCounter = out_16_bits_writeData_groupCounter_0;
  assign out_17_valid = out_17_valid_0;
  assign out_17_bits_ffoByOther = out_17_bits_ffoByOther_0;
  assign out_17_bits_writeData_data = out_17_bits_writeData_data_0;
  assign out_17_bits_writeData_mask = out_17_bits_writeData_mask_0;
  assign out_17_bits_writeData_groupCounter = out_17_bits_writeData_groupCounter_0;
  assign out_18_valid = out_18_valid_0;
  assign out_18_bits_ffoByOther = out_18_bits_ffoByOther_0;
  assign out_18_bits_writeData_data = out_18_bits_writeData_data_0;
  assign out_18_bits_writeData_mask = out_18_bits_writeData_mask_0;
  assign out_18_bits_writeData_groupCounter = out_18_bits_writeData_groupCounter_0;
  assign out_19_valid = out_19_valid_0;
  assign out_19_bits_ffoByOther = out_19_bits_ffoByOther_0;
  assign out_19_bits_writeData_data = out_19_bits_writeData_data_0;
  assign out_19_bits_writeData_mask = out_19_bits_writeData_mask_0;
  assign out_19_bits_writeData_groupCounter = out_19_bits_writeData_groupCounter_0;
  assign out_20_valid = out_20_valid_0;
  assign out_20_bits_ffoByOther = out_20_bits_ffoByOther_0;
  assign out_20_bits_writeData_data = out_20_bits_writeData_data_0;
  assign out_20_bits_writeData_mask = out_20_bits_writeData_mask_0;
  assign out_20_bits_writeData_groupCounter = out_20_bits_writeData_groupCounter_0;
  assign out_21_valid = out_21_valid_0;
  assign out_21_bits_ffoByOther = out_21_bits_ffoByOther_0;
  assign out_21_bits_writeData_data = out_21_bits_writeData_data_0;
  assign out_21_bits_writeData_mask = out_21_bits_writeData_mask_0;
  assign out_21_bits_writeData_groupCounter = out_21_bits_writeData_groupCounter_0;
  assign out_22_valid = out_22_valid_0;
  assign out_22_bits_ffoByOther = out_22_bits_ffoByOther_0;
  assign out_22_bits_writeData_data = out_22_bits_writeData_data_0;
  assign out_22_bits_writeData_mask = out_22_bits_writeData_mask_0;
  assign out_22_bits_writeData_groupCounter = out_22_bits_writeData_groupCounter_0;
  assign out_23_valid = out_23_valid_0;
  assign out_23_bits_ffoByOther = out_23_bits_ffoByOther_0;
  assign out_23_bits_writeData_data = out_23_bits_writeData_data_0;
  assign out_23_bits_writeData_mask = out_23_bits_writeData_mask_0;
  assign out_23_bits_writeData_groupCounter = out_23_bits_writeData_groupCounter_0;
  assign out_24_valid = out_24_valid_0;
  assign out_24_bits_ffoByOther = out_24_bits_ffoByOther_0;
  assign out_24_bits_writeData_data = out_24_bits_writeData_data_0;
  assign out_24_bits_writeData_mask = out_24_bits_writeData_mask_0;
  assign out_24_bits_writeData_groupCounter = out_24_bits_writeData_groupCounter_0;
  assign out_25_valid = out_25_valid_0;
  assign out_25_bits_ffoByOther = out_25_bits_ffoByOther_0;
  assign out_25_bits_writeData_data = out_25_bits_writeData_data_0;
  assign out_25_bits_writeData_mask = out_25_bits_writeData_mask_0;
  assign out_25_bits_writeData_groupCounter = out_25_bits_writeData_groupCounter_0;
  assign out_26_valid = out_26_valid_0;
  assign out_26_bits_ffoByOther = out_26_bits_ffoByOther_0;
  assign out_26_bits_writeData_data = out_26_bits_writeData_data_0;
  assign out_26_bits_writeData_mask = out_26_bits_writeData_mask_0;
  assign out_26_bits_writeData_groupCounter = out_26_bits_writeData_groupCounter_0;
  assign out_27_valid = out_27_valid_0;
  assign out_27_bits_ffoByOther = out_27_bits_ffoByOther_0;
  assign out_27_bits_writeData_data = out_27_bits_writeData_data_0;
  assign out_27_bits_writeData_mask = out_27_bits_writeData_mask_0;
  assign out_27_bits_writeData_groupCounter = out_27_bits_writeData_groupCounter_0;
  assign out_28_valid = out_28_valid_0;
  assign out_28_bits_ffoByOther = out_28_bits_ffoByOther_0;
  assign out_28_bits_writeData_data = out_28_bits_writeData_data_0;
  assign out_28_bits_writeData_mask = out_28_bits_writeData_mask_0;
  assign out_28_bits_writeData_groupCounter = out_28_bits_writeData_groupCounter_0;
  assign out_29_valid = out_29_valid_0;
  assign out_29_bits_ffoByOther = out_29_bits_ffoByOther_0;
  assign out_29_bits_writeData_data = out_29_bits_writeData_data_0;
  assign out_29_bits_writeData_mask = out_29_bits_writeData_mask_0;
  assign out_29_bits_writeData_groupCounter = out_29_bits_writeData_groupCounter_0;
  assign out_30_valid = out_30_valid_0;
  assign out_30_bits_ffoByOther = out_30_bits_ffoByOther_0;
  assign out_30_bits_writeData_data = out_30_bits_writeData_data_0;
  assign out_30_bits_writeData_mask = out_30_bits_writeData_mask_0;
  assign out_30_bits_writeData_groupCounter = out_30_bits_writeData_groupCounter_0;
  assign out_31_valid = out_31_valid_0;
  assign out_31_bits_ffoByOther = out_31_bits_ffoByOther_0;
  assign out_31_bits_writeData_data = out_31_bits_writeData_data_0;
  assign out_31_bits_writeData_mask = out_31_bits_writeData_mask_0;
  assign out_31_bits_writeData_groupCounter = out_31_bits_writeData_groupCounter_0;
  assign readChannel_0_valid = readChannel_0_valid_0;
  assign readChannel_0_bits_vs = readChannel_0_bits_vs_0;
  assign readChannel_0_bits_offset = readChannel_0_bits_offset_0;
  assign readChannel_1_valid = readChannel_1_valid_0;
  assign readChannel_1_bits_vs = readChannel_1_bits_vs_0;
  assign readChannel_1_bits_offset = readChannel_1_bits_offset_0;
  assign readChannel_2_valid = readChannel_2_valid_0;
  assign readChannel_2_bits_vs = readChannel_2_bits_vs_0;
  assign readChannel_2_bits_offset = readChannel_2_bits_offset_0;
  assign readChannel_3_valid = readChannel_3_valid_0;
  assign readChannel_3_bits_vs = readChannel_3_bits_vs_0;
  assign readChannel_3_bits_offset = readChannel_3_bits_offset_0;
  assign readChannel_4_valid = readChannel_4_valid_0;
  assign readChannel_4_bits_vs = readChannel_4_bits_vs_0;
  assign readChannel_4_bits_offset = readChannel_4_bits_offset_0;
  assign readChannel_5_valid = readChannel_5_valid_0;
  assign readChannel_5_bits_vs = readChannel_5_bits_vs_0;
  assign readChannel_5_bits_offset = readChannel_5_bits_offset_0;
  assign readChannel_6_valid = readChannel_6_valid_0;
  assign readChannel_6_bits_vs = readChannel_6_bits_vs_0;
  assign readChannel_6_bits_offset = readChannel_6_bits_offset_0;
  assign readChannel_7_valid = readChannel_7_valid_0;
  assign readChannel_7_bits_vs = readChannel_7_bits_vs_0;
  assign readChannel_7_bits_offset = readChannel_7_bits_offset_0;
  assign readChannel_8_valid = readChannel_8_valid_0;
  assign readChannel_8_bits_vs = readChannel_8_bits_vs_0;
  assign readChannel_8_bits_offset = readChannel_8_bits_offset_0;
  assign readChannel_9_valid = readChannel_9_valid_0;
  assign readChannel_9_bits_vs = readChannel_9_bits_vs_0;
  assign readChannel_9_bits_offset = readChannel_9_bits_offset_0;
  assign readChannel_10_valid = readChannel_10_valid_0;
  assign readChannel_10_bits_vs = readChannel_10_bits_vs_0;
  assign readChannel_10_bits_offset = readChannel_10_bits_offset_0;
  assign readChannel_11_valid = readChannel_11_valid_0;
  assign readChannel_11_bits_vs = readChannel_11_bits_vs_0;
  assign readChannel_11_bits_offset = readChannel_11_bits_offset_0;
  assign readChannel_12_valid = readChannel_12_valid_0;
  assign readChannel_12_bits_vs = readChannel_12_bits_vs_0;
  assign readChannel_12_bits_offset = readChannel_12_bits_offset_0;
  assign readChannel_13_valid = readChannel_13_valid_0;
  assign readChannel_13_bits_vs = readChannel_13_bits_vs_0;
  assign readChannel_13_bits_offset = readChannel_13_bits_offset_0;
  assign readChannel_14_valid = readChannel_14_valid_0;
  assign readChannel_14_bits_vs = readChannel_14_bits_vs_0;
  assign readChannel_14_bits_offset = readChannel_14_bits_offset_0;
  assign readChannel_15_valid = readChannel_15_valid_0;
  assign readChannel_15_bits_vs = readChannel_15_bits_vs_0;
  assign readChannel_15_bits_offset = readChannel_15_bits_offset_0;
  assign readChannel_16_valid = readChannel_16_valid_0;
  assign readChannel_16_bits_vs = readChannel_16_bits_vs_0;
  assign readChannel_16_bits_offset = readChannel_16_bits_offset_0;
  assign readChannel_17_valid = readChannel_17_valid_0;
  assign readChannel_17_bits_vs = readChannel_17_bits_vs_0;
  assign readChannel_17_bits_offset = readChannel_17_bits_offset_0;
  assign readChannel_18_valid = readChannel_18_valid_0;
  assign readChannel_18_bits_vs = readChannel_18_bits_vs_0;
  assign readChannel_18_bits_offset = readChannel_18_bits_offset_0;
  assign readChannel_19_valid = readChannel_19_valid_0;
  assign readChannel_19_bits_vs = readChannel_19_bits_vs_0;
  assign readChannel_19_bits_offset = readChannel_19_bits_offset_0;
  assign readChannel_20_valid = readChannel_20_valid_0;
  assign readChannel_20_bits_vs = readChannel_20_bits_vs_0;
  assign readChannel_20_bits_offset = readChannel_20_bits_offset_0;
  assign readChannel_21_valid = readChannel_21_valid_0;
  assign readChannel_21_bits_vs = readChannel_21_bits_vs_0;
  assign readChannel_21_bits_offset = readChannel_21_bits_offset_0;
  assign readChannel_22_valid = readChannel_22_valid_0;
  assign readChannel_22_bits_vs = readChannel_22_bits_vs_0;
  assign readChannel_22_bits_offset = readChannel_22_bits_offset_0;
  assign readChannel_23_valid = readChannel_23_valid_0;
  assign readChannel_23_bits_vs = readChannel_23_bits_vs_0;
  assign readChannel_23_bits_offset = readChannel_23_bits_offset_0;
  assign readChannel_24_valid = readChannel_24_valid_0;
  assign readChannel_24_bits_vs = readChannel_24_bits_vs_0;
  assign readChannel_24_bits_offset = readChannel_24_bits_offset_0;
  assign readChannel_25_valid = readChannel_25_valid_0;
  assign readChannel_25_bits_vs = readChannel_25_bits_vs_0;
  assign readChannel_25_bits_offset = readChannel_25_bits_offset_0;
  assign readChannel_26_valid = readChannel_26_valid_0;
  assign readChannel_26_bits_vs = readChannel_26_bits_vs_0;
  assign readChannel_26_bits_offset = readChannel_26_bits_offset_0;
  assign readChannel_27_valid = readChannel_27_valid_0;
  assign readChannel_27_bits_vs = readChannel_27_bits_vs_0;
  assign readChannel_27_bits_offset = readChannel_27_bits_offset_0;
  assign readChannel_28_valid = readChannel_28_valid_0;
  assign readChannel_28_bits_vs = readChannel_28_bits_vs_0;
  assign readChannel_28_bits_offset = readChannel_28_bits_offset_0;
  assign readChannel_29_valid = readChannel_29_valid_0;
  assign readChannel_29_bits_vs = readChannel_29_bits_vs_0;
  assign readChannel_29_bits_offset = readChannel_29_bits_offset_0;
  assign readChannel_30_valid = readChannel_30_valid_0;
  assign readChannel_30_bits_vs = readChannel_30_bits_vs_0;
  assign readChannel_30_bits_offset = readChannel_30_bits_offset_0;
  assign readChannel_31_valid = readChannel_31_valid_0;
  assign readChannel_31_bits_vs = readChannel_31_bits_vs_0;
  assign readChannel_31_bits_offset = readChannel_31_bits_offset_0;
  assign stageClear =
    stageClearVec_0 & stageClearVec_1 & stageClearVec_2 & stageClearVec_3 & stageClearVec_4 & stageClearVec_5 & stageClearVec_6 & stageClearVec_7 & stageClearVec_8 & stageClearVec_9 & stageClearVec_10 & stageClearVec_11 & stageClearVec_12
    & stageClearVec_13 & stageClearVec_14 & stageClearVec_15 & stageClearVec_16 & stageClearVec_17 & stageClearVec_18 & stageClearVec_19 & stageClearVec_20 & stageClearVec_21 & stageClearVec_22 & stageClearVec_23 & stageClearVec_24
    & stageClearVec_25 & stageClearVec_26 & stageClearVec_27 & stageClearVec_28 & stageClearVec_29 & stageClearVec_30 & stageClearVec_31;
endmodule

