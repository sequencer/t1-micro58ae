module QDS(
  input  [6:0] input_partialReminderCarry,
               input_partialReminderSum,
  input  [2:0] input_partialDivider,
  output [4:0] output_selectedQuotientOH
);

  wire [7:0][6:0] _GEN = '{7'h6A, 7'h6C, 7'h6C, 7'h6E, 7'h70, 7'h70, 7'h72, 7'h74};
  wire [7:0][6:0] _GEN_0 = '{7'h78, 7'h78, 7'h7A, 7'h7A, 7'h7C, 7'h7C, 7'h7C, 7'h7C};
  wire [7:0][6:0] _GEN_1 = '{7'h8, 7'h8, 7'h8, 7'h6, 7'h6, 7'h6, 7'h5, 7'h4};
  wire [7:0][6:0] _GEN_2 = '{7'h17, 7'h16, 7'h14, 7'h12, 7'h11, 7'h10, 7'hE, 7'hD};
  wire [6:0]      selectRom_0_0 = 7'h74;
  wire [6:0]      selectRom_0_2 = 7'h4;
  wire [6:0]      selectRom_0_3 = 7'hD;
  wire [6:0]      selectRom_1_0 = 7'h72;
  wire [6:0]      selectRom_1_2 = 7'h5;
  wire [6:0]      selectRom_1_3 = 7'hE;
  wire [6:0]      selectRom_2_3 = 7'h10;
  wire [6:0]      selectRom_2_0 = 7'h70;
  wire [6:0]      selectRom_3_0 = 7'h70;
  wire [6:0]      selectRom_0_1 = 7'h7C;
  wire [6:0]      selectRom_1_1 = 7'h7C;
  wire [6:0]      selectRom_2_1 = 7'h7C;
  wire [6:0]      selectRom_3_1 = 7'h7C;
  wire [6:0]      selectRom_3_3 = 7'h11;
  wire [6:0]      selectRom_4_0 = 7'h6E;
  wire [6:0]      selectRom_2_2 = 7'h6;
  wire [6:0]      selectRom_3_2 = 7'h6;
  wire [6:0]      selectRom_4_2 = 7'h6;
  wire [6:0]      selectRom_4_3 = 7'h12;
  wire [6:0]      selectRom_4_1 = 7'h7A;
  wire [6:0]      selectRom_5_1 = 7'h7A;
  wire [6:0]      selectRom_5_3 = 7'h14;
  wire [6:0]      selectRom_5_0 = 7'h6C;
  wire [6:0]      selectRom_6_0 = 7'h6C;
  wire [6:0]      selectRom_6_3 = 7'h16;
  wire [6:0]      selectRom_7_0 = 7'h6A;
  wire [6:0]      selectRom_6_1 = 7'h78;
  wire [6:0]      selectRom_7_1 = 7'h78;
  wire [6:0]      selectRom_5_2 = 7'h8;
  wire [6:0]      selectRom_6_2 = 7'h8;
  wire [6:0]      selectRom_7_2 = 7'h8;
  wire [6:0]      selectRom_7_3 = 7'h17;
  wire [6:0]      yTruncate = input_partialReminderCarry + input_partialReminderSum;
  wire            selectPoints_fillBit = yTruncate[6];
  wire            selectPoints_fillBit_2 = yTruncate[6];
  wire            selectPoints_fillBit_4 = yTruncate[6];
  wire            selectPoints_fillBit_6 = yTruncate[6];
  wire            selectPoints_fillBit_1 = _GEN[input_partialDivider][6];
  wire [7:0]      _selectPoints_T_2 = {selectPoints_fillBit, yTruncate} + {selectPoints_fillBit_1, _GEN[input_partialDivider]};
  wire            selectPoints_fillBit_3 = _GEN_0[input_partialDivider][6];
  wire [7:0]      _selectPoints_T_7 = {selectPoints_fillBit_2, yTruncate} + {selectPoints_fillBit_3, _GEN_0[input_partialDivider]};
  wire            selectPoints_fillBit_5 = _GEN_1[input_partialDivider][6];
  wire [7:0]      _selectPoints_T_12 = {selectPoints_fillBit_4, yTruncate} + {selectPoints_fillBit_5, _GEN_1[input_partialDivider]};
  wire            selectPoints_fillBit_7 = _GEN_2[input_partialDivider][6];
  wire [7:0]      _selectPoints_T_17 = {selectPoints_fillBit_6, yTruncate} + {selectPoints_fillBit_7, _GEN_2[input_partialDivider]};
  wire [1:0]      selectPoints_lo = {_selectPoints_T_7[7], _selectPoints_T_2[7]};
  wire [1:0]      selectPoints_hi = {_selectPoints_T_17[7], _selectPoints_T_12[7]};
  wire [3:0]      selectPoints = {selectPoints_hi, selectPoints_lo};
  wire [3:0]      output_selectedQuotientOH_plaInput = selectPoints;
  wire [3:0]      output_selectedQuotientOH_invInputs = ~output_selectedQuotientOH_plaInput;
  wire [4:0]      output_selectedQuotientOH_invMatrixOutputs;
  wire            output_selectedQuotientOH_andMatrixOutputs_andMatrixInput_0 = output_selectedQuotientOH_invInputs[0];
  wire            output_selectedQuotientOH_andMatrixOutputs_1_2 = output_selectedQuotientOH_andMatrixOutputs_andMatrixInput_0;
  wire            output_selectedQuotientOH_andMatrixOutputs_andMatrixInput_0_1 = output_selectedQuotientOH_invInputs[1];
  wire            output_selectedQuotientOH_andMatrixOutputs_andMatrixInput_1 = output_selectedQuotientOH_invInputs[1];
  wire            output_selectedQuotientOH_andMatrixOutputs_2_2 = output_selectedQuotientOH_andMatrixOutputs_andMatrixInput_0_1;
  wire            output_selectedQuotientOH_andMatrixOutputs_andMatrixInput_0_2 = output_selectedQuotientOH_invInputs[2];
  wire            output_selectedQuotientOH_andMatrixOutputs_andMatrixInput_2 = output_selectedQuotientOH_invInputs[2];
  wire            output_selectedQuotientOH_andMatrixOutputs_4_2 = output_selectedQuotientOH_andMatrixOutputs_andMatrixInput_0_2;
  wire            output_selectedQuotientOH_andMatrixOutputs_andMatrixInput_0_3 = output_selectedQuotientOH_invInputs[3];
  wire            output_selectedQuotientOH_andMatrixOutputs_andMatrixInput_3 = output_selectedQuotientOH_invInputs[3];
  wire            output_selectedQuotientOH_andMatrixOutputs_0_2 = output_selectedQuotientOH_andMatrixOutputs_andMatrixInput_0_3;
  wire            output_selectedQuotientOH_andMatrixOutputs_andMatrixInput_0_4 = output_selectedQuotientOH_plaInput[0];
  wire            output_selectedQuotientOH_andMatrixOutputs_andMatrixInput_0_5 = output_selectedQuotientOH_plaInput[0];
  wire            output_selectedQuotientOH_andMatrixOutputs_andMatrixInput_0_6 = output_selectedQuotientOH_plaInput[0];
  wire            output_selectedQuotientOH_andMatrixOutputs_3_2 = &{output_selectedQuotientOH_andMatrixOutputs_andMatrixInput_0_4, output_selectedQuotientOH_andMatrixOutputs_andMatrixInput_1};
  wire            output_selectedQuotientOH_andMatrixOutputs_andMatrixInput_1_1 = output_selectedQuotientOH_plaInput[1];
  wire            output_selectedQuotientOH_andMatrixOutputs_andMatrixInput_1_2 = output_selectedQuotientOH_plaInput[1];
  wire [1:0]      output_selectedQuotientOH_andMatrixOutputs_hi = {output_selectedQuotientOH_andMatrixOutputs_andMatrixInput_0_5, output_selectedQuotientOH_andMatrixOutputs_andMatrixInput_1_1};
  wire            output_selectedQuotientOH_andMatrixOutputs_6_2 = &{output_selectedQuotientOH_andMatrixOutputs_hi, output_selectedQuotientOH_andMatrixOutputs_andMatrixInput_2};
  wire            output_selectedQuotientOH_andMatrixOutputs_andMatrixInput_2_1 = output_selectedQuotientOH_plaInput[2];
  wire [1:0]      output_selectedQuotientOH_andMatrixOutputs_lo = {output_selectedQuotientOH_andMatrixOutputs_andMatrixInput_2_1, output_selectedQuotientOH_andMatrixOutputs_andMatrixInput_3};
  wire [1:0]      output_selectedQuotientOH_andMatrixOutputs_hi_1 = {output_selectedQuotientOH_andMatrixOutputs_andMatrixInput_0_6, output_selectedQuotientOH_andMatrixOutputs_andMatrixInput_1_2};
  wire            output_selectedQuotientOH_andMatrixOutputs_5_2 = &{output_selectedQuotientOH_andMatrixOutputs_hi_1, output_selectedQuotientOH_andMatrixOutputs_lo};
  wire [1:0]      output_selectedQuotientOH_orMatrixOutputs_lo = {output_selectedQuotientOH_andMatrixOutputs_4_2, output_selectedQuotientOH_andMatrixOutputs_0_2};
  wire [1:0]      output_selectedQuotientOH_orMatrixOutputs_hi = {output_selectedQuotientOH_andMatrixOutputs_1_2, output_selectedQuotientOH_andMatrixOutputs_2_2};
  wire [1:0]      output_selectedQuotientOH_orMatrixOutputs_lo_1 = {output_selectedQuotientOH_andMatrixOutputs_5_2, |{output_selectedQuotientOH_orMatrixOutputs_hi, output_selectedQuotientOH_orMatrixOutputs_lo}};
  wire [1:0]      output_selectedQuotientOH_orMatrixOutputs_hi_hi = {output_selectedQuotientOH_andMatrixOutputs_1_2, output_selectedQuotientOH_andMatrixOutputs_3_2};
  wire [2:0]      output_selectedQuotientOH_orMatrixOutputs_hi_1 = {output_selectedQuotientOH_orMatrixOutputs_hi_hi, output_selectedQuotientOH_andMatrixOutputs_6_2};
  wire [4:0]      output_selectedQuotientOH_orMatrixOutputs = {output_selectedQuotientOH_orMatrixOutputs_hi_1, output_selectedQuotientOH_orMatrixOutputs_lo_1};
  wire [1:0]      output_selectedQuotientOH_invMatrixOutputs_lo = {output_selectedQuotientOH_orMatrixOutputs[1], ~(output_selectedQuotientOH_orMatrixOutputs[0])};
  wire [1:0]      output_selectedQuotientOH_invMatrixOutputs_hi_hi = output_selectedQuotientOH_orMatrixOutputs[4:3];
  wire [2:0]      output_selectedQuotientOH_invMatrixOutputs_hi = {output_selectedQuotientOH_invMatrixOutputs_hi_hi, output_selectedQuotientOH_orMatrixOutputs[2]};
  assign output_selectedQuotientOH_invMatrixOutputs = {output_selectedQuotientOH_invMatrixOutputs_hi, output_selectedQuotientOH_invMatrixOutputs_lo};
  wire [4:0]      output_selectedQuotientOH_plaOutput = output_selectedQuotientOH_invMatrixOutputs;
  assign output_selectedQuotientOH = output_selectedQuotientOH_plaOutput;
endmodule

