
// Include register initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for register randomization.

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_
module T1TokenManager(
  input        clock,
               reset,
               instructionIssue_valid,
  input  [2:0] instructionIssue_bits_instructionIndex,
  input        instructionIssue_bits_writeV0,
               instructionIssue_bits_useV0AsMask,
               instructionIssue_bits_toLane,
               instructionIssue_bits_toMask,
               lsuWriteV0_0_valid,
  input  [2:0] lsuWriteV0_0_bits,
  input        lsuWriteV0_1_valid,
  input  [2:0] lsuWriteV0_1_bits,
  input        lsuWriteV0_2_valid,
  input  [2:0] lsuWriteV0_2_bits,
  input        lsuWriteV0_3_valid,
  input  [2:0] lsuWriteV0_3_bits,
  input        lsuWriteV0_4_valid,
  input  [2:0] lsuWriteV0_4_bits,
  input        lsuWriteV0_5_valid,
  input  [2:0] lsuWriteV0_5_bits,
  input        lsuWriteV0_6_valid,
  input  [2:0] lsuWriteV0_6_bits,
  input        lsuWriteV0_7_valid,
  input  [2:0] lsuWriteV0_7_bits,
  input        lsuWriteV0_8_valid,
  input  [2:0] lsuWriteV0_8_bits,
  input        lsuWriteV0_9_valid,
  input  [2:0] lsuWriteV0_9_bits,
  input        lsuWriteV0_10_valid,
  input  [2:0] lsuWriteV0_10_bits,
  input        lsuWriteV0_11_valid,
  input  [2:0] lsuWriteV0_11_bits,
  input        lsuWriteV0_12_valid,
  input  [2:0] lsuWriteV0_12_bits,
  input        lsuWriteV0_13_valid,
  input  [2:0] lsuWriteV0_13_bits,
  input        lsuWriteV0_14_valid,
  input  [2:0] lsuWriteV0_14_bits,
  input        lsuWriteV0_15_valid,
  input  [2:0] lsuWriteV0_15_bits,
  output       issueAllow,
  input  [7:0] instructionFinish_0,
               instructionFinish_1,
               instructionFinish_2,
               instructionFinish_3,
               instructionFinish_4,
               instructionFinish_5,
               instructionFinish_6,
               instructionFinish_7,
               instructionFinish_8,
               instructionFinish_9,
               instructionFinish_10,
               instructionFinish_11,
               instructionFinish_12,
               instructionFinish_13,
               instructionFinish_14,
               instructionFinish_15,
  output [7:0] v0WriteValid,
  input        maskUnitFree
);

  wire [7:0] issueIndex1H = 8'h1 << instructionIssue_bits_instructionIndex;
  wire [7:0] v0WriteValidVec_lsuWriteSet = lsuWriteV0_0_valid ? 8'h1 << lsuWriteV0_0_bits : 8'h0;
  wire       _maskUnitWriteV0_set_T = instructionIssue_valid & instructionIssue_bits_writeV0;
  wire       _GEN = _maskUnitWriteV0_set_T & instructionIssue_bits_toLane;
  wire       v0WriteValidVec_v0WriteIssue;
  assign v0WriteValidVec_v0WriteIssue = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_1;
  assign v0WriteValidVec_v0WriteIssue_1 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_2;
  assign v0WriteValidVec_v0WriteIssue_2 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_3;
  assign v0WriteValidVec_v0WriteIssue_3 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_4;
  assign v0WriteValidVec_v0WriteIssue_4 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_5;
  assign v0WriteValidVec_v0WriteIssue_5 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_6;
  assign v0WriteValidVec_v0WriteIssue_6 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_7;
  assign v0WriteValidVec_v0WriteIssue_7 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_8;
  assign v0WriteValidVec_v0WriteIssue_8 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_9;
  assign v0WriteValidVec_v0WriteIssue_9 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_10;
  assign v0WriteValidVec_v0WriteIssue_10 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_11;
  assign v0WriteValidVec_v0WriteIssue_11 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_12;
  assign v0WriteValidVec_v0WriteIssue_12 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_13;
  assign v0WriteValidVec_v0WriteIssue_13 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_14;
  assign v0WriteValidVec_v0WriteIssue_14 = _GEN;
  wire       v0WriteValidVec_v0WriteIssue_15;
  assign v0WriteValidVec_v0WriteIssue_15 = _GEN;
  wire [7:0] v0WriteValidVec_updateOH = v0WriteValidVec_v0WriteIssue ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res;
  reg        v0WriteValidVec_res_1;
  reg        v0WriteValidVec_res_2;
  reg        v0WriteValidVec_res_3;
  reg        v0WriteValidVec_res_4;
  reg        v0WriteValidVec_res_5;
  reg        v0WriteValidVec_res_6;
  reg        v0WriteValidVec_res_7;
  wire [1:0] v0WriteValidVec_lo_lo = {v0WriteValidVec_res_1, v0WriteValidVec_res};
  wire [1:0] v0WriteValidVec_lo_hi = {v0WriteValidVec_res_3, v0WriteValidVec_res_2};
  wire [3:0] v0WriteValidVec_lo = {v0WriteValidVec_lo_hi, v0WriteValidVec_lo_lo};
  wire [1:0] v0WriteValidVec_hi_lo = {v0WriteValidVec_res_5, v0WriteValidVec_res_4};
  wire [1:0] v0WriteValidVec_hi_hi = {v0WriteValidVec_res_7, v0WriteValidVec_res_6};
  wire [3:0] v0WriteValidVec_hi = {v0WriteValidVec_hi_hi, v0WriteValidVec_hi_lo};
  wire [7:0] v0WriteValidVec_0 = {v0WriteValidVec_hi, v0WriteValidVec_lo};
  wire [7:0] v0WriteValidVec_lsuWriteSet_1 = lsuWriteV0_1_valid ? 8'h1 << lsuWriteV0_1_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_1 = v0WriteValidVec_v0WriteIssue_1 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_8;
  reg        v0WriteValidVec_res_9;
  reg        v0WriteValidVec_res_10;
  reg        v0WriteValidVec_res_11;
  reg        v0WriteValidVec_res_12;
  reg        v0WriteValidVec_res_13;
  reg        v0WriteValidVec_res_14;
  reg        v0WriteValidVec_res_15;
  wire [1:0] v0WriteValidVec_lo_lo_1 = {v0WriteValidVec_res_9, v0WriteValidVec_res_8};
  wire [1:0] v0WriteValidVec_lo_hi_1 = {v0WriteValidVec_res_11, v0WriteValidVec_res_10};
  wire [3:0] v0WriteValidVec_lo_1 = {v0WriteValidVec_lo_hi_1, v0WriteValidVec_lo_lo_1};
  wire [1:0] v0WriteValidVec_hi_lo_1 = {v0WriteValidVec_res_13, v0WriteValidVec_res_12};
  wire [1:0] v0WriteValidVec_hi_hi_1 = {v0WriteValidVec_res_15, v0WriteValidVec_res_14};
  wire [3:0] v0WriteValidVec_hi_1 = {v0WriteValidVec_hi_hi_1, v0WriteValidVec_hi_lo_1};
  wire [7:0] v0WriteValidVec_1 = {v0WriteValidVec_hi_1, v0WriteValidVec_lo_1};
  wire [7:0] v0WriteValidVec_lsuWriteSet_2 = lsuWriteV0_2_valid ? 8'h1 << lsuWriteV0_2_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_2 = v0WriteValidVec_v0WriteIssue_2 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_16;
  reg        v0WriteValidVec_res_17;
  reg        v0WriteValidVec_res_18;
  reg        v0WriteValidVec_res_19;
  reg        v0WriteValidVec_res_20;
  reg        v0WriteValidVec_res_21;
  reg        v0WriteValidVec_res_22;
  reg        v0WriteValidVec_res_23;
  wire [1:0] v0WriteValidVec_lo_lo_2 = {v0WriteValidVec_res_17, v0WriteValidVec_res_16};
  wire [1:0] v0WriteValidVec_lo_hi_2 = {v0WriteValidVec_res_19, v0WriteValidVec_res_18};
  wire [3:0] v0WriteValidVec_lo_2 = {v0WriteValidVec_lo_hi_2, v0WriteValidVec_lo_lo_2};
  wire [1:0] v0WriteValidVec_hi_lo_2 = {v0WriteValidVec_res_21, v0WriteValidVec_res_20};
  wire [1:0] v0WriteValidVec_hi_hi_2 = {v0WriteValidVec_res_23, v0WriteValidVec_res_22};
  wire [3:0] v0WriteValidVec_hi_2 = {v0WriteValidVec_hi_hi_2, v0WriteValidVec_hi_lo_2};
  wire [7:0] v0WriteValidVec_2 = {v0WriteValidVec_hi_2, v0WriteValidVec_lo_2};
  wire [7:0] v0WriteValidVec_lsuWriteSet_3 = lsuWriteV0_3_valid ? 8'h1 << lsuWriteV0_3_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_3 = v0WriteValidVec_v0WriteIssue_3 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_24;
  reg        v0WriteValidVec_res_25;
  reg        v0WriteValidVec_res_26;
  reg        v0WriteValidVec_res_27;
  reg        v0WriteValidVec_res_28;
  reg        v0WriteValidVec_res_29;
  reg        v0WriteValidVec_res_30;
  reg        v0WriteValidVec_res_31;
  wire [1:0] v0WriteValidVec_lo_lo_3 = {v0WriteValidVec_res_25, v0WriteValidVec_res_24};
  wire [1:0] v0WriteValidVec_lo_hi_3 = {v0WriteValidVec_res_27, v0WriteValidVec_res_26};
  wire [3:0] v0WriteValidVec_lo_3 = {v0WriteValidVec_lo_hi_3, v0WriteValidVec_lo_lo_3};
  wire [1:0] v0WriteValidVec_hi_lo_3 = {v0WriteValidVec_res_29, v0WriteValidVec_res_28};
  wire [1:0] v0WriteValidVec_hi_hi_3 = {v0WriteValidVec_res_31, v0WriteValidVec_res_30};
  wire [3:0] v0WriteValidVec_hi_3 = {v0WriteValidVec_hi_hi_3, v0WriteValidVec_hi_lo_3};
  wire [7:0] v0WriteValidVec_3 = {v0WriteValidVec_hi_3, v0WriteValidVec_lo_3};
  wire [7:0] v0WriteValidVec_lsuWriteSet_4 = lsuWriteV0_4_valid ? 8'h1 << lsuWriteV0_4_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_4 = v0WriteValidVec_v0WriteIssue_4 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_32;
  reg        v0WriteValidVec_res_33;
  reg        v0WriteValidVec_res_34;
  reg        v0WriteValidVec_res_35;
  reg        v0WriteValidVec_res_36;
  reg        v0WriteValidVec_res_37;
  reg        v0WriteValidVec_res_38;
  reg        v0WriteValidVec_res_39;
  wire [1:0] v0WriteValidVec_lo_lo_4 = {v0WriteValidVec_res_33, v0WriteValidVec_res_32};
  wire [1:0] v0WriteValidVec_lo_hi_4 = {v0WriteValidVec_res_35, v0WriteValidVec_res_34};
  wire [3:0] v0WriteValidVec_lo_4 = {v0WriteValidVec_lo_hi_4, v0WriteValidVec_lo_lo_4};
  wire [1:0] v0WriteValidVec_hi_lo_4 = {v0WriteValidVec_res_37, v0WriteValidVec_res_36};
  wire [1:0] v0WriteValidVec_hi_hi_4 = {v0WriteValidVec_res_39, v0WriteValidVec_res_38};
  wire [3:0] v0WriteValidVec_hi_4 = {v0WriteValidVec_hi_hi_4, v0WriteValidVec_hi_lo_4};
  wire [7:0] v0WriteValidVec_4 = {v0WriteValidVec_hi_4, v0WriteValidVec_lo_4};
  wire [7:0] v0WriteValidVec_lsuWriteSet_5 = lsuWriteV0_5_valid ? 8'h1 << lsuWriteV0_5_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_5 = v0WriteValidVec_v0WriteIssue_5 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_40;
  reg        v0WriteValidVec_res_41;
  reg        v0WriteValidVec_res_42;
  reg        v0WriteValidVec_res_43;
  reg        v0WriteValidVec_res_44;
  reg        v0WriteValidVec_res_45;
  reg        v0WriteValidVec_res_46;
  reg        v0WriteValidVec_res_47;
  wire [1:0] v0WriteValidVec_lo_lo_5 = {v0WriteValidVec_res_41, v0WriteValidVec_res_40};
  wire [1:0] v0WriteValidVec_lo_hi_5 = {v0WriteValidVec_res_43, v0WriteValidVec_res_42};
  wire [3:0] v0WriteValidVec_lo_5 = {v0WriteValidVec_lo_hi_5, v0WriteValidVec_lo_lo_5};
  wire [1:0] v0WriteValidVec_hi_lo_5 = {v0WriteValidVec_res_45, v0WriteValidVec_res_44};
  wire [1:0] v0WriteValidVec_hi_hi_5 = {v0WriteValidVec_res_47, v0WriteValidVec_res_46};
  wire [3:0] v0WriteValidVec_hi_5 = {v0WriteValidVec_hi_hi_5, v0WriteValidVec_hi_lo_5};
  wire [7:0] v0WriteValidVec_5 = {v0WriteValidVec_hi_5, v0WriteValidVec_lo_5};
  wire [7:0] v0WriteValidVec_lsuWriteSet_6 = lsuWriteV0_6_valid ? 8'h1 << lsuWriteV0_6_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_6 = v0WriteValidVec_v0WriteIssue_6 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_48;
  reg        v0WriteValidVec_res_49;
  reg        v0WriteValidVec_res_50;
  reg        v0WriteValidVec_res_51;
  reg        v0WriteValidVec_res_52;
  reg        v0WriteValidVec_res_53;
  reg        v0WriteValidVec_res_54;
  reg        v0WriteValidVec_res_55;
  wire [1:0] v0WriteValidVec_lo_lo_6 = {v0WriteValidVec_res_49, v0WriteValidVec_res_48};
  wire [1:0] v0WriteValidVec_lo_hi_6 = {v0WriteValidVec_res_51, v0WriteValidVec_res_50};
  wire [3:0] v0WriteValidVec_lo_6 = {v0WriteValidVec_lo_hi_6, v0WriteValidVec_lo_lo_6};
  wire [1:0] v0WriteValidVec_hi_lo_6 = {v0WriteValidVec_res_53, v0WriteValidVec_res_52};
  wire [1:0] v0WriteValidVec_hi_hi_6 = {v0WriteValidVec_res_55, v0WriteValidVec_res_54};
  wire [3:0] v0WriteValidVec_hi_6 = {v0WriteValidVec_hi_hi_6, v0WriteValidVec_hi_lo_6};
  wire [7:0] v0WriteValidVec_6 = {v0WriteValidVec_hi_6, v0WriteValidVec_lo_6};
  wire [7:0] v0WriteValidVec_lsuWriteSet_7 = lsuWriteV0_7_valid ? 8'h1 << lsuWriteV0_7_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_7 = v0WriteValidVec_v0WriteIssue_7 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_56;
  reg        v0WriteValidVec_res_57;
  reg        v0WriteValidVec_res_58;
  reg        v0WriteValidVec_res_59;
  reg        v0WriteValidVec_res_60;
  reg        v0WriteValidVec_res_61;
  reg        v0WriteValidVec_res_62;
  reg        v0WriteValidVec_res_63;
  wire [1:0] v0WriteValidVec_lo_lo_7 = {v0WriteValidVec_res_57, v0WriteValidVec_res_56};
  wire [1:0] v0WriteValidVec_lo_hi_7 = {v0WriteValidVec_res_59, v0WriteValidVec_res_58};
  wire [3:0] v0WriteValidVec_lo_7 = {v0WriteValidVec_lo_hi_7, v0WriteValidVec_lo_lo_7};
  wire [1:0] v0WriteValidVec_hi_lo_7 = {v0WriteValidVec_res_61, v0WriteValidVec_res_60};
  wire [1:0] v0WriteValidVec_hi_hi_7 = {v0WriteValidVec_res_63, v0WriteValidVec_res_62};
  wire [3:0] v0WriteValidVec_hi_7 = {v0WriteValidVec_hi_hi_7, v0WriteValidVec_hi_lo_7};
  wire [7:0] v0WriteValidVec_7 = {v0WriteValidVec_hi_7, v0WriteValidVec_lo_7};
  wire [7:0] v0WriteValidVec_lsuWriteSet_8 = lsuWriteV0_8_valid ? 8'h1 << lsuWriteV0_8_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_8 = v0WriteValidVec_v0WriteIssue_8 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_64;
  reg        v0WriteValidVec_res_65;
  reg        v0WriteValidVec_res_66;
  reg        v0WriteValidVec_res_67;
  reg        v0WriteValidVec_res_68;
  reg        v0WriteValidVec_res_69;
  reg        v0WriteValidVec_res_70;
  reg        v0WriteValidVec_res_71;
  wire [1:0] v0WriteValidVec_lo_lo_8 = {v0WriteValidVec_res_65, v0WriteValidVec_res_64};
  wire [1:0] v0WriteValidVec_lo_hi_8 = {v0WriteValidVec_res_67, v0WriteValidVec_res_66};
  wire [3:0] v0WriteValidVec_lo_8 = {v0WriteValidVec_lo_hi_8, v0WriteValidVec_lo_lo_8};
  wire [1:0] v0WriteValidVec_hi_lo_8 = {v0WriteValidVec_res_69, v0WriteValidVec_res_68};
  wire [1:0] v0WriteValidVec_hi_hi_8 = {v0WriteValidVec_res_71, v0WriteValidVec_res_70};
  wire [3:0] v0WriteValidVec_hi_8 = {v0WriteValidVec_hi_hi_8, v0WriteValidVec_hi_lo_8};
  wire [7:0] v0WriteValidVec_8 = {v0WriteValidVec_hi_8, v0WriteValidVec_lo_8};
  wire [7:0] v0WriteValidVec_lsuWriteSet_9 = lsuWriteV0_9_valid ? 8'h1 << lsuWriteV0_9_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_9 = v0WriteValidVec_v0WriteIssue_9 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_72;
  reg        v0WriteValidVec_res_73;
  reg        v0WriteValidVec_res_74;
  reg        v0WriteValidVec_res_75;
  reg        v0WriteValidVec_res_76;
  reg        v0WriteValidVec_res_77;
  reg        v0WriteValidVec_res_78;
  reg        v0WriteValidVec_res_79;
  wire [1:0] v0WriteValidVec_lo_lo_9 = {v0WriteValidVec_res_73, v0WriteValidVec_res_72};
  wire [1:0] v0WriteValidVec_lo_hi_9 = {v0WriteValidVec_res_75, v0WriteValidVec_res_74};
  wire [3:0] v0WriteValidVec_lo_9 = {v0WriteValidVec_lo_hi_9, v0WriteValidVec_lo_lo_9};
  wire [1:0] v0WriteValidVec_hi_lo_9 = {v0WriteValidVec_res_77, v0WriteValidVec_res_76};
  wire [1:0] v0WriteValidVec_hi_hi_9 = {v0WriteValidVec_res_79, v0WriteValidVec_res_78};
  wire [3:0] v0WriteValidVec_hi_9 = {v0WriteValidVec_hi_hi_9, v0WriteValidVec_hi_lo_9};
  wire [7:0] v0WriteValidVec_9 = {v0WriteValidVec_hi_9, v0WriteValidVec_lo_9};
  wire [7:0] v0WriteValidVec_lsuWriteSet_10 = lsuWriteV0_10_valid ? 8'h1 << lsuWriteV0_10_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_10 = v0WriteValidVec_v0WriteIssue_10 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_80;
  reg        v0WriteValidVec_res_81;
  reg        v0WriteValidVec_res_82;
  reg        v0WriteValidVec_res_83;
  reg        v0WriteValidVec_res_84;
  reg        v0WriteValidVec_res_85;
  reg        v0WriteValidVec_res_86;
  reg        v0WriteValidVec_res_87;
  wire [1:0] v0WriteValidVec_lo_lo_10 = {v0WriteValidVec_res_81, v0WriteValidVec_res_80};
  wire [1:0] v0WriteValidVec_lo_hi_10 = {v0WriteValidVec_res_83, v0WriteValidVec_res_82};
  wire [3:0] v0WriteValidVec_lo_10 = {v0WriteValidVec_lo_hi_10, v0WriteValidVec_lo_lo_10};
  wire [1:0] v0WriteValidVec_hi_lo_10 = {v0WriteValidVec_res_85, v0WriteValidVec_res_84};
  wire [1:0] v0WriteValidVec_hi_hi_10 = {v0WriteValidVec_res_87, v0WriteValidVec_res_86};
  wire [3:0] v0WriteValidVec_hi_10 = {v0WriteValidVec_hi_hi_10, v0WriteValidVec_hi_lo_10};
  wire [7:0] v0WriteValidVec_10 = {v0WriteValidVec_hi_10, v0WriteValidVec_lo_10};
  wire [7:0] v0WriteValidVec_lsuWriteSet_11 = lsuWriteV0_11_valid ? 8'h1 << lsuWriteV0_11_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_11 = v0WriteValidVec_v0WriteIssue_11 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_88;
  reg        v0WriteValidVec_res_89;
  reg        v0WriteValidVec_res_90;
  reg        v0WriteValidVec_res_91;
  reg        v0WriteValidVec_res_92;
  reg        v0WriteValidVec_res_93;
  reg        v0WriteValidVec_res_94;
  reg        v0WriteValidVec_res_95;
  wire [1:0] v0WriteValidVec_lo_lo_11 = {v0WriteValidVec_res_89, v0WriteValidVec_res_88};
  wire [1:0] v0WriteValidVec_lo_hi_11 = {v0WriteValidVec_res_91, v0WriteValidVec_res_90};
  wire [3:0] v0WriteValidVec_lo_11 = {v0WriteValidVec_lo_hi_11, v0WriteValidVec_lo_lo_11};
  wire [1:0] v0WriteValidVec_hi_lo_11 = {v0WriteValidVec_res_93, v0WriteValidVec_res_92};
  wire [1:0] v0WriteValidVec_hi_hi_11 = {v0WriteValidVec_res_95, v0WriteValidVec_res_94};
  wire [3:0] v0WriteValidVec_hi_11 = {v0WriteValidVec_hi_hi_11, v0WriteValidVec_hi_lo_11};
  wire [7:0] v0WriteValidVec_11 = {v0WriteValidVec_hi_11, v0WriteValidVec_lo_11};
  wire [7:0] v0WriteValidVec_lsuWriteSet_12 = lsuWriteV0_12_valid ? 8'h1 << lsuWriteV0_12_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_12 = v0WriteValidVec_v0WriteIssue_12 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_96;
  reg        v0WriteValidVec_res_97;
  reg        v0WriteValidVec_res_98;
  reg        v0WriteValidVec_res_99;
  reg        v0WriteValidVec_res_100;
  reg        v0WriteValidVec_res_101;
  reg        v0WriteValidVec_res_102;
  reg        v0WriteValidVec_res_103;
  wire [1:0] v0WriteValidVec_lo_lo_12 = {v0WriteValidVec_res_97, v0WriteValidVec_res_96};
  wire [1:0] v0WriteValidVec_lo_hi_12 = {v0WriteValidVec_res_99, v0WriteValidVec_res_98};
  wire [3:0] v0WriteValidVec_lo_12 = {v0WriteValidVec_lo_hi_12, v0WriteValidVec_lo_lo_12};
  wire [1:0] v0WriteValidVec_hi_lo_12 = {v0WriteValidVec_res_101, v0WriteValidVec_res_100};
  wire [1:0] v0WriteValidVec_hi_hi_12 = {v0WriteValidVec_res_103, v0WriteValidVec_res_102};
  wire [3:0] v0WriteValidVec_hi_12 = {v0WriteValidVec_hi_hi_12, v0WriteValidVec_hi_lo_12};
  wire [7:0] v0WriteValidVec_12 = {v0WriteValidVec_hi_12, v0WriteValidVec_lo_12};
  wire [7:0] v0WriteValidVec_lsuWriteSet_13 = lsuWriteV0_13_valid ? 8'h1 << lsuWriteV0_13_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_13 = v0WriteValidVec_v0WriteIssue_13 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_104;
  reg        v0WriteValidVec_res_105;
  reg        v0WriteValidVec_res_106;
  reg        v0WriteValidVec_res_107;
  reg        v0WriteValidVec_res_108;
  reg        v0WriteValidVec_res_109;
  reg        v0WriteValidVec_res_110;
  reg        v0WriteValidVec_res_111;
  wire [1:0] v0WriteValidVec_lo_lo_13 = {v0WriteValidVec_res_105, v0WriteValidVec_res_104};
  wire [1:0] v0WriteValidVec_lo_hi_13 = {v0WriteValidVec_res_107, v0WriteValidVec_res_106};
  wire [3:0] v0WriteValidVec_lo_13 = {v0WriteValidVec_lo_hi_13, v0WriteValidVec_lo_lo_13};
  wire [1:0] v0WriteValidVec_hi_lo_13 = {v0WriteValidVec_res_109, v0WriteValidVec_res_108};
  wire [1:0] v0WriteValidVec_hi_hi_13 = {v0WriteValidVec_res_111, v0WriteValidVec_res_110};
  wire [3:0] v0WriteValidVec_hi_13 = {v0WriteValidVec_hi_hi_13, v0WriteValidVec_hi_lo_13};
  wire [7:0] v0WriteValidVec_13 = {v0WriteValidVec_hi_13, v0WriteValidVec_lo_13};
  wire [7:0] v0WriteValidVec_lsuWriteSet_14 = lsuWriteV0_14_valid ? 8'h1 << lsuWriteV0_14_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_14 = v0WriteValidVec_v0WriteIssue_14 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_112;
  reg        v0WriteValidVec_res_113;
  reg        v0WriteValidVec_res_114;
  reg        v0WriteValidVec_res_115;
  reg        v0WriteValidVec_res_116;
  reg        v0WriteValidVec_res_117;
  reg        v0WriteValidVec_res_118;
  reg        v0WriteValidVec_res_119;
  wire [1:0] v0WriteValidVec_lo_lo_14 = {v0WriteValidVec_res_113, v0WriteValidVec_res_112};
  wire [1:0] v0WriteValidVec_lo_hi_14 = {v0WriteValidVec_res_115, v0WriteValidVec_res_114};
  wire [3:0] v0WriteValidVec_lo_14 = {v0WriteValidVec_lo_hi_14, v0WriteValidVec_lo_lo_14};
  wire [1:0] v0WriteValidVec_hi_lo_14 = {v0WriteValidVec_res_117, v0WriteValidVec_res_116};
  wire [1:0] v0WriteValidVec_hi_hi_14 = {v0WriteValidVec_res_119, v0WriteValidVec_res_118};
  wire [3:0] v0WriteValidVec_hi_14 = {v0WriteValidVec_hi_hi_14, v0WriteValidVec_hi_lo_14};
  wire [7:0] v0WriteValidVec_14 = {v0WriteValidVec_hi_14, v0WriteValidVec_lo_14};
  wire [7:0] v0WriteValidVec_lsuWriteSet_15 = lsuWriteV0_15_valid ? 8'h1 << lsuWriteV0_15_bits : 8'h0;
  wire [7:0] v0WriteValidVec_updateOH_15 = v0WriteValidVec_v0WriteIssue_15 ? issueIndex1H : 8'h0;
  reg        v0WriteValidVec_res_120;
  reg        v0WriteValidVec_res_121;
  reg        v0WriteValidVec_res_122;
  reg        v0WriteValidVec_res_123;
  reg        v0WriteValidVec_res_124;
  reg        v0WriteValidVec_res_125;
  reg        v0WriteValidVec_res_126;
  reg        v0WriteValidVec_res_127;
  wire [1:0] v0WriteValidVec_lo_lo_15 = {v0WriteValidVec_res_121, v0WriteValidVec_res_120};
  wire [1:0] v0WriteValidVec_lo_hi_15 = {v0WriteValidVec_res_123, v0WriteValidVec_res_122};
  wire [3:0] v0WriteValidVec_lo_15 = {v0WriteValidVec_lo_hi_15, v0WriteValidVec_lo_lo_15};
  wire [1:0] v0WriteValidVec_hi_lo_15 = {v0WriteValidVec_res_125, v0WriteValidVec_res_124};
  wire [1:0] v0WriteValidVec_hi_hi_15 = {v0WriteValidVec_res_127, v0WriteValidVec_res_126};
  wire [3:0] v0WriteValidVec_hi_15 = {v0WriteValidVec_hi_hi_15, v0WriteValidVec_hi_lo_15};
  wire [7:0] v0WriteValidVec_15 = {v0WriteValidVec_hi_15, v0WriteValidVec_lo_15};
  wire       _GEN_0 = instructionIssue_valid & instructionIssue_bits_useV0AsMask & instructionIssue_bits_toLane;
  wire       useV0AsMaskToken_useV0Issue;
  assign useV0AsMaskToken_useV0Issue = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_1;
  assign useV0AsMaskToken_useV0Issue_1 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_2;
  assign useV0AsMaskToken_useV0Issue_2 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_3;
  assign useV0AsMaskToken_useV0Issue_3 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_4;
  assign useV0AsMaskToken_useV0Issue_4 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_5;
  assign useV0AsMaskToken_useV0Issue_5 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_6;
  assign useV0AsMaskToken_useV0Issue_6 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_7;
  assign useV0AsMaskToken_useV0Issue_7 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_8;
  assign useV0AsMaskToken_useV0Issue_8 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_9;
  assign useV0AsMaskToken_useV0Issue_9 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_10;
  assign useV0AsMaskToken_useV0Issue_10 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_11;
  assign useV0AsMaskToken_useV0Issue_11 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_12;
  assign useV0AsMaskToken_useV0Issue_12 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_13;
  assign useV0AsMaskToken_useV0Issue_13 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_14;
  assign useV0AsMaskToken_useV0Issue_14 = _GEN_0;
  wire       useV0AsMaskToken_useV0Issue_15;
  assign useV0AsMaskToken_useV0Issue_15 = _GEN_0;
  wire [7:0] useV0AsMaskToken_updateOH = useV0AsMaskToken_useV0Issue ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res;
  reg        useV0AsMaskToken_res_1;
  reg        useV0AsMaskToken_res_2;
  reg        useV0AsMaskToken_res_3;
  reg        useV0AsMaskToken_res_4;
  reg        useV0AsMaskToken_res_5;
  reg        useV0AsMaskToken_res_6;
  reg        useV0AsMaskToken_res_7;
  wire [1:0] useV0AsMaskToken_lo_lo = {useV0AsMaskToken_res_1, useV0AsMaskToken_res};
  wire [1:0] useV0AsMaskToken_lo_hi = {useV0AsMaskToken_res_3, useV0AsMaskToken_res_2};
  wire [3:0] useV0AsMaskToken_lo = {useV0AsMaskToken_lo_hi, useV0AsMaskToken_lo_lo};
  wire [1:0] useV0AsMaskToken_hi_lo = {useV0AsMaskToken_res_5, useV0AsMaskToken_res_4};
  wire [1:0] useV0AsMaskToken_hi_hi = {useV0AsMaskToken_res_7, useV0AsMaskToken_res_6};
  wire [3:0] useV0AsMaskToken_hi = {useV0AsMaskToken_hi_hi, useV0AsMaskToken_hi_lo};
  wire [7:0] useV0AsMaskToken_updateOH_1 = useV0AsMaskToken_useV0Issue_1 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_8;
  reg        useV0AsMaskToken_res_9;
  reg        useV0AsMaskToken_res_10;
  reg        useV0AsMaskToken_res_11;
  reg        useV0AsMaskToken_res_12;
  reg        useV0AsMaskToken_res_13;
  reg        useV0AsMaskToken_res_14;
  reg        useV0AsMaskToken_res_15;
  wire [1:0] useV0AsMaskToken_lo_lo_1 = {useV0AsMaskToken_res_9, useV0AsMaskToken_res_8};
  wire [1:0] useV0AsMaskToken_lo_hi_1 = {useV0AsMaskToken_res_11, useV0AsMaskToken_res_10};
  wire [3:0] useV0AsMaskToken_lo_1 = {useV0AsMaskToken_lo_hi_1, useV0AsMaskToken_lo_lo_1};
  wire [1:0] useV0AsMaskToken_hi_lo_1 = {useV0AsMaskToken_res_13, useV0AsMaskToken_res_12};
  wire [1:0] useV0AsMaskToken_hi_hi_1 = {useV0AsMaskToken_res_15, useV0AsMaskToken_res_14};
  wire [3:0] useV0AsMaskToken_hi_1 = {useV0AsMaskToken_hi_hi_1, useV0AsMaskToken_hi_lo_1};
  wire [7:0] useV0AsMaskToken_updateOH_2 = useV0AsMaskToken_useV0Issue_2 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_16;
  reg        useV0AsMaskToken_res_17;
  reg        useV0AsMaskToken_res_18;
  reg        useV0AsMaskToken_res_19;
  reg        useV0AsMaskToken_res_20;
  reg        useV0AsMaskToken_res_21;
  reg        useV0AsMaskToken_res_22;
  reg        useV0AsMaskToken_res_23;
  wire [1:0] useV0AsMaskToken_lo_lo_2 = {useV0AsMaskToken_res_17, useV0AsMaskToken_res_16};
  wire [1:0] useV0AsMaskToken_lo_hi_2 = {useV0AsMaskToken_res_19, useV0AsMaskToken_res_18};
  wire [3:0] useV0AsMaskToken_lo_2 = {useV0AsMaskToken_lo_hi_2, useV0AsMaskToken_lo_lo_2};
  wire [1:0] useV0AsMaskToken_hi_lo_2 = {useV0AsMaskToken_res_21, useV0AsMaskToken_res_20};
  wire [1:0] useV0AsMaskToken_hi_hi_2 = {useV0AsMaskToken_res_23, useV0AsMaskToken_res_22};
  wire [3:0] useV0AsMaskToken_hi_2 = {useV0AsMaskToken_hi_hi_2, useV0AsMaskToken_hi_lo_2};
  wire [7:0] useV0AsMaskToken_updateOH_3 = useV0AsMaskToken_useV0Issue_3 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_24;
  reg        useV0AsMaskToken_res_25;
  reg        useV0AsMaskToken_res_26;
  reg        useV0AsMaskToken_res_27;
  reg        useV0AsMaskToken_res_28;
  reg        useV0AsMaskToken_res_29;
  reg        useV0AsMaskToken_res_30;
  reg        useV0AsMaskToken_res_31;
  wire [1:0] useV0AsMaskToken_lo_lo_3 = {useV0AsMaskToken_res_25, useV0AsMaskToken_res_24};
  wire [1:0] useV0AsMaskToken_lo_hi_3 = {useV0AsMaskToken_res_27, useV0AsMaskToken_res_26};
  wire [3:0] useV0AsMaskToken_lo_3 = {useV0AsMaskToken_lo_hi_3, useV0AsMaskToken_lo_lo_3};
  wire [1:0] useV0AsMaskToken_hi_lo_3 = {useV0AsMaskToken_res_29, useV0AsMaskToken_res_28};
  wire [1:0] useV0AsMaskToken_hi_hi_3 = {useV0AsMaskToken_res_31, useV0AsMaskToken_res_30};
  wire [3:0] useV0AsMaskToken_hi_3 = {useV0AsMaskToken_hi_hi_3, useV0AsMaskToken_hi_lo_3};
  wire [7:0] useV0AsMaskToken_updateOH_4 = useV0AsMaskToken_useV0Issue_4 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_32;
  reg        useV0AsMaskToken_res_33;
  reg        useV0AsMaskToken_res_34;
  reg        useV0AsMaskToken_res_35;
  reg        useV0AsMaskToken_res_36;
  reg        useV0AsMaskToken_res_37;
  reg        useV0AsMaskToken_res_38;
  reg        useV0AsMaskToken_res_39;
  wire [1:0] useV0AsMaskToken_lo_lo_4 = {useV0AsMaskToken_res_33, useV0AsMaskToken_res_32};
  wire [1:0] useV0AsMaskToken_lo_hi_4 = {useV0AsMaskToken_res_35, useV0AsMaskToken_res_34};
  wire [3:0] useV0AsMaskToken_lo_4 = {useV0AsMaskToken_lo_hi_4, useV0AsMaskToken_lo_lo_4};
  wire [1:0] useV0AsMaskToken_hi_lo_4 = {useV0AsMaskToken_res_37, useV0AsMaskToken_res_36};
  wire [1:0] useV0AsMaskToken_hi_hi_4 = {useV0AsMaskToken_res_39, useV0AsMaskToken_res_38};
  wire [3:0] useV0AsMaskToken_hi_4 = {useV0AsMaskToken_hi_hi_4, useV0AsMaskToken_hi_lo_4};
  wire [7:0] useV0AsMaskToken_updateOH_5 = useV0AsMaskToken_useV0Issue_5 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_40;
  reg        useV0AsMaskToken_res_41;
  reg        useV0AsMaskToken_res_42;
  reg        useV0AsMaskToken_res_43;
  reg        useV0AsMaskToken_res_44;
  reg        useV0AsMaskToken_res_45;
  reg        useV0AsMaskToken_res_46;
  reg        useV0AsMaskToken_res_47;
  wire [1:0] useV0AsMaskToken_lo_lo_5 = {useV0AsMaskToken_res_41, useV0AsMaskToken_res_40};
  wire [1:0] useV0AsMaskToken_lo_hi_5 = {useV0AsMaskToken_res_43, useV0AsMaskToken_res_42};
  wire [3:0] useV0AsMaskToken_lo_5 = {useV0AsMaskToken_lo_hi_5, useV0AsMaskToken_lo_lo_5};
  wire [1:0] useV0AsMaskToken_hi_lo_5 = {useV0AsMaskToken_res_45, useV0AsMaskToken_res_44};
  wire [1:0] useV0AsMaskToken_hi_hi_5 = {useV0AsMaskToken_res_47, useV0AsMaskToken_res_46};
  wire [3:0] useV0AsMaskToken_hi_5 = {useV0AsMaskToken_hi_hi_5, useV0AsMaskToken_hi_lo_5};
  wire [7:0] useV0AsMaskToken_updateOH_6 = useV0AsMaskToken_useV0Issue_6 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_48;
  reg        useV0AsMaskToken_res_49;
  reg        useV0AsMaskToken_res_50;
  reg        useV0AsMaskToken_res_51;
  reg        useV0AsMaskToken_res_52;
  reg        useV0AsMaskToken_res_53;
  reg        useV0AsMaskToken_res_54;
  reg        useV0AsMaskToken_res_55;
  wire [1:0] useV0AsMaskToken_lo_lo_6 = {useV0AsMaskToken_res_49, useV0AsMaskToken_res_48};
  wire [1:0] useV0AsMaskToken_lo_hi_6 = {useV0AsMaskToken_res_51, useV0AsMaskToken_res_50};
  wire [3:0] useV0AsMaskToken_lo_6 = {useV0AsMaskToken_lo_hi_6, useV0AsMaskToken_lo_lo_6};
  wire [1:0] useV0AsMaskToken_hi_lo_6 = {useV0AsMaskToken_res_53, useV0AsMaskToken_res_52};
  wire [1:0] useV0AsMaskToken_hi_hi_6 = {useV0AsMaskToken_res_55, useV0AsMaskToken_res_54};
  wire [3:0] useV0AsMaskToken_hi_6 = {useV0AsMaskToken_hi_hi_6, useV0AsMaskToken_hi_lo_6};
  wire [7:0] useV0AsMaskToken_updateOH_7 = useV0AsMaskToken_useV0Issue_7 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_56;
  reg        useV0AsMaskToken_res_57;
  reg        useV0AsMaskToken_res_58;
  reg        useV0AsMaskToken_res_59;
  reg        useV0AsMaskToken_res_60;
  reg        useV0AsMaskToken_res_61;
  reg        useV0AsMaskToken_res_62;
  reg        useV0AsMaskToken_res_63;
  wire [1:0] useV0AsMaskToken_lo_lo_7 = {useV0AsMaskToken_res_57, useV0AsMaskToken_res_56};
  wire [1:0] useV0AsMaskToken_lo_hi_7 = {useV0AsMaskToken_res_59, useV0AsMaskToken_res_58};
  wire [3:0] useV0AsMaskToken_lo_7 = {useV0AsMaskToken_lo_hi_7, useV0AsMaskToken_lo_lo_7};
  wire [1:0] useV0AsMaskToken_hi_lo_7 = {useV0AsMaskToken_res_61, useV0AsMaskToken_res_60};
  wire [1:0] useV0AsMaskToken_hi_hi_7 = {useV0AsMaskToken_res_63, useV0AsMaskToken_res_62};
  wire [3:0] useV0AsMaskToken_hi_7 = {useV0AsMaskToken_hi_hi_7, useV0AsMaskToken_hi_lo_7};
  wire [7:0] useV0AsMaskToken_updateOH_8 = useV0AsMaskToken_useV0Issue_8 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_64;
  reg        useV0AsMaskToken_res_65;
  reg        useV0AsMaskToken_res_66;
  reg        useV0AsMaskToken_res_67;
  reg        useV0AsMaskToken_res_68;
  reg        useV0AsMaskToken_res_69;
  reg        useV0AsMaskToken_res_70;
  reg        useV0AsMaskToken_res_71;
  wire [1:0] useV0AsMaskToken_lo_lo_8 = {useV0AsMaskToken_res_65, useV0AsMaskToken_res_64};
  wire [1:0] useV0AsMaskToken_lo_hi_8 = {useV0AsMaskToken_res_67, useV0AsMaskToken_res_66};
  wire [3:0] useV0AsMaskToken_lo_8 = {useV0AsMaskToken_lo_hi_8, useV0AsMaskToken_lo_lo_8};
  wire [1:0] useV0AsMaskToken_hi_lo_8 = {useV0AsMaskToken_res_69, useV0AsMaskToken_res_68};
  wire [1:0] useV0AsMaskToken_hi_hi_8 = {useV0AsMaskToken_res_71, useV0AsMaskToken_res_70};
  wire [3:0] useV0AsMaskToken_hi_8 = {useV0AsMaskToken_hi_hi_8, useV0AsMaskToken_hi_lo_8};
  wire [7:0] useV0AsMaskToken_updateOH_9 = useV0AsMaskToken_useV0Issue_9 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_72;
  reg        useV0AsMaskToken_res_73;
  reg        useV0AsMaskToken_res_74;
  reg        useV0AsMaskToken_res_75;
  reg        useV0AsMaskToken_res_76;
  reg        useV0AsMaskToken_res_77;
  reg        useV0AsMaskToken_res_78;
  reg        useV0AsMaskToken_res_79;
  wire [1:0] useV0AsMaskToken_lo_lo_9 = {useV0AsMaskToken_res_73, useV0AsMaskToken_res_72};
  wire [1:0] useV0AsMaskToken_lo_hi_9 = {useV0AsMaskToken_res_75, useV0AsMaskToken_res_74};
  wire [3:0] useV0AsMaskToken_lo_9 = {useV0AsMaskToken_lo_hi_9, useV0AsMaskToken_lo_lo_9};
  wire [1:0] useV0AsMaskToken_hi_lo_9 = {useV0AsMaskToken_res_77, useV0AsMaskToken_res_76};
  wire [1:0] useV0AsMaskToken_hi_hi_9 = {useV0AsMaskToken_res_79, useV0AsMaskToken_res_78};
  wire [3:0] useV0AsMaskToken_hi_9 = {useV0AsMaskToken_hi_hi_9, useV0AsMaskToken_hi_lo_9};
  wire [7:0] useV0AsMaskToken_updateOH_10 = useV0AsMaskToken_useV0Issue_10 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_80;
  reg        useV0AsMaskToken_res_81;
  reg        useV0AsMaskToken_res_82;
  reg        useV0AsMaskToken_res_83;
  reg        useV0AsMaskToken_res_84;
  reg        useV0AsMaskToken_res_85;
  reg        useV0AsMaskToken_res_86;
  reg        useV0AsMaskToken_res_87;
  wire [1:0] useV0AsMaskToken_lo_lo_10 = {useV0AsMaskToken_res_81, useV0AsMaskToken_res_80};
  wire [1:0] useV0AsMaskToken_lo_hi_10 = {useV0AsMaskToken_res_83, useV0AsMaskToken_res_82};
  wire [3:0] useV0AsMaskToken_lo_10 = {useV0AsMaskToken_lo_hi_10, useV0AsMaskToken_lo_lo_10};
  wire [1:0] useV0AsMaskToken_hi_lo_10 = {useV0AsMaskToken_res_85, useV0AsMaskToken_res_84};
  wire [1:0] useV0AsMaskToken_hi_hi_10 = {useV0AsMaskToken_res_87, useV0AsMaskToken_res_86};
  wire [3:0] useV0AsMaskToken_hi_10 = {useV0AsMaskToken_hi_hi_10, useV0AsMaskToken_hi_lo_10};
  wire [7:0] useV0AsMaskToken_updateOH_11 = useV0AsMaskToken_useV0Issue_11 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_88;
  reg        useV0AsMaskToken_res_89;
  reg        useV0AsMaskToken_res_90;
  reg        useV0AsMaskToken_res_91;
  reg        useV0AsMaskToken_res_92;
  reg        useV0AsMaskToken_res_93;
  reg        useV0AsMaskToken_res_94;
  reg        useV0AsMaskToken_res_95;
  wire [1:0] useV0AsMaskToken_lo_lo_11 = {useV0AsMaskToken_res_89, useV0AsMaskToken_res_88};
  wire [1:0] useV0AsMaskToken_lo_hi_11 = {useV0AsMaskToken_res_91, useV0AsMaskToken_res_90};
  wire [3:0] useV0AsMaskToken_lo_11 = {useV0AsMaskToken_lo_hi_11, useV0AsMaskToken_lo_lo_11};
  wire [1:0] useV0AsMaskToken_hi_lo_11 = {useV0AsMaskToken_res_93, useV0AsMaskToken_res_92};
  wire [1:0] useV0AsMaskToken_hi_hi_11 = {useV0AsMaskToken_res_95, useV0AsMaskToken_res_94};
  wire [3:0] useV0AsMaskToken_hi_11 = {useV0AsMaskToken_hi_hi_11, useV0AsMaskToken_hi_lo_11};
  wire [7:0] useV0AsMaskToken_updateOH_12 = useV0AsMaskToken_useV0Issue_12 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_96;
  reg        useV0AsMaskToken_res_97;
  reg        useV0AsMaskToken_res_98;
  reg        useV0AsMaskToken_res_99;
  reg        useV0AsMaskToken_res_100;
  reg        useV0AsMaskToken_res_101;
  reg        useV0AsMaskToken_res_102;
  reg        useV0AsMaskToken_res_103;
  wire [1:0] useV0AsMaskToken_lo_lo_12 = {useV0AsMaskToken_res_97, useV0AsMaskToken_res_96};
  wire [1:0] useV0AsMaskToken_lo_hi_12 = {useV0AsMaskToken_res_99, useV0AsMaskToken_res_98};
  wire [3:0] useV0AsMaskToken_lo_12 = {useV0AsMaskToken_lo_hi_12, useV0AsMaskToken_lo_lo_12};
  wire [1:0] useV0AsMaskToken_hi_lo_12 = {useV0AsMaskToken_res_101, useV0AsMaskToken_res_100};
  wire [1:0] useV0AsMaskToken_hi_hi_12 = {useV0AsMaskToken_res_103, useV0AsMaskToken_res_102};
  wire [3:0] useV0AsMaskToken_hi_12 = {useV0AsMaskToken_hi_hi_12, useV0AsMaskToken_hi_lo_12};
  wire [7:0] useV0AsMaskToken_updateOH_13 = useV0AsMaskToken_useV0Issue_13 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_104;
  reg        useV0AsMaskToken_res_105;
  reg        useV0AsMaskToken_res_106;
  reg        useV0AsMaskToken_res_107;
  reg        useV0AsMaskToken_res_108;
  reg        useV0AsMaskToken_res_109;
  reg        useV0AsMaskToken_res_110;
  reg        useV0AsMaskToken_res_111;
  wire [1:0] useV0AsMaskToken_lo_lo_13 = {useV0AsMaskToken_res_105, useV0AsMaskToken_res_104};
  wire [1:0] useV0AsMaskToken_lo_hi_13 = {useV0AsMaskToken_res_107, useV0AsMaskToken_res_106};
  wire [3:0] useV0AsMaskToken_lo_13 = {useV0AsMaskToken_lo_hi_13, useV0AsMaskToken_lo_lo_13};
  wire [1:0] useV0AsMaskToken_hi_lo_13 = {useV0AsMaskToken_res_109, useV0AsMaskToken_res_108};
  wire [1:0] useV0AsMaskToken_hi_hi_13 = {useV0AsMaskToken_res_111, useV0AsMaskToken_res_110};
  wire [3:0] useV0AsMaskToken_hi_13 = {useV0AsMaskToken_hi_hi_13, useV0AsMaskToken_hi_lo_13};
  wire [7:0] useV0AsMaskToken_updateOH_14 = useV0AsMaskToken_useV0Issue_14 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_112;
  reg        useV0AsMaskToken_res_113;
  reg        useV0AsMaskToken_res_114;
  reg        useV0AsMaskToken_res_115;
  reg        useV0AsMaskToken_res_116;
  reg        useV0AsMaskToken_res_117;
  reg        useV0AsMaskToken_res_118;
  reg        useV0AsMaskToken_res_119;
  wire [1:0] useV0AsMaskToken_lo_lo_14 = {useV0AsMaskToken_res_113, useV0AsMaskToken_res_112};
  wire [1:0] useV0AsMaskToken_lo_hi_14 = {useV0AsMaskToken_res_115, useV0AsMaskToken_res_114};
  wire [3:0] useV0AsMaskToken_lo_14 = {useV0AsMaskToken_lo_hi_14, useV0AsMaskToken_lo_lo_14};
  wire [1:0] useV0AsMaskToken_hi_lo_14 = {useV0AsMaskToken_res_117, useV0AsMaskToken_res_116};
  wire [1:0] useV0AsMaskToken_hi_hi_14 = {useV0AsMaskToken_res_119, useV0AsMaskToken_res_118};
  wire [3:0] useV0AsMaskToken_hi_14 = {useV0AsMaskToken_hi_hi_14, useV0AsMaskToken_hi_lo_14};
  wire [7:0] useV0AsMaskToken_updateOH_15 = useV0AsMaskToken_useV0Issue_15 ? issueIndex1H : 8'h0;
  reg        useV0AsMaskToken_res_120;
  reg        useV0AsMaskToken_res_121;
  reg        useV0AsMaskToken_res_122;
  reg        useV0AsMaskToken_res_123;
  reg        useV0AsMaskToken_res_124;
  reg        useV0AsMaskToken_res_125;
  reg        useV0AsMaskToken_res_126;
  reg        useV0AsMaskToken_res_127;
  wire [1:0] useV0AsMaskToken_lo_lo_15 = {useV0AsMaskToken_res_121, useV0AsMaskToken_res_120};
  wire [1:0] useV0AsMaskToken_lo_hi_15 = {useV0AsMaskToken_res_123, useV0AsMaskToken_res_122};
  wire [3:0] useV0AsMaskToken_lo_15 = {useV0AsMaskToken_lo_hi_15, useV0AsMaskToken_lo_lo_15};
  wire [1:0] useV0AsMaskToken_hi_lo_15 = {useV0AsMaskToken_res_125, useV0AsMaskToken_res_124};
  wire [1:0] useV0AsMaskToken_hi_hi_15 = {useV0AsMaskToken_res_127, useV0AsMaskToken_res_126};
  wire [3:0] useV0AsMaskToken_hi_15 = {useV0AsMaskToken_hi_hi_15, useV0AsMaskToken_hi_lo_15};
  wire [7:0] useV0AsMaskToken =
    {useV0AsMaskToken_hi, useV0AsMaskToken_lo} | {useV0AsMaskToken_hi_1, useV0AsMaskToken_lo_1} | {useV0AsMaskToken_hi_2, useV0AsMaskToken_lo_2} | {useV0AsMaskToken_hi_3, useV0AsMaskToken_lo_3}
    | {useV0AsMaskToken_hi_4, useV0AsMaskToken_lo_4} | {useV0AsMaskToken_hi_5, useV0AsMaskToken_lo_5} | {useV0AsMaskToken_hi_6, useV0AsMaskToken_lo_6} | {useV0AsMaskToken_hi_7, useV0AsMaskToken_lo_7}
    | {useV0AsMaskToken_hi_8, useV0AsMaskToken_lo_8} | {useV0AsMaskToken_hi_9, useV0AsMaskToken_lo_9} | {useV0AsMaskToken_hi_10, useV0AsMaskToken_lo_10} | {useV0AsMaskToken_hi_11, useV0AsMaskToken_lo_11}
    | {useV0AsMaskToken_hi_12, useV0AsMaskToken_lo_12} | {useV0AsMaskToken_hi_13, useV0AsMaskToken_lo_13} | {useV0AsMaskToken_hi_14, useV0AsMaskToken_lo_14} | {useV0AsMaskToken_hi_15, useV0AsMaskToken_lo_15};
  wire       maskUnitWriteV0_set = _maskUnitWriteV0_set_T & instructionIssue_bits_toMask;
  reg        maskUnitWriteV0;
  wire [7:0] _v0WriteValid_output =
    v0WriteValidVec_0 | v0WriteValidVec_1 | v0WriteValidVec_2 | v0WriteValidVec_3 | v0WriteValidVec_4 | v0WriteValidVec_5 | v0WriteValidVec_6 | v0WriteValidVec_7 | v0WriteValidVec_8 | v0WriteValidVec_9 | v0WriteValidVec_10
    | v0WriteValidVec_11 | v0WriteValidVec_12 | v0WriteValidVec_13 | v0WriteValidVec_14 | v0WriteValidVec_15;
  wire       v0Conflict = instructionIssue_bits_writeV0 & (|useV0AsMaskToken) | instructionIssue_bits_useV0AsMask & ((|_v0WriteValid_output) | maskUnitWriteV0);
  always @(posedge clock) begin
    if (reset) begin
      v0WriteValidVec_res <= 1'h0;
      v0WriteValidVec_res_1 <= 1'h0;
      v0WriteValidVec_res_2 <= 1'h0;
      v0WriteValidVec_res_3 <= 1'h0;
      v0WriteValidVec_res_4 <= 1'h0;
      v0WriteValidVec_res_5 <= 1'h0;
      v0WriteValidVec_res_6 <= 1'h0;
      v0WriteValidVec_res_7 <= 1'h0;
      v0WriteValidVec_res_8 <= 1'h0;
      v0WriteValidVec_res_9 <= 1'h0;
      v0WriteValidVec_res_10 <= 1'h0;
      v0WriteValidVec_res_11 <= 1'h0;
      v0WriteValidVec_res_12 <= 1'h0;
      v0WriteValidVec_res_13 <= 1'h0;
      v0WriteValidVec_res_14 <= 1'h0;
      v0WriteValidVec_res_15 <= 1'h0;
      v0WriteValidVec_res_16 <= 1'h0;
      v0WriteValidVec_res_17 <= 1'h0;
      v0WriteValidVec_res_18 <= 1'h0;
      v0WriteValidVec_res_19 <= 1'h0;
      v0WriteValidVec_res_20 <= 1'h0;
      v0WriteValidVec_res_21 <= 1'h0;
      v0WriteValidVec_res_22 <= 1'h0;
      v0WriteValidVec_res_23 <= 1'h0;
      v0WriteValidVec_res_24 <= 1'h0;
      v0WriteValidVec_res_25 <= 1'h0;
      v0WriteValidVec_res_26 <= 1'h0;
      v0WriteValidVec_res_27 <= 1'h0;
      v0WriteValidVec_res_28 <= 1'h0;
      v0WriteValidVec_res_29 <= 1'h0;
      v0WriteValidVec_res_30 <= 1'h0;
      v0WriteValidVec_res_31 <= 1'h0;
      v0WriteValidVec_res_32 <= 1'h0;
      v0WriteValidVec_res_33 <= 1'h0;
      v0WriteValidVec_res_34 <= 1'h0;
      v0WriteValidVec_res_35 <= 1'h0;
      v0WriteValidVec_res_36 <= 1'h0;
      v0WriteValidVec_res_37 <= 1'h0;
      v0WriteValidVec_res_38 <= 1'h0;
      v0WriteValidVec_res_39 <= 1'h0;
      v0WriteValidVec_res_40 <= 1'h0;
      v0WriteValidVec_res_41 <= 1'h0;
      v0WriteValidVec_res_42 <= 1'h0;
      v0WriteValidVec_res_43 <= 1'h0;
      v0WriteValidVec_res_44 <= 1'h0;
      v0WriteValidVec_res_45 <= 1'h0;
      v0WriteValidVec_res_46 <= 1'h0;
      v0WriteValidVec_res_47 <= 1'h0;
      v0WriteValidVec_res_48 <= 1'h0;
      v0WriteValidVec_res_49 <= 1'h0;
      v0WriteValidVec_res_50 <= 1'h0;
      v0WriteValidVec_res_51 <= 1'h0;
      v0WriteValidVec_res_52 <= 1'h0;
      v0WriteValidVec_res_53 <= 1'h0;
      v0WriteValidVec_res_54 <= 1'h0;
      v0WriteValidVec_res_55 <= 1'h0;
      v0WriteValidVec_res_56 <= 1'h0;
      v0WriteValidVec_res_57 <= 1'h0;
      v0WriteValidVec_res_58 <= 1'h0;
      v0WriteValidVec_res_59 <= 1'h0;
      v0WriteValidVec_res_60 <= 1'h0;
      v0WriteValidVec_res_61 <= 1'h0;
      v0WriteValidVec_res_62 <= 1'h0;
      v0WriteValidVec_res_63 <= 1'h0;
      v0WriteValidVec_res_64 <= 1'h0;
      v0WriteValidVec_res_65 <= 1'h0;
      v0WriteValidVec_res_66 <= 1'h0;
      v0WriteValidVec_res_67 <= 1'h0;
      v0WriteValidVec_res_68 <= 1'h0;
      v0WriteValidVec_res_69 <= 1'h0;
      v0WriteValidVec_res_70 <= 1'h0;
      v0WriteValidVec_res_71 <= 1'h0;
      v0WriteValidVec_res_72 <= 1'h0;
      v0WriteValidVec_res_73 <= 1'h0;
      v0WriteValidVec_res_74 <= 1'h0;
      v0WriteValidVec_res_75 <= 1'h0;
      v0WriteValidVec_res_76 <= 1'h0;
      v0WriteValidVec_res_77 <= 1'h0;
      v0WriteValidVec_res_78 <= 1'h0;
      v0WriteValidVec_res_79 <= 1'h0;
      v0WriteValidVec_res_80 <= 1'h0;
      v0WriteValidVec_res_81 <= 1'h0;
      v0WriteValidVec_res_82 <= 1'h0;
      v0WriteValidVec_res_83 <= 1'h0;
      v0WriteValidVec_res_84 <= 1'h0;
      v0WriteValidVec_res_85 <= 1'h0;
      v0WriteValidVec_res_86 <= 1'h0;
      v0WriteValidVec_res_87 <= 1'h0;
      v0WriteValidVec_res_88 <= 1'h0;
      v0WriteValidVec_res_89 <= 1'h0;
      v0WriteValidVec_res_90 <= 1'h0;
      v0WriteValidVec_res_91 <= 1'h0;
      v0WriteValidVec_res_92 <= 1'h0;
      v0WriteValidVec_res_93 <= 1'h0;
      v0WriteValidVec_res_94 <= 1'h0;
      v0WriteValidVec_res_95 <= 1'h0;
      v0WriteValidVec_res_96 <= 1'h0;
      v0WriteValidVec_res_97 <= 1'h0;
      v0WriteValidVec_res_98 <= 1'h0;
      v0WriteValidVec_res_99 <= 1'h0;
      v0WriteValidVec_res_100 <= 1'h0;
      v0WriteValidVec_res_101 <= 1'h0;
      v0WriteValidVec_res_102 <= 1'h0;
      v0WriteValidVec_res_103 <= 1'h0;
      v0WriteValidVec_res_104 <= 1'h0;
      v0WriteValidVec_res_105 <= 1'h0;
      v0WriteValidVec_res_106 <= 1'h0;
      v0WriteValidVec_res_107 <= 1'h0;
      v0WriteValidVec_res_108 <= 1'h0;
      v0WriteValidVec_res_109 <= 1'h0;
      v0WriteValidVec_res_110 <= 1'h0;
      v0WriteValidVec_res_111 <= 1'h0;
      v0WriteValidVec_res_112 <= 1'h0;
      v0WriteValidVec_res_113 <= 1'h0;
      v0WriteValidVec_res_114 <= 1'h0;
      v0WriteValidVec_res_115 <= 1'h0;
      v0WriteValidVec_res_116 <= 1'h0;
      v0WriteValidVec_res_117 <= 1'h0;
      v0WriteValidVec_res_118 <= 1'h0;
      v0WriteValidVec_res_119 <= 1'h0;
      v0WriteValidVec_res_120 <= 1'h0;
      v0WriteValidVec_res_121 <= 1'h0;
      v0WriteValidVec_res_122 <= 1'h0;
      v0WriteValidVec_res_123 <= 1'h0;
      v0WriteValidVec_res_124 <= 1'h0;
      v0WriteValidVec_res_125 <= 1'h0;
      v0WriteValidVec_res_126 <= 1'h0;
      v0WriteValidVec_res_127 <= 1'h0;
      useV0AsMaskToken_res <= 1'h0;
      useV0AsMaskToken_res_1 <= 1'h0;
      useV0AsMaskToken_res_2 <= 1'h0;
      useV0AsMaskToken_res_3 <= 1'h0;
      useV0AsMaskToken_res_4 <= 1'h0;
      useV0AsMaskToken_res_5 <= 1'h0;
      useV0AsMaskToken_res_6 <= 1'h0;
      useV0AsMaskToken_res_7 <= 1'h0;
      useV0AsMaskToken_res_8 <= 1'h0;
      useV0AsMaskToken_res_9 <= 1'h0;
      useV0AsMaskToken_res_10 <= 1'h0;
      useV0AsMaskToken_res_11 <= 1'h0;
      useV0AsMaskToken_res_12 <= 1'h0;
      useV0AsMaskToken_res_13 <= 1'h0;
      useV0AsMaskToken_res_14 <= 1'h0;
      useV0AsMaskToken_res_15 <= 1'h0;
      useV0AsMaskToken_res_16 <= 1'h0;
      useV0AsMaskToken_res_17 <= 1'h0;
      useV0AsMaskToken_res_18 <= 1'h0;
      useV0AsMaskToken_res_19 <= 1'h0;
      useV0AsMaskToken_res_20 <= 1'h0;
      useV0AsMaskToken_res_21 <= 1'h0;
      useV0AsMaskToken_res_22 <= 1'h0;
      useV0AsMaskToken_res_23 <= 1'h0;
      useV0AsMaskToken_res_24 <= 1'h0;
      useV0AsMaskToken_res_25 <= 1'h0;
      useV0AsMaskToken_res_26 <= 1'h0;
      useV0AsMaskToken_res_27 <= 1'h0;
      useV0AsMaskToken_res_28 <= 1'h0;
      useV0AsMaskToken_res_29 <= 1'h0;
      useV0AsMaskToken_res_30 <= 1'h0;
      useV0AsMaskToken_res_31 <= 1'h0;
      useV0AsMaskToken_res_32 <= 1'h0;
      useV0AsMaskToken_res_33 <= 1'h0;
      useV0AsMaskToken_res_34 <= 1'h0;
      useV0AsMaskToken_res_35 <= 1'h0;
      useV0AsMaskToken_res_36 <= 1'h0;
      useV0AsMaskToken_res_37 <= 1'h0;
      useV0AsMaskToken_res_38 <= 1'h0;
      useV0AsMaskToken_res_39 <= 1'h0;
      useV0AsMaskToken_res_40 <= 1'h0;
      useV0AsMaskToken_res_41 <= 1'h0;
      useV0AsMaskToken_res_42 <= 1'h0;
      useV0AsMaskToken_res_43 <= 1'h0;
      useV0AsMaskToken_res_44 <= 1'h0;
      useV0AsMaskToken_res_45 <= 1'h0;
      useV0AsMaskToken_res_46 <= 1'h0;
      useV0AsMaskToken_res_47 <= 1'h0;
      useV0AsMaskToken_res_48 <= 1'h0;
      useV0AsMaskToken_res_49 <= 1'h0;
      useV0AsMaskToken_res_50 <= 1'h0;
      useV0AsMaskToken_res_51 <= 1'h0;
      useV0AsMaskToken_res_52 <= 1'h0;
      useV0AsMaskToken_res_53 <= 1'h0;
      useV0AsMaskToken_res_54 <= 1'h0;
      useV0AsMaskToken_res_55 <= 1'h0;
      useV0AsMaskToken_res_56 <= 1'h0;
      useV0AsMaskToken_res_57 <= 1'h0;
      useV0AsMaskToken_res_58 <= 1'h0;
      useV0AsMaskToken_res_59 <= 1'h0;
      useV0AsMaskToken_res_60 <= 1'h0;
      useV0AsMaskToken_res_61 <= 1'h0;
      useV0AsMaskToken_res_62 <= 1'h0;
      useV0AsMaskToken_res_63 <= 1'h0;
      useV0AsMaskToken_res_64 <= 1'h0;
      useV0AsMaskToken_res_65 <= 1'h0;
      useV0AsMaskToken_res_66 <= 1'h0;
      useV0AsMaskToken_res_67 <= 1'h0;
      useV0AsMaskToken_res_68 <= 1'h0;
      useV0AsMaskToken_res_69 <= 1'h0;
      useV0AsMaskToken_res_70 <= 1'h0;
      useV0AsMaskToken_res_71 <= 1'h0;
      useV0AsMaskToken_res_72 <= 1'h0;
      useV0AsMaskToken_res_73 <= 1'h0;
      useV0AsMaskToken_res_74 <= 1'h0;
      useV0AsMaskToken_res_75 <= 1'h0;
      useV0AsMaskToken_res_76 <= 1'h0;
      useV0AsMaskToken_res_77 <= 1'h0;
      useV0AsMaskToken_res_78 <= 1'h0;
      useV0AsMaskToken_res_79 <= 1'h0;
      useV0AsMaskToken_res_80 <= 1'h0;
      useV0AsMaskToken_res_81 <= 1'h0;
      useV0AsMaskToken_res_82 <= 1'h0;
      useV0AsMaskToken_res_83 <= 1'h0;
      useV0AsMaskToken_res_84 <= 1'h0;
      useV0AsMaskToken_res_85 <= 1'h0;
      useV0AsMaskToken_res_86 <= 1'h0;
      useV0AsMaskToken_res_87 <= 1'h0;
      useV0AsMaskToken_res_88 <= 1'h0;
      useV0AsMaskToken_res_89 <= 1'h0;
      useV0AsMaskToken_res_90 <= 1'h0;
      useV0AsMaskToken_res_91 <= 1'h0;
      useV0AsMaskToken_res_92 <= 1'h0;
      useV0AsMaskToken_res_93 <= 1'h0;
      useV0AsMaskToken_res_94 <= 1'h0;
      useV0AsMaskToken_res_95 <= 1'h0;
      useV0AsMaskToken_res_96 <= 1'h0;
      useV0AsMaskToken_res_97 <= 1'h0;
      useV0AsMaskToken_res_98 <= 1'h0;
      useV0AsMaskToken_res_99 <= 1'h0;
      useV0AsMaskToken_res_100 <= 1'h0;
      useV0AsMaskToken_res_101 <= 1'h0;
      useV0AsMaskToken_res_102 <= 1'h0;
      useV0AsMaskToken_res_103 <= 1'h0;
      useV0AsMaskToken_res_104 <= 1'h0;
      useV0AsMaskToken_res_105 <= 1'h0;
      useV0AsMaskToken_res_106 <= 1'h0;
      useV0AsMaskToken_res_107 <= 1'h0;
      useV0AsMaskToken_res_108 <= 1'h0;
      useV0AsMaskToken_res_109 <= 1'h0;
      useV0AsMaskToken_res_110 <= 1'h0;
      useV0AsMaskToken_res_111 <= 1'h0;
      useV0AsMaskToken_res_112 <= 1'h0;
      useV0AsMaskToken_res_113 <= 1'h0;
      useV0AsMaskToken_res_114 <= 1'h0;
      useV0AsMaskToken_res_115 <= 1'h0;
      useV0AsMaskToken_res_116 <= 1'h0;
      useV0AsMaskToken_res_117 <= 1'h0;
      useV0AsMaskToken_res_118 <= 1'h0;
      useV0AsMaskToken_res_119 <= 1'h0;
      useV0AsMaskToken_res_120 <= 1'h0;
      useV0AsMaskToken_res_121 <= 1'h0;
      useV0AsMaskToken_res_122 <= 1'h0;
      useV0AsMaskToken_res_123 <= 1'h0;
      useV0AsMaskToken_res_124 <= 1'h0;
      useV0AsMaskToken_res_125 <= 1'h0;
      useV0AsMaskToken_res_126 <= 1'h0;
      useV0AsMaskToken_res_127 <= 1'h0;
      maskUnitWriteV0 <= 1'h0;
    end
    else begin
      automatic logic [7:0] _v0WriteValidVec_T = v0WriteValidVec_updateOH | v0WriteValidVec_lsuWriteSet;
      automatic logic [7:0] _v0WriteValidVec_T_25 = v0WriteValidVec_updateOH_1 | v0WriteValidVec_lsuWriteSet_1;
      automatic logic [7:0] _v0WriteValidVec_T_50 = v0WriteValidVec_updateOH_2 | v0WriteValidVec_lsuWriteSet_2;
      automatic logic [7:0] _v0WriteValidVec_T_75 = v0WriteValidVec_updateOH_3 | v0WriteValidVec_lsuWriteSet_3;
      automatic logic [7:0] _v0WriteValidVec_T_100 = v0WriteValidVec_updateOH_4 | v0WriteValidVec_lsuWriteSet_4;
      automatic logic [7:0] _v0WriteValidVec_T_125 = v0WriteValidVec_updateOH_5 | v0WriteValidVec_lsuWriteSet_5;
      automatic logic [7:0] _v0WriteValidVec_T_150 = v0WriteValidVec_updateOH_6 | v0WriteValidVec_lsuWriteSet_6;
      automatic logic [7:0] _v0WriteValidVec_T_175 = v0WriteValidVec_updateOH_7 | v0WriteValidVec_lsuWriteSet_7;
      automatic logic [7:0] _v0WriteValidVec_T_200 = v0WriteValidVec_updateOH_8 | v0WriteValidVec_lsuWriteSet_8;
      automatic logic [7:0] _v0WriteValidVec_T_225 = v0WriteValidVec_updateOH_9 | v0WriteValidVec_lsuWriteSet_9;
      automatic logic [7:0] _v0WriteValidVec_T_250 = v0WriteValidVec_updateOH_10 | v0WriteValidVec_lsuWriteSet_10;
      automatic logic [7:0] _v0WriteValidVec_T_275 = v0WriteValidVec_updateOH_11 | v0WriteValidVec_lsuWriteSet_11;
      automatic logic [7:0] _v0WriteValidVec_T_300 = v0WriteValidVec_updateOH_12 | v0WriteValidVec_lsuWriteSet_12;
      automatic logic [7:0] _v0WriteValidVec_T_325 = v0WriteValidVec_updateOH_13 | v0WriteValidVec_lsuWriteSet_13;
      automatic logic [7:0] _v0WriteValidVec_T_350 = v0WriteValidVec_updateOH_14 | v0WriteValidVec_lsuWriteSet_14;
      automatic logic [7:0] _v0WriteValidVec_T_375 = v0WriteValidVec_updateOH_15 | v0WriteValidVec_lsuWriteSet_15;
      if (_v0WriteValidVec_T[0] | instructionFinish_0[0])
        v0WriteValidVec_res <= _v0WriteValidVec_T[0];
      if (_v0WriteValidVec_T[1] | instructionFinish_0[1])
        v0WriteValidVec_res_1 <= _v0WriteValidVec_T[1];
      if (_v0WriteValidVec_T[2] | instructionFinish_0[2])
        v0WriteValidVec_res_2 <= _v0WriteValidVec_T[2];
      if (_v0WriteValidVec_T[3] | instructionFinish_0[3])
        v0WriteValidVec_res_3 <= _v0WriteValidVec_T[3];
      if (_v0WriteValidVec_T[4] | instructionFinish_0[4])
        v0WriteValidVec_res_4 <= _v0WriteValidVec_T[4];
      if (_v0WriteValidVec_T[5] | instructionFinish_0[5])
        v0WriteValidVec_res_5 <= _v0WriteValidVec_T[5];
      if (_v0WriteValidVec_T[6] | instructionFinish_0[6])
        v0WriteValidVec_res_6 <= _v0WriteValidVec_T[6];
      if (_v0WriteValidVec_T[7] | instructionFinish_0[7])
        v0WriteValidVec_res_7 <= _v0WriteValidVec_T[7];
      if (_v0WriteValidVec_T_25[0] | instructionFinish_1[0])
        v0WriteValidVec_res_8 <= _v0WriteValidVec_T_25[0];
      if (_v0WriteValidVec_T_25[1] | instructionFinish_1[1])
        v0WriteValidVec_res_9 <= _v0WriteValidVec_T_25[1];
      if (_v0WriteValidVec_T_25[2] | instructionFinish_1[2])
        v0WriteValidVec_res_10 <= _v0WriteValidVec_T_25[2];
      if (_v0WriteValidVec_T_25[3] | instructionFinish_1[3])
        v0WriteValidVec_res_11 <= _v0WriteValidVec_T_25[3];
      if (_v0WriteValidVec_T_25[4] | instructionFinish_1[4])
        v0WriteValidVec_res_12 <= _v0WriteValidVec_T_25[4];
      if (_v0WriteValidVec_T_25[5] | instructionFinish_1[5])
        v0WriteValidVec_res_13 <= _v0WriteValidVec_T_25[5];
      if (_v0WriteValidVec_T_25[6] | instructionFinish_1[6])
        v0WriteValidVec_res_14 <= _v0WriteValidVec_T_25[6];
      if (_v0WriteValidVec_T_25[7] | instructionFinish_1[7])
        v0WriteValidVec_res_15 <= _v0WriteValidVec_T_25[7];
      if (_v0WriteValidVec_T_50[0] | instructionFinish_2[0])
        v0WriteValidVec_res_16 <= _v0WriteValidVec_T_50[0];
      if (_v0WriteValidVec_T_50[1] | instructionFinish_2[1])
        v0WriteValidVec_res_17 <= _v0WriteValidVec_T_50[1];
      if (_v0WriteValidVec_T_50[2] | instructionFinish_2[2])
        v0WriteValidVec_res_18 <= _v0WriteValidVec_T_50[2];
      if (_v0WriteValidVec_T_50[3] | instructionFinish_2[3])
        v0WriteValidVec_res_19 <= _v0WriteValidVec_T_50[3];
      if (_v0WriteValidVec_T_50[4] | instructionFinish_2[4])
        v0WriteValidVec_res_20 <= _v0WriteValidVec_T_50[4];
      if (_v0WriteValidVec_T_50[5] | instructionFinish_2[5])
        v0WriteValidVec_res_21 <= _v0WriteValidVec_T_50[5];
      if (_v0WriteValidVec_T_50[6] | instructionFinish_2[6])
        v0WriteValidVec_res_22 <= _v0WriteValidVec_T_50[6];
      if (_v0WriteValidVec_T_50[7] | instructionFinish_2[7])
        v0WriteValidVec_res_23 <= _v0WriteValidVec_T_50[7];
      if (_v0WriteValidVec_T_75[0] | instructionFinish_3[0])
        v0WriteValidVec_res_24 <= _v0WriteValidVec_T_75[0];
      if (_v0WriteValidVec_T_75[1] | instructionFinish_3[1])
        v0WriteValidVec_res_25 <= _v0WriteValidVec_T_75[1];
      if (_v0WriteValidVec_T_75[2] | instructionFinish_3[2])
        v0WriteValidVec_res_26 <= _v0WriteValidVec_T_75[2];
      if (_v0WriteValidVec_T_75[3] | instructionFinish_3[3])
        v0WriteValidVec_res_27 <= _v0WriteValidVec_T_75[3];
      if (_v0WriteValidVec_T_75[4] | instructionFinish_3[4])
        v0WriteValidVec_res_28 <= _v0WriteValidVec_T_75[4];
      if (_v0WriteValidVec_T_75[5] | instructionFinish_3[5])
        v0WriteValidVec_res_29 <= _v0WriteValidVec_T_75[5];
      if (_v0WriteValidVec_T_75[6] | instructionFinish_3[6])
        v0WriteValidVec_res_30 <= _v0WriteValidVec_T_75[6];
      if (_v0WriteValidVec_T_75[7] | instructionFinish_3[7])
        v0WriteValidVec_res_31 <= _v0WriteValidVec_T_75[7];
      if (_v0WriteValidVec_T_100[0] | instructionFinish_4[0])
        v0WriteValidVec_res_32 <= _v0WriteValidVec_T_100[0];
      if (_v0WriteValidVec_T_100[1] | instructionFinish_4[1])
        v0WriteValidVec_res_33 <= _v0WriteValidVec_T_100[1];
      if (_v0WriteValidVec_T_100[2] | instructionFinish_4[2])
        v0WriteValidVec_res_34 <= _v0WriteValidVec_T_100[2];
      if (_v0WriteValidVec_T_100[3] | instructionFinish_4[3])
        v0WriteValidVec_res_35 <= _v0WriteValidVec_T_100[3];
      if (_v0WriteValidVec_T_100[4] | instructionFinish_4[4])
        v0WriteValidVec_res_36 <= _v0WriteValidVec_T_100[4];
      if (_v0WriteValidVec_T_100[5] | instructionFinish_4[5])
        v0WriteValidVec_res_37 <= _v0WriteValidVec_T_100[5];
      if (_v0WriteValidVec_T_100[6] | instructionFinish_4[6])
        v0WriteValidVec_res_38 <= _v0WriteValidVec_T_100[6];
      if (_v0WriteValidVec_T_100[7] | instructionFinish_4[7])
        v0WriteValidVec_res_39 <= _v0WriteValidVec_T_100[7];
      if (_v0WriteValidVec_T_125[0] | instructionFinish_5[0])
        v0WriteValidVec_res_40 <= _v0WriteValidVec_T_125[0];
      if (_v0WriteValidVec_T_125[1] | instructionFinish_5[1])
        v0WriteValidVec_res_41 <= _v0WriteValidVec_T_125[1];
      if (_v0WriteValidVec_T_125[2] | instructionFinish_5[2])
        v0WriteValidVec_res_42 <= _v0WriteValidVec_T_125[2];
      if (_v0WriteValidVec_T_125[3] | instructionFinish_5[3])
        v0WriteValidVec_res_43 <= _v0WriteValidVec_T_125[3];
      if (_v0WriteValidVec_T_125[4] | instructionFinish_5[4])
        v0WriteValidVec_res_44 <= _v0WriteValidVec_T_125[4];
      if (_v0WriteValidVec_T_125[5] | instructionFinish_5[5])
        v0WriteValidVec_res_45 <= _v0WriteValidVec_T_125[5];
      if (_v0WriteValidVec_T_125[6] | instructionFinish_5[6])
        v0WriteValidVec_res_46 <= _v0WriteValidVec_T_125[6];
      if (_v0WriteValidVec_T_125[7] | instructionFinish_5[7])
        v0WriteValidVec_res_47 <= _v0WriteValidVec_T_125[7];
      if (_v0WriteValidVec_T_150[0] | instructionFinish_6[0])
        v0WriteValidVec_res_48 <= _v0WriteValidVec_T_150[0];
      if (_v0WriteValidVec_T_150[1] | instructionFinish_6[1])
        v0WriteValidVec_res_49 <= _v0WriteValidVec_T_150[1];
      if (_v0WriteValidVec_T_150[2] | instructionFinish_6[2])
        v0WriteValidVec_res_50 <= _v0WriteValidVec_T_150[2];
      if (_v0WriteValidVec_T_150[3] | instructionFinish_6[3])
        v0WriteValidVec_res_51 <= _v0WriteValidVec_T_150[3];
      if (_v0WriteValidVec_T_150[4] | instructionFinish_6[4])
        v0WriteValidVec_res_52 <= _v0WriteValidVec_T_150[4];
      if (_v0WriteValidVec_T_150[5] | instructionFinish_6[5])
        v0WriteValidVec_res_53 <= _v0WriteValidVec_T_150[5];
      if (_v0WriteValidVec_T_150[6] | instructionFinish_6[6])
        v0WriteValidVec_res_54 <= _v0WriteValidVec_T_150[6];
      if (_v0WriteValidVec_T_150[7] | instructionFinish_6[7])
        v0WriteValidVec_res_55 <= _v0WriteValidVec_T_150[7];
      if (_v0WriteValidVec_T_175[0] | instructionFinish_7[0])
        v0WriteValidVec_res_56 <= _v0WriteValidVec_T_175[0];
      if (_v0WriteValidVec_T_175[1] | instructionFinish_7[1])
        v0WriteValidVec_res_57 <= _v0WriteValidVec_T_175[1];
      if (_v0WriteValidVec_T_175[2] | instructionFinish_7[2])
        v0WriteValidVec_res_58 <= _v0WriteValidVec_T_175[2];
      if (_v0WriteValidVec_T_175[3] | instructionFinish_7[3])
        v0WriteValidVec_res_59 <= _v0WriteValidVec_T_175[3];
      if (_v0WriteValidVec_T_175[4] | instructionFinish_7[4])
        v0WriteValidVec_res_60 <= _v0WriteValidVec_T_175[4];
      if (_v0WriteValidVec_T_175[5] | instructionFinish_7[5])
        v0WriteValidVec_res_61 <= _v0WriteValidVec_T_175[5];
      if (_v0WriteValidVec_T_175[6] | instructionFinish_7[6])
        v0WriteValidVec_res_62 <= _v0WriteValidVec_T_175[6];
      if (_v0WriteValidVec_T_175[7] | instructionFinish_7[7])
        v0WriteValidVec_res_63 <= _v0WriteValidVec_T_175[7];
      if (_v0WriteValidVec_T_200[0] | instructionFinish_8[0])
        v0WriteValidVec_res_64 <= _v0WriteValidVec_T_200[0];
      if (_v0WriteValidVec_T_200[1] | instructionFinish_8[1])
        v0WriteValidVec_res_65 <= _v0WriteValidVec_T_200[1];
      if (_v0WriteValidVec_T_200[2] | instructionFinish_8[2])
        v0WriteValidVec_res_66 <= _v0WriteValidVec_T_200[2];
      if (_v0WriteValidVec_T_200[3] | instructionFinish_8[3])
        v0WriteValidVec_res_67 <= _v0WriteValidVec_T_200[3];
      if (_v0WriteValidVec_T_200[4] | instructionFinish_8[4])
        v0WriteValidVec_res_68 <= _v0WriteValidVec_T_200[4];
      if (_v0WriteValidVec_T_200[5] | instructionFinish_8[5])
        v0WriteValidVec_res_69 <= _v0WriteValidVec_T_200[5];
      if (_v0WriteValidVec_T_200[6] | instructionFinish_8[6])
        v0WriteValidVec_res_70 <= _v0WriteValidVec_T_200[6];
      if (_v0WriteValidVec_T_200[7] | instructionFinish_8[7])
        v0WriteValidVec_res_71 <= _v0WriteValidVec_T_200[7];
      if (_v0WriteValidVec_T_225[0] | instructionFinish_9[0])
        v0WriteValidVec_res_72 <= _v0WriteValidVec_T_225[0];
      if (_v0WriteValidVec_T_225[1] | instructionFinish_9[1])
        v0WriteValidVec_res_73 <= _v0WriteValidVec_T_225[1];
      if (_v0WriteValidVec_T_225[2] | instructionFinish_9[2])
        v0WriteValidVec_res_74 <= _v0WriteValidVec_T_225[2];
      if (_v0WriteValidVec_T_225[3] | instructionFinish_9[3])
        v0WriteValidVec_res_75 <= _v0WriteValidVec_T_225[3];
      if (_v0WriteValidVec_T_225[4] | instructionFinish_9[4])
        v0WriteValidVec_res_76 <= _v0WriteValidVec_T_225[4];
      if (_v0WriteValidVec_T_225[5] | instructionFinish_9[5])
        v0WriteValidVec_res_77 <= _v0WriteValidVec_T_225[5];
      if (_v0WriteValidVec_T_225[6] | instructionFinish_9[6])
        v0WriteValidVec_res_78 <= _v0WriteValidVec_T_225[6];
      if (_v0WriteValidVec_T_225[7] | instructionFinish_9[7])
        v0WriteValidVec_res_79 <= _v0WriteValidVec_T_225[7];
      if (_v0WriteValidVec_T_250[0] | instructionFinish_10[0])
        v0WriteValidVec_res_80 <= _v0WriteValidVec_T_250[0];
      if (_v0WriteValidVec_T_250[1] | instructionFinish_10[1])
        v0WriteValidVec_res_81 <= _v0WriteValidVec_T_250[1];
      if (_v0WriteValidVec_T_250[2] | instructionFinish_10[2])
        v0WriteValidVec_res_82 <= _v0WriteValidVec_T_250[2];
      if (_v0WriteValidVec_T_250[3] | instructionFinish_10[3])
        v0WriteValidVec_res_83 <= _v0WriteValidVec_T_250[3];
      if (_v0WriteValidVec_T_250[4] | instructionFinish_10[4])
        v0WriteValidVec_res_84 <= _v0WriteValidVec_T_250[4];
      if (_v0WriteValidVec_T_250[5] | instructionFinish_10[5])
        v0WriteValidVec_res_85 <= _v0WriteValidVec_T_250[5];
      if (_v0WriteValidVec_T_250[6] | instructionFinish_10[6])
        v0WriteValidVec_res_86 <= _v0WriteValidVec_T_250[6];
      if (_v0WriteValidVec_T_250[7] | instructionFinish_10[7])
        v0WriteValidVec_res_87 <= _v0WriteValidVec_T_250[7];
      if (_v0WriteValidVec_T_275[0] | instructionFinish_11[0])
        v0WriteValidVec_res_88 <= _v0WriteValidVec_T_275[0];
      if (_v0WriteValidVec_T_275[1] | instructionFinish_11[1])
        v0WriteValidVec_res_89 <= _v0WriteValidVec_T_275[1];
      if (_v0WriteValidVec_T_275[2] | instructionFinish_11[2])
        v0WriteValidVec_res_90 <= _v0WriteValidVec_T_275[2];
      if (_v0WriteValidVec_T_275[3] | instructionFinish_11[3])
        v0WriteValidVec_res_91 <= _v0WriteValidVec_T_275[3];
      if (_v0WriteValidVec_T_275[4] | instructionFinish_11[4])
        v0WriteValidVec_res_92 <= _v0WriteValidVec_T_275[4];
      if (_v0WriteValidVec_T_275[5] | instructionFinish_11[5])
        v0WriteValidVec_res_93 <= _v0WriteValidVec_T_275[5];
      if (_v0WriteValidVec_T_275[6] | instructionFinish_11[6])
        v0WriteValidVec_res_94 <= _v0WriteValidVec_T_275[6];
      if (_v0WriteValidVec_T_275[7] | instructionFinish_11[7])
        v0WriteValidVec_res_95 <= _v0WriteValidVec_T_275[7];
      if (_v0WriteValidVec_T_300[0] | instructionFinish_12[0])
        v0WriteValidVec_res_96 <= _v0WriteValidVec_T_300[0];
      if (_v0WriteValidVec_T_300[1] | instructionFinish_12[1])
        v0WriteValidVec_res_97 <= _v0WriteValidVec_T_300[1];
      if (_v0WriteValidVec_T_300[2] | instructionFinish_12[2])
        v0WriteValidVec_res_98 <= _v0WriteValidVec_T_300[2];
      if (_v0WriteValidVec_T_300[3] | instructionFinish_12[3])
        v0WriteValidVec_res_99 <= _v0WriteValidVec_T_300[3];
      if (_v0WriteValidVec_T_300[4] | instructionFinish_12[4])
        v0WriteValidVec_res_100 <= _v0WriteValidVec_T_300[4];
      if (_v0WriteValidVec_T_300[5] | instructionFinish_12[5])
        v0WriteValidVec_res_101 <= _v0WriteValidVec_T_300[5];
      if (_v0WriteValidVec_T_300[6] | instructionFinish_12[6])
        v0WriteValidVec_res_102 <= _v0WriteValidVec_T_300[6];
      if (_v0WriteValidVec_T_300[7] | instructionFinish_12[7])
        v0WriteValidVec_res_103 <= _v0WriteValidVec_T_300[7];
      if (_v0WriteValidVec_T_325[0] | instructionFinish_13[0])
        v0WriteValidVec_res_104 <= _v0WriteValidVec_T_325[0];
      if (_v0WriteValidVec_T_325[1] | instructionFinish_13[1])
        v0WriteValidVec_res_105 <= _v0WriteValidVec_T_325[1];
      if (_v0WriteValidVec_T_325[2] | instructionFinish_13[2])
        v0WriteValidVec_res_106 <= _v0WriteValidVec_T_325[2];
      if (_v0WriteValidVec_T_325[3] | instructionFinish_13[3])
        v0WriteValidVec_res_107 <= _v0WriteValidVec_T_325[3];
      if (_v0WriteValidVec_T_325[4] | instructionFinish_13[4])
        v0WriteValidVec_res_108 <= _v0WriteValidVec_T_325[4];
      if (_v0WriteValidVec_T_325[5] | instructionFinish_13[5])
        v0WriteValidVec_res_109 <= _v0WriteValidVec_T_325[5];
      if (_v0WriteValidVec_T_325[6] | instructionFinish_13[6])
        v0WriteValidVec_res_110 <= _v0WriteValidVec_T_325[6];
      if (_v0WriteValidVec_T_325[7] | instructionFinish_13[7])
        v0WriteValidVec_res_111 <= _v0WriteValidVec_T_325[7];
      if (_v0WriteValidVec_T_350[0] | instructionFinish_14[0])
        v0WriteValidVec_res_112 <= _v0WriteValidVec_T_350[0];
      if (_v0WriteValidVec_T_350[1] | instructionFinish_14[1])
        v0WriteValidVec_res_113 <= _v0WriteValidVec_T_350[1];
      if (_v0WriteValidVec_T_350[2] | instructionFinish_14[2])
        v0WriteValidVec_res_114 <= _v0WriteValidVec_T_350[2];
      if (_v0WriteValidVec_T_350[3] | instructionFinish_14[3])
        v0WriteValidVec_res_115 <= _v0WriteValidVec_T_350[3];
      if (_v0WriteValidVec_T_350[4] | instructionFinish_14[4])
        v0WriteValidVec_res_116 <= _v0WriteValidVec_T_350[4];
      if (_v0WriteValidVec_T_350[5] | instructionFinish_14[5])
        v0WriteValidVec_res_117 <= _v0WriteValidVec_T_350[5];
      if (_v0WriteValidVec_T_350[6] | instructionFinish_14[6])
        v0WriteValidVec_res_118 <= _v0WriteValidVec_T_350[6];
      if (_v0WriteValidVec_T_350[7] | instructionFinish_14[7])
        v0WriteValidVec_res_119 <= _v0WriteValidVec_T_350[7];
      if (_v0WriteValidVec_T_375[0] | instructionFinish_15[0])
        v0WriteValidVec_res_120 <= _v0WriteValidVec_T_375[0];
      if (_v0WriteValidVec_T_375[1] | instructionFinish_15[1])
        v0WriteValidVec_res_121 <= _v0WriteValidVec_T_375[1];
      if (_v0WriteValidVec_T_375[2] | instructionFinish_15[2])
        v0WriteValidVec_res_122 <= _v0WriteValidVec_T_375[2];
      if (_v0WriteValidVec_T_375[3] | instructionFinish_15[3])
        v0WriteValidVec_res_123 <= _v0WriteValidVec_T_375[3];
      if (_v0WriteValidVec_T_375[4] | instructionFinish_15[4])
        v0WriteValidVec_res_124 <= _v0WriteValidVec_T_375[4];
      if (_v0WriteValidVec_T_375[5] | instructionFinish_15[5])
        v0WriteValidVec_res_125 <= _v0WriteValidVec_T_375[5];
      if (_v0WriteValidVec_T_375[6] | instructionFinish_15[6])
        v0WriteValidVec_res_126 <= _v0WriteValidVec_T_375[6];
      if (_v0WriteValidVec_T_375[7] | instructionFinish_15[7])
        v0WriteValidVec_res_127 <= _v0WriteValidVec_T_375[7];
      if (useV0AsMaskToken_updateOH[0] | instructionFinish_0[0])
        useV0AsMaskToken_res <= useV0AsMaskToken_updateOH[0];
      if (useV0AsMaskToken_updateOH[1] | instructionFinish_0[1])
        useV0AsMaskToken_res_1 <= useV0AsMaskToken_updateOH[1];
      if (useV0AsMaskToken_updateOH[2] | instructionFinish_0[2])
        useV0AsMaskToken_res_2 <= useV0AsMaskToken_updateOH[2];
      if (useV0AsMaskToken_updateOH[3] | instructionFinish_0[3])
        useV0AsMaskToken_res_3 <= useV0AsMaskToken_updateOH[3];
      if (useV0AsMaskToken_updateOH[4] | instructionFinish_0[4])
        useV0AsMaskToken_res_4 <= useV0AsMaskToken_updateOH[4];
      if (useV0AsMaskToken_updateOH[5] | instructionFinish_0[5])
        useV0AsMaskToken_res_5 <= useV0AsMaskToken_updateOH[5];
      if (useV0AsMaskToken_updateOH[6] | instructionFinish_0[6])
        useV0AsMaskToken_res_6 <= useV0AsMaskToken_updateOH[6];
      if (useV0AsMaskToken_updateOH[7] | instructionFinish_0[7])
        useV0AsMaskToken_res_7 <= useV0AsMaskToken_updateOH[7];
      if (useV0AsMaskToken_updateOH_1[0] | instructionFinish_1[0])
        useV0AsMaskToken_res_8 <= useV0AsMaskToken_updateOH_1[0];
      if (useV0AsMaskToken_updateOH_1[1] | instructionFinish_1[1])
        useV0AsMaskToken_res_9 <= useV0AsMaskToken_updateOH_1[1];
      if (useV0AsMaskToken_updateOH_1[2] | instructionFinish_1[2])
        useV0AsMaskToken_res_10 <= useV0AsMaskToken_updateOH_1[2];
      if (useV0AsMaskToken_updateOH_1[3] | instructionFinish_1[3])
        useV0AsMaskToken_res_11 <= useV0AsMaskToken_updateOH_1[3];
      if (useV0AsMaskToken_updateOH_1[4] | instructionFinish_1[4])
        useV0AsMaskToken_res_12 <= useV0AsMaskToken_updateOH_1[4];
      if (useV0AsMaskToken_updateOH_1[5] | instructionFinish_1[5])
        useV0AsMaskToken_res_13 <= useV0AsMaskToken_updateOH_1[5];
      if (useV0AsMaskToken_updateOH_1[6] | instructionFinish_1[6])
        useV0AsMaskToken_res_14 <= useV0AsMaskToken_updateOH_1[6];
      if (useV0AsMaskToken_updateOH_1[7] | instructionFinish_1[7])
        useV0AsMaskToken_res_15 <= useV0AsMaskToken_updateOH_1[7];
      if (useV0AsMaskToken_updateOH_2[0] | instructionFinish_2[0])
        useV0AsMaskToken_res_16 <= useV0AsMaskToken_updateOH_2[0];
      if (useV0AsMaskToken_updateOH_2[1] | instructionFinish_2[1])
        useV0AsMaskToken_res_17 <= useV0AsMaskToken_updateOH_2[1];
      if (useV0AsMaskToken_updateOH_2[2] | instructionFinish_2[2])
        useV0AsMaskToken_res_18 <= useV0AsMaskToken_updateOH_2[2];
      if (useV0AsMaskToken_updateOH_2[3] | instructionFinish_2[3])
        useV0AsMaskToken_res_19 <= useV0AsMaskToken_updateOH_2[3];
      if (useV0AsMaskToken_updateOH_2[4] | instructionFinish_2[4])
        useV0AsMaskToken_res_20 <= useV0AsMaskToken_updateOH_2[4];
      if (useV0AsMaskToken_updateOH_2[5] | instructionFinish_2[5])
        useV0AsMaskToken_res_21 <= useV0AsMaskToken_updateOH_2[5];
      if (useV0AsMaskToken_updateOH_2[6] | instructionFinish_2[6])
        useV0AsMaskToken_res_22 <= useV0AsMaskToken_updateOH_2[6];
      if (useV0AsMaskToken_updateOH_2[7] | instructionFinish_2[7])
        useV0AsMaskToken_res_23 <= useV0AsMaskToken_updateOH_2[7];
      if (useV0AsMaskToken_updateOH_3[0] | instructionFinish_3[0])
        useV0AsMaskToken_res_24 <= useV0AsMaskToken_updateOH_3[0];
      if (useV0AsMaskToken_updateOH_3[1] | instructionFinish_3[1])
        useV0AsMaskToken_res_25 <= useV0AsMaskToken_updateOH_3[1];
      if (useV0AsMaskToken_updateOH_3[2] | instructionFinish_3[2])
        useV0AsMaskToken_res_26 <= useV0AsMaskToken_updateOH_3[2];
      if (useV0AsMaskToken_updateOH_3[3] | instructionFinish_3[3])
        useV0AsMaskToken_res_27 <= useV0AsMaskToken_updateOH_3[3];
      if (useV0AsMaskToken_updateOH_3[4] | instructionFinish_3[4])
        useV0AsMaskToken_res_28 <= useV0AsMaskToken_updateOH_3[4];
      if (useV0AsMaskToken_updateOH_3[5] | instructionFinish_3[5])
        useV0AsMaskToken_res_29 <= useV0AsMaskToken_updateOH_3[5];
      if (useV0AsMaskToken_updateOH_3[6] | instructionFinish_3[6])
        useV0AsMaskToken_res_30 <= useV0AsMaskToken_updateOH_3[6];
      if (useV0AsMaskToken_updateOH_3[7] | instructionFinish_3[7])
        useV0AsMaskToken_res_31 <= useV0AsMaskToken_updateOH_3[7];
      if (useV0AsMaskToken_updateOH_4[0] | instructionFinish_4[0])
        useV0AsMaskToken_res_32 <= useV0AsMaskToken_updateOH_4[0];
      if (useV0AsMaskToken_updateOH_4[1] | instructionFinish_4[1])
        useV0AsMaskToken_res_33 <= useV0AsMaskToken_updateOH_4[1];
      if (useV0AsMaskToken_updateOH_4[2] | instructionFinish_4[2])
        useV0AsMaskToken_res_34 <= useV0AsMaskToken_updateOH_4[2];
      if (useV0AsMaskToken_updateOH_4[3] | instructionFinish_4[3])
        useV0AsMaskToken_res_35 <= useV0AsMaskToken_updateOH_4[3];
      if (useV0AsMaskToken_updateOH_4[4] | instructionFinish_4[4])
        useV0AsMaskToken_res_36 <= useV0AsMaskToken_updateOH_4[4];
      if (useV0AsMaskToken_updateOH_4[5] | instructionFinish_4[5])
        useV0AsMaskToken_res_37 <= useV0AsMaskToken_updateOH_4[5];
      if (useV0AsMaskToken_updateOH_4[6] | instructionFinish_4[6])
        useV0AsMaskToken_res_38 <= useV0AsMaskToken_updateOH_4[6];
      if (useV0AsMaskToken_updateOH_4[7] | instructionFinish_4[7])
        useV0AsMaskToken_res_39 <= useV0AsMaskToken_updateOH_4[7];
      if (useV0AsMaskToken_updateOH_5[0] | instructionFinish_5[0])
        useV0AsMaskToken_res_40 <= useV0AsMaskToken_updateOH_5[0];
      if (useV0AsMaskToken_updateOH_5[1] | instructionFinish_5[1])
        useV0AsMaskToken_res_41 <= useV0AsMaskToken_updateOH_5[1];
      if (useV0AsMaskToken_updateOH_5[2] | instructionFinish_5[2])
        useV0AsMaskToken_res_42 <= useV0AsMaskToken_updateOH_5[2];
      if (useV0AsMaskToken_updateOH_5[3] | instructionFinish_5[3])
        useV0AsMaskToken_res_43 <= useV0AsMaskToken_updateOH_5[3];
      if (useV0AsMaskToken_updateOH_5[4] | instructionFinish_5[4])
        useV0AsMaskToken_res_44 <= useV0AsMaskToken_updateOH_5[4];
      if (useV0AsMaskToken_updateOH_5[5] | instructionFinish_5[5])
        useV0AsMaskToken_res_45 <= useV0AsMaskToken_updateOH_5[5];
      if (useV0AsMaskToken_updateOH_5[6] | instructionFinish_5[6])
        useV0AsMaskToken_res_46 <= useV0AsMaskToken_updateOH_5[6];
      if (useV0AsMaskToken_updateOH_5[7] | instructionFinish_5[7])
        useV0AsMaskToken_res_47 <= useV0AsMaskToken_updateOH_5[7];
      if (useV0AsMaskToken_updateOH_6[0] | instructionFinish_6[0])
        useV0AsMaskToken_res_48 <= useV0AsMaskToken_updateOH_6[0];
      if (useV0AsMaskToken_updateOH_6[1] | instructionFinish_6[1])
        useV0AsMaskToken_res_49 <= useV0AsMaskToken_updateOH_6[1];
      if (useV0AsMaskToken_updateOH_6[2] | instructionFinish_6[2])
        useV0AsMaskToken_res_50 <= useV0AsMaskToken_updateOH_6[2];
      if (useV0AsMaskToken_updateOH_6[3] | instructionFinish_6[3])
        useV0AsMaskToken_res_51 <= useV0AsMaskToken_updateOH_6[3];
      if (useV0AsMaskToken_updateOH_6[4] | instructionFinish_6[4])
        useV0AsMaskToken_res_52 <= useV0AsMaskToken_updateOH_6[4];
      if (useV0AsMaskToken_updateOH_6[5] | instructionFinish_6[5])
        useV0AsMaskToken_res_53 <= useV0AsMaskToken_updateOH_6[5];
      if (useV0AsMaskToken_updateOH_6[6] | instructionFinish_6[6])
        useV0AsMaskToken_res_54 <= useV0AsMaskToken_updateOH_6[6];
      if (useV0AsMaskToken_updateOH_6[7] | instructionFinish_6[7])
        useV0AsMaskToken_res_55 <= useV0AsMaskToken_updateOH_6[7];
      if (useV0AsMaskToken_updateOH_7[0] | instructionFinish_7[0])
        useV0AsMaskToken_res_56 <= useV0AsMaskToken_updateOH_7[0];
      if (useV0AsMaskToken_updateOH_7[1] | instructionFinish_7[1])
        useV0AsMaskToken_res_57 <= useV0AsMaskToken_updateOH_7[1];
      if (useV0AsMaskToken_updateOH_7[2] | instructionFinish_7[2])
        useV0AsMaskToken_res_58 <= useV0AsMaskToken_updateOH_7[2];
      if (useV0AsMaskToken_updateOH_7[3] | instructionFinish_7[3])
        useV0AsMaskToken_res_59 <= useV0AsMaskToken_updateOH_7[3];
      if (useV0AsMaskToken_updateOH_7[4] | instructionFinish_7[4])
        useV0AsMaskToken_res_60 <= useV0AsMaskToken_updateOH_7[4];
      if (useV0AsMaskToken_updateOH_7[5] | instructionFinish_7[5])
        useV0AsMaskToken_res_61 <= useV0AsMaskToken_updateOH_7[5];
      if (useV0AsMaskToken_updateOH_7[6] | instructionFinish_7[6])
        useV0AsMaskToken_res_62 <= useV0AsMaskToken_updateOH_7[6];
      if (useV0AsMaskToken_updateOH_7[7] | instructionFinish_7[7])
        useV0AsMaskToken_res_63 <= useV0AsMaskToken_updateOH_7[7];
      if (useV0AsMaskToken_updateOH_8[0] | instructionFinish_8[0])
        useV0AsMaskToken_res_64 <= useV0AsMaskToken_updateOH_8[0];
      if (useV0AsMaskToken_updateOH_8[1] | instructionFinish_8[1])
        useV0AsMaskToken_res_65 <= useV0AsMaskToken_updateOH_8[1];
      if (useV0AsMaskToken_updateOH_8[2] | instructionFinish_8[2])
        useV0AsMaskToken_res_66 <= useV0AsMaskToken_updateOH_8[2];
      if (useV0AsMaskToken_updateOH_8[3] | instructionFinish_8[3])
        useV0AsMaskToken_res_67 <= useV0AsMaskToken_updateOH_8[3];
      if (useV0AsMaskToken_updateOH_8[4] | instructionFinish_8[4])
        useV0AsMaskToken_res_68 <= useV0AsMaskToken_updateOH_8[4];
      if (useV0AsMaskToken_updateOH_8[5] | instructionFinish_8[5])
        useV0AsMaskToken_res_69 <= useV0AsMaskToken_updateOH_8[5];
      if (useV0AsMaskToken_updateOH_8[6] | instructionFinish_8[6])
        useV0AsMaskToken_res_70 <= useV0AsMaskToken_updateOH_8[6];
      if (useV0AsMaskToken_updateOH_8[7] | instructionFinish_8[7])
        useV0AsMaskToken_res_71 <= useV0AsMaskToken_updateOH_8[7];
      if (useV0AsMaskToken_updateOH_9[0] | instructionFinish_9[0])
        useV0AsMaskToken_res_72 <= useV0AsMaskToken_updateOH_9[0];
      if (useV0AsMaskToken_updateOH_9[1] | instructionFinish_9[1])
        useV0AsMaskToken_res_73 <= useV0AsMaskToken_updateOH_9[1];
      if (useV0AsMaskToken_updateOH_9[2] | instructionFinish_9[2])
        useV0AsMaskToken_res_74 <= useV0AsMaskToken_updateOH_9[2];
      if (useV0AsMaskToken_updateOH_9[3] | instructionFinish_9[3])
        useV0AsMaskToken_res_75 <= useV0AsMaskToken_updateOH_9[3];
      if (useV0AsMaskToken_updateOH_9[4] | instructionFinish_9[4])
        useV0AsMaskToken_res_76 <= useV0AsMaskToken_updateOH_9[4];
      if (useV0AsMaskToken_updateOH_9[5] | instructionFinish_9[5])
        useV0AsMaskToken_res_77 <= useV0AsMaskToken_updateOH_9[5];
      if (useV0AsMaskToken_updateOH_9[6] | instructionFinish_9[6])
        useV0AsMaskToken_res_78 <= useV0AsMaskToken_updateOH_9[6];
      if (useV0AsMaskToken_updateOH_9[7] | instructionFinish_9[7])
        useV0AsMaskToken_res_79 <= useV0AsMaskToken_updateOH_9[7];
      if (useV0AsMaskToken_updateOH_10[0] | instructionFinish_10[0])
        useV0AsMaskToken_res_80 <= useV0AsMaskToken_updateOH_10[0];
      if (useV0AsMaskToken_updateOH_10[1] | instructionFinish_10[1])
        useV0AsMaskToken_res_81 <= useV0AsMaskToken_updateOH_10[1];
      if (useV0AsMaskToken_updateOH_10[2] | instructionFinish_10[2])
        useV0AsMaskToken_res_82 <= useV0AsMaskToken_updateOH_10[2];
      if (useV0AsMaskToken_updateOH_10[3] | instructionFinish_10[3])
        useV0AsMaskToken_res_83 <= useV0AsMaskToken_updateOH_10[3];
      if (useV0AsMaskToken_updateOH_10[4] | instructionFinish_10[4])
        useV0AsMaskToken_res_84 <= useV0AsMaskToken_updateOH_10[4];
      if (useV0AsMaskToken_updateOH_10[5] | instructionFinish_10[5])
        useV0AsMaskToken_res_85 <= useV0AsMaskToken_updateOH_10[5];
      if (useV0AsMaskToken_updateOH_10[6] | instructionFinish_10[6])
        useV0AsMaskToken_res_86 <= useV0AsMaskToken_updateOH_10[6];
      if (useV0AsMaskToken_updateOH_10[7] | instructionFinish_10[7])
        useV0AsMaskToken_res_87 <= useV0AsMaskToken_updateOH_10[7];
      if (useV0AsMaskToken_updateOH_11[0] | instructionFinish_11[0])
        useV0AsMaskToken_res_88 <= useV0AsMaskToken_updateOH_11[0];
      if (useV0AsMaskToken_updateOH_11[1] | instructionFinish_11[1])
        useV0AsMaskToken_res_89 <= useV0AsMaskToken_updateOH_11[1];
      if (useV0AsMaskToken_updateOH_11[2] | instructionFinish_11[2])
        useV0AsMaskToken_res_90 <= useV0AsMaskToken_updateOH_11[2];
      if (useV0AsMaskToken_updateOH_11[3] | instructionFinish_11[3])
        useV0AsMaskToken_res_91 <= useV0AsMaskToken_updateOH_11[3];
      if (useV0AsMaskToken_updateOH_11[4] | instructionFinish_11[4])
        useV0AsMaskToken_res_92 <= useV0AsMaskToken_updateOH_11[4];
      if (useV0AsMaskToken_updateOH_11[5] | instructionFinish_11[5])
        useV0AsMaskToken_res_93 <= useV0AsMaskToken_updateOH_11[5];
      if (useV0AsMaskToken_updateOH_11[6] | instructionFinish_11[6])
        useV0AsMaskToken_res_94 <= useV0AsMaskToken_updateOH_11[6];
      if (useV0AsMaskToken_updateOH_11[7] | instructionFinish_11[7])
        useV0AsMaskToken_res_95 <= useV0AsMaskToken_updateOH_11[7];
      if (useV0AsMaskToken_updateOH_12[0] | instructionFinish_12[0])
        useV0AsMaskToken_res_96 <= useV0AsMaskToken_updateOH_12[0];
      if (useV0AsMaskToken_updateOH_12[1] | instructionFinish_12[1])
        useV0AsMaskToken_res_97 <= useV0AsMaskToken_updateOH_12[1];
      if (useV0AsMaskToken_updateOH_12[2] | instructionFinish_12[2])
        useV0AsMaskToken_res_98 <= useV0AsMaskToken_updateOH_12[2];
      if (useV0AsMaskToken_updateOH_12[3] | instructionFinish_12[3])
        useV0AsMaskToken_res_99 <= useV0AsMaskToken_updateOH_12[3];
      if (useV0AsMaskToken_updateOH_12[4] | instructionFinish_12[4])
        useV0AsMaskToken_res_100 <= useV0AsMaskToken_updateOH_12[4];
      if (useV0AsMaskToken_updateOH_12[5] | instructionFinish_12[5])
        useV0AsMaskToken_res_101 <= useV0AsMaskToken_updateOH_12[5];
      if (useV0AsMaskToken_updateOH_12[6] | instructionFinish_12[6])
        useV0AsMaskToken_res_102 <= useV0AsMaskToken_updateOH_12[6];
      if (useV0AsMaskToken_updateOH_12[7] | instructionFinish_12[7])
        useV0AsMaskToken_res_103 <= useV0AsMaskToken_updateOH_12[7];
      if (useV0AsMaskToken_updateOH_13[0] | instructionFinish_13[0])
        useV0AsMaskToken_res_104 <= useV0AsMaskToken_updateOH_13[0];
      if (useV0AsMaskToken_updateOH_13[1] | instructionFinish_13[1])
        useV0AsMaskToken_res_105 <= useV0AsMaskToken_updateOH_13[1];
      if (useV0AsMaskToken_updateOH_13[2] | instructionFinish_13[2])
        useV0AsMaskToken_res_106 <= useV0AsMaskToken_updateOH_13[2];
      if (useV0AsMaskToken_updateOH_13[3] | instructionFinish_13[3])
        useV0AsMaskToken_res_107 <= useV0AsMaskToken_updateOH_13[3];
      if (useV0AsMaskToken_updateOH_13[4] | instructionFinish_13[4])
        useV0AsMaskToken_res_108 <= useV0AsMaskToken_updateOH_13[4];
      if (useV0AsMaskToken_updateOH_13[5] | instructionFinish_13[5])
        useV0AsMaskToken_res_109 <= useV0AsMaskToken_updateOH_13[5];
      if (useV0AsMaskToken_updateOH_13[6] | instructionFinish_13[6])
        useV0AsMaskToken_res_110 <= useV0AsMaskToken_updateOH_13[6];
      if (useV0AsMaskToken_updateOH_13[7] | instructionFinish_13[7])
        useV0AsMaskToken_res_111 <= useV0AsMaskToken_updateOH_13[7];
      if (useV0AsMaskToken_updateOH_14[0] | instructionFinish_14[0])
        useV0AsMaskToken_res_112 <= useV0AsMaskToken_updateOH_14[0];
      if (useV0AsMaskToken_updateOH_14[1] | instructionFinish_14[1])
        useV0AsMaskToken_res_113 <= useV0AsMaskToken_updateOH_14[1];
      if (useV0AsMaskToken_updateOH_14[2] | instructionFinish_14[2])
        useV0AsMaskToken_res_114 <= useV0AsMaskToken_updateOH_14[2];
      if (useV0AsMaskToken_updateOH_14[3] | instructionFinish_14[3])
        useV0AsMaskToken_res_115 <= useV0AsMaskToken_updateOH_14[3];
      if (useV0AsMaskToken_updateOH_14[4] | instructionFinish_14[4])
        useV0AsMaskToken_res_116 <= useV0AsMaskToken_updateOH_14[4];
      if (useV0AsMaskToken_updateOH_14[5] | instructionFinish_14[5])
        useV0AsMaskToken_res_117 <= useV0AsMaskToken_updateOH_14[5];
      if (useV0AsMaskToken_updateOH_14[6] | instructionFinish_14[6])
        useV0AsMaskToken_res_118 <= useV0AsMaskToken_updateOH_14[6];
      if (useV0AsMaskToken_updateOH_14[7] | instructionFinish_14[7])
        useV0AsMaskToken_res_119 <= useV0AsMaskToken_updateOH_14[7];
      if (useV0AsMaskToken_updateOH_15[0] | instructionFinish_15[0])
        useV0AsMaskToken_res_120 <= useV0AsMaskToken_updateOH_15[0];
      if (useV0AsMaskToken_updateOH_15[1] | instructionFinish_15[1])
        useV0AsMaskToken_res_121 <= useV0AsMaskToken_updateOH_15[1];
      if (useV0AsMaskToken_updateOH_15[2] | instructionFinish_15[2])
        useV0AsMaskToken_res_122 <= useV0AsMaskToken_updateOH_15[2];
      if (useV0AsMaskToken_updateOH_15[3] | instructionFinish_15[3])
        useV0AsMaskToken_res_123 <= useV0AsMaskToken_updateOH_15[3];
      if (useV0AsMaskToken_updateOH_15[4] | instructionFinish_15[4])
        useV0AsMaskToken_res_124 <= useV0AsMaskToken_updateOH_15[4];
      if (useV0AsMaskToken_updateOH_15[5] | instructionFinish_15[5])
        useV0AsMaskToken_res_125 <= useV0AsMaskToken_updateOH_15[5];
      if (useV0AsMaskToken_updateOH_15[6] | instructionFinish_15[6])
        useV0AsMaskToken_res_126 <= useV0AsMaskToken_updateOH_15[6];
      if (useV0AsMaskToken_updateOH_15[7] | instructionFinish_15[7])
        useV0AsMaskToken_res_127 <= useV0AsMaskToken_updateOH_15[7];
      if (maskUnitWriteV0_set | maskUnitFree)
        maskUnitWriteV0 <= maskUnitWriteV0_set;
    end
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:8];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [3:0] i = 4'h0; i < 4'h9; i += 4'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        v0WriteValidVec_res = _RANDOM[4'h0][0];
        v0WriteValidVec_res_1 = _RANDOM[4'h0][1];
        v0WriteValidVec_res_2 = _RANDOM[4'h0][2];
        v0WriteValidVec_res_3 = _RANDOM[4'h0][3];
        v0WriteValidVec_res_4 = _RANDOM[4'h0][4];
        v0WriteValidVec_res_5 = _RANDOM[4'h0][5];
        v0WriteValidVec_res_6 = _RANDOM[4'h0][6];
        v0WriteValidVec_res_7 = _RANDOM[4'h0][7];
        v0WriteValidVec_res_8 = _RANDOM[4'h0][8];
        v0WriteValidVec_res_9 = _RANDOM[4'h0][9];
        v0WriteValidVec_res_10 = _RANDOM[4'h0][10];
        v0WriteValidVec_res_11 = _RANDOM[4'h0][11];
        v0WriteValidVec_res_12 = _RANDOM[4'h0][12];
        v0WriteValidVec_res_13 = _RANDOM[4'h0][13];
        v0WriteValidVec_res_14 = _RANDOM[4'h0][14];
        v0WriteValidVec_res_15 = _RANDOM[4'h0][15];
        v0WriteValidVec_res_16 = _RANDOM[4'h0][16];
        v0WriteValidVec_res_17 = _RANDOM[4'h0][17];
        v0WriteValidVec_res_18 = _RANDOM[4'h0][18];
        v0WriteValidVec_res_19 = _RANDOM[4'h0][19];
        v0WriteValidVec_res_20 = _RANDOM[4'h0][20];
        v0WriteValidVec_res_21 = _RANDOM[4'h0][21];
        v0WriteValidVec_res_22 = _RANDOM[4'h0][22];
        v0WriteValidVec_res_23 = _RANDOM[4'h0][23];
        v0WriteValidVec_res_24 = _RANDOM[4'h0][24];
        v0WriteValidVec_res_25 = _RANDOM[4'h0][25];
        v0WriteValidVec_res_26 = _RANDOM[4'h0][26];
        v0WriteValidVec_res_27 = _RANDOM[4'h0][27];
        v0WriteValidVec_res_28 = _RANDOM[4'h0][28];
        v0WriteValidVec_res_29 = _RANDOM[4'h0][29];
        v0WriteValidVec_res_30 = _RANDOM[4'h0][30];
        v0WriteValidVec_res_31 = _RANDOM[4'h0][31];
        v0WriteValidVec_res_32 = _RANDOM[4'h1][0];
        v0WriteValidVec_res_33 = _RANDOM[4'h1][1];
        v0WriteValidVec_res_34 = _RANDOM[4'h1][2];
        v0WriteValidVec_res_35 = _RANDOM[4'h1][3];
        v0WriteValidVec_res_36 = _RANDOM[4'h1][4];
        v0WriteValidVec_res_37 = _RANDOM[4'h1][5];
        v0WriteValidVec_res_38 = _RANDOM[4'h1][6];
        v0WriteValidVec_res_39 = _RANDOM[4'h1][7];
        v0WriteValidVec_res_40 = _RANDOM[4'h1][8];
        v0WriteValidVec_res_41 = _RANDOM[4'h1][9];
        v0WriteValidVec_res_42 = _RANDOM[4'h1][10];
        v0WriteValidVec_res_43 = _RANDOM[4'h1][11];
        v0WriteValidVec_res_44 = _RANDOM[4'h1][12];
        v0WriteValidVec_res_45 = _RANDOM[4'h1][13];
        v0WriteValidVec_res_46 = _RANDOM[4'h1][14];
        v0WriteValidVec_res_47 = _RANDOM[4'h1][15];
        v0WriteValidVec_res_48 = _RANDOM[4'h1][16];
        v0WriteValidVec_res_49 = _RANDOM[4'h1][17];
        v0WriteValidVec_res_50 = _RANDOM[4'h1][18];
        v0WriteValidVec_res_51 = _RANDOM[4'h1][19];
        v0WriteValidVec_res_52 = _RANDOM[4'h1][20];
        v0WriteValidVec_res_53 = _RANDOM[4'h1][21];
        v0WriteValidVec_res_54 = _RANDOM[4'h1][22];
        v0WriteValidVec_res_55 = _RANDOM[4'h1][23];
        v0WriteValidVec_res_56 = _RANDOM[4'h1][24];
        v0WriteValidVec_res_57 = _RANDOM[4'h1][25];
        v0WriteValidVec_res_58 = _RANDOM[4'h1][26];
        v0WriteValidVec_res_59 = _RANDOM[4'h1][27];
        v0WriteValidVec_res_60 = _RANDOM[4'h1][28];
        v0WriteValidVec_res_61 = _RANDOM[4'h1][29];
        v0WriteValidVec_res_62 = _RANDOM[4'h1][30];
        v0WriteValidVec_res_63 = _RANDOM[4'h1][31];
        v0WriteValidVec_res_64 = _RANDOM[4'h2][0];
        v0WriteValidVec_res_65 = _RANDOM[4'h2][1];
        v0WriteValidVec_res_66 = _RANDOM[4'h2][2];
        v0WriteValidVec_res_67 = _RANDOM[4'h2][3];
        v0WriteValidVec_res_68 = _RANDOM[4'h2][4];
        v0WriteValidVec_res_69 = _RANDOM[4'h2][5];
        v0WriteValidVec_res_70 = _RANDOM[4'h2][6];
        v0WriteValidVec_res_71 = _RANDOM[4'h2][7];
        v0WriteValidVec_res_72 = _RANDOM[4'h2][8];
        v0WriteValidVec_res_73 = _RANDOM[4'h2][9];
        v0WriteValidVec_res_74 = _RANDOM[4'h2][10];
        v0WriteValidVec_res_75 = _RANDOM[4'h2][11];
        v0WriteValidVec_res_76 = _RANDOM[4'h2][12];
        v0WriteValidVec_res_77 = _RANDOM[4'h2][13];
        v0WriteValidVec_res_78 = _RANDOM[4'h2][14];
        v0WriteValidVec_res_79 = _RANDOM[4'h2][15];
        v0WriteValidVec_res_80 = _RANDOM[4'h2][16];
        v0WriteValidVec_res_81 = _RANDOM[4'h2][17];
        v0WriteValidVec_res_82 = _RANDOM[4'h2][18];
        v0WriteValidVec_res_83 = _RANDOM[4'h2][19];
        v0WriteValidVec_res_84 = _RANDOM[4'h2][20];
        v0WriteValidVec_res_85 = _RANDOM[4'h2][21];
        v0WriteValidVec_res_86 = _RANDOM[4'h2][22];
        v0WriteValidVec_res_87 = _RANDOM[4'h2][23];
        v0WriteValidVec_res_88 = _RANDOM[4'h2][24];
        v0WriteValidVec_res_89 = _RANDOM[4'h2][25];
        v0WriteValidVec_res_90 = _RANDOM[4'h2][26];
        v0WriteValidVec_res_91 = _RANDOM[4'h2][27];
        v0WriteValidVec_res_92 = _RANDOM[4'h2][28];
        v0WriteValidVec_res_93 = _RANDOM[4'h2][29];
        v0WriteValidVec_res_94 = _RANDOM[4'h2][30];
        v0WriteValidVec_res_95 = _RANDOM[4'h2][31];
        v0WriteValidVec_res_96 = _RANDOM[4'h3][0];
        v0WriteValidVec_res_97 = _RANDOM[4'h3][1];
        v0WriteValidVec_res_98 = _RANDOM[4'h3][2];
        v0WriteValidVec_res_99 = _RANDOM[4'h3][3];
        v0WriteValidVec_res_100 = _RANDOM[4'h3][4];
        v0WriteValidVec_res_101 = _RANDOM[4'h3][5];
        v0WriteValidVec_res_102 = _RANDOM[4'h3][6];
        v0WriteValidVec_res_103 = _RANDOM[4'h3][7];
        v0WriteValidVec_res_104 = _RANDOM[4'h3][8];
        v0WriteValidVec_res_105 = _RANDOM[4'h3][9];
        v0WriteValidVec_res_106 = _RANDOM[4'h3][10];
        v0WriteValidVec_res_107 = _RANDOM[4'h3][11];
        v0WriteValidVec_res_108 = _RANDOM[4'h3][12];
        v0WriteValidVec_res_109 = _RANDOM[4'h3][13];
        v0WriteValidVec_res_110 = _RANDOM[4'h3][14];
        v0WriteValidVec_res_111 = _RANDOM[4'h3][15];
        v0WriteValidVec_res_112 = _RANDOM[4'h3][16];
        v0WriteValidVec_res_113 = _RANDOM[4'h3][17];
        v0WriteValidVec_res_114 = _RANDOM[4'h3][18];
        v0WriteValidVec_res_115 = _RANDOM[4'h3][19];
        v0WriteValidVec_res_116 = _RANDOM[4'h3][20];
        v0WriteValidVec_res_117 = _RANDOM[4'h3][21];
        v0WriteValidVec_res_118 = _RANDOM[4'h3][22];
        v0WriteValidVec_res_119 = _RANDOM[4'h3][23];
        v0WriteValidVec_res_120 = _RANDOM[4'h3][24];
        v0WriteValidVec_res_121 = _RANDOM[4'h3][25];
        v0WriteValidVec_res_122 = _RANDOM[4'h3][26];
        v0WriteValidVec_res_123 = _RANDOM[4'h3][27];
        v0WriteValidVec_res_124 = _RANDOM[4'h3][28];
        v0WriteValidVec_res_125 = _RANDOM[4'h3][29];
        v0WriteValidVec_res_126 = _RANDOM[4'h3][30];
        v0WriteValidVec_res_127 = _RANDOM[4'h3][31];
        useV0AsMaskToken_res = _RANDOM[4'h4][0];
        useV0AsMaskToken_res_1 = _RANDOM[4'h4][1];
        useV0AsMaskToken_res_2 = _RANDOM[4'h4][2];
        useV0AsMaskToken_res_3 = _RANDOM[4'h4][3];
        useV0AsMaskToken_res_4 = _RANDOM[4'h4][4];
        useV0AsMaskToken_res_5 = _RANDOM[4'h4][5];
        useV0AsMaskToken_res_6 = _RANDOM[4'h4][6];
        useV0AsMaskToken_res_7 = _RANDOM[4'h4][7];
        useV0AsMaskToken_res_8 = _RANDOM[4'h4][8];
        useV0AsMaskToken_res_9 = _RANDOM[4'h4][9];
        useV0AsMaskToken_res_10 = _RANDOM[4'h4][10];
        useV0AsMaskToken_res_11 = _RANDOM[4'h4][11];
        useV0AsMaskToken_res_12 = _RANDOM[4'h4][12];
        useV0AsMaskToken_res_13 = _RANDOM[4'h4][13];
        useV0AsMaskToken_res_14 = _RANDOM[4'h4][14];
        useV0AsMaskToken_res_15 = _RANDOM[4'h4][15];
        useV0AsMaskToken_res_16 = _RANDOM[4'h4][16];
        useV0AsMaskToken_res_17 = _RANDOM[4'h4][17];
        useV0AsMaskToken_res_18 = _RANDOM[4'h4][18];
        useV0AsMaskToken_res_19 = _RANDOM[4'h4][19];
        useV0AsMaskToken_res_20 = _RANDOM[4'h4][20];
        useV0AsMaskToken_res_21 = _RANDOM[4'h4][21];
        useV0AsMaskToken_res_22 = _RANDOM[4'h4][22];
        useV0AsMaskToken_res_23 = _RANDOM[4'h4][23];
        useV0AsMaskToken_res_24 = _RANDOM[4'h4][24];
        useV0AsMaskToken_res_25 = _RANDOM[4'h4][25];
        useV0AsMaskToken_res_26 = _RANDOM[4'h4][26];
        useV0AsMaskToken_res_27 = _RANDOM[4'h4][27];
        useV0AsMaskToken_res_28 = _RANDOM[4'h4][28];
        useV0AsMaskToken_res_29 = _RANDOM[4'h4][29];
        useV0AsMaskToken_res_30 = _RANDOM[4'h4][30];
        useV0AsMaskToken_res_31 = _RANDOM[4'h4][31];
        useV0AsMaskToken_res_32 = _RANDOM[4'h5][0];
        useV0AsMaskToken_res_33 = _RANDOM[4'h5][1];
        useV0AsMaskToken_res_34 = _RANDOM[4'h5][2];
        useV0AsMaskToken_res_35 = _RANDOM[4'h5][3];
        useV0AsMaskToken_res_36 = _RANDOM[4'h5][4];
        useV0AsMaskToken_res_37 = _RANDOM[4'h5][5];
        useV0AsMaskToken_res_38 = _RANDOM[4'h5][6];
        useV0AsMaskToken_res_39 = _RANDOM[4'h5][7];
        useV0AsMaskToken_res_40 = _RANDOM[4'h5][8];
        useV0AsMaskToken_res_41 = _RANDOM[4'h5][9];
        useV0AsMaskToken_res_42 = _RANDOM[4'h5][10];
        useV0AsMaskToken_res_43 = _RANDOM[4'h5][11];
        useV0AsMaskToken_res_44 = _RANDOM[4'h5][12];
        useV0AsMaskToken_res_45 = _RANDOM[4'h5][13];
        useV0AsMaskToken_res_46 = _RANDOM[4'h5][14];
        useV0AsMaskToken_res_47 = _RANDOM[4'h5][15];
        useV0AsMaskToken_res_48 = _RANDOM[4'h5][16];
        useV0AsMaskToken_res_49 = _RANDOM[4'h5][17];
        useV0AsMaskToken_res_50 = _RANDOM[4'h5][18];
        useV0AsMaskToken_res_51 = _RANDOM[4'h5][19];
        useV0AsMaskToken_res_52 = _RANDOM[4'h5][20];
        useV0AsMaskToken_res_53 = _RANDOM[4'h5][21];
        useV0AsMaskToken_res_54 = _RANDOM[4'h5][22];
        useV0AsMaskToken_res_55 = _RANDOM[4'h5][23];
        useV0AsMaskToken_res_56 = _RANDOM[4'h5][24];
        useV0AsMaskToken_res_57 = _RANDOM[4'h5][25];
        useV0AsMaskToken_res_58 = _RANDOM[4'h5][26];
        useV0AsMaskToken_res_59 = _RANDOM[4'h5][27];
        useV0AsMaskToken_res_60 = _RANDOM[4'h5][28];
        useV0AsMaskToken_res_61 = _RANDOM[4'h5][29];
        useV0AsMaskToken_res_62 = _RANDOM[4'h5][30];
        useV0AsMaskToken_res_63 = _RANDOM[4'h5][31];
        useV0AsMaskToken_res_64 = _RANDOM[4'h6][0];
        useV0AsMaskToken_res_65 = _RANDOM[4'h6][1];
        useV0AsMaskToken_res_66 = _RANDOM[4'h6][2];
        useV0AsMaskToken_res_67 = _RANDOM[4'h6][3];
        useV0AsMaskToken_res_68 = _RANDOM[4'h6][4];
        useV0AsMaskToken_res_69 = _RANDOM[4'h6][5];
        useV0AsMaskToken_res_70 = _RANDOM[4'h6][6];
        useV0AsMaskToken_res_71 = _RANDOM[4'h6][7];
        useV0AsMaskToken_res_72 = _RANDOM[4'h6][8];
        useV0AsMaskToken_res_73 = _RANDOM[4'h6][9];
        useV0AsMaskToken_res_74 = _RANDOM[4'h6][10];
        useV0AsMaskToken_res_75 = _RANDOM[4'h6][11];
        useV0AsMaskToken_res_76 = _RANDOM[4'h6][12];
        useV0AsMaskToken_res_77 = _RANDOM[4'h6][13];
        useV0AsMaskToken_res_78 = _RANDOM[4'h6][14];
        useV0AsMaskToken_res_79 = _RANDOM[4'h6][15];
        useV0AsMaskToken_res_80 = _RANDOM[4'h6][16];
        useV0AsMaskToken_res_81 = _RANDOM[4'h6][17];
        useV0AsMaskToken_res_82 = _RANDOM[4'h6][18];
        useV0AsMaskToken_res_83 = _RANDOM[4'h6][19];
        useV0AsMaskToken_res_84 = _RANDOM[4'h6][20];
        useV0AsMaskToken_res_85 = _RANDOM[4'h6][21];
        useV0AsMaskToken_res_86 = _RANDOM[4'h6][22];
        useV0AsMaskToken_res_87 = _RANDOM[4'h6][23];
        useV0AsMaskToken_res_88 = _RANDOM[4'h6][24];
        useV0AsMaskToken_res_89 = _RANDOM[4'h6][25];
        useV0AsMaskToken_res_90 = _RANDOM[4'h6][26];
        useV0AsMaskToken_res_91 = _RANDOM[4'h6][27];
        useV0AsMaskToken_res_92 = _RANDOM[4'h6][28];
        useV0AsMaskToken_res_93 = _RANDOM[4'h6][29];
        useV0AsMaskToken_res_94 = _RANDOM[4'h6][30];
        useV0AsMaskToken_res_95 = _RANDOM[4'h6][31];
        useV0AsMaskToken_res_96 = _RANDOM[4'h7][0];
        useV0AsMaskToken_res_97 = _RANDOM[4'h7][1];
        useV0AsMaskToken_res_98 = _RANDOM[4'h7][2];
        useV0AsMaskToken_res_99 = _RANDOM[4'h7][3];
        useV0AsMaskToken_res_100 = _RANDOM[4'h7][4];
        useV0AsMaskToken_res_101 = _RANDOM[4'h7][5];
        useV0AsMaskToken_res_102 = _RANDOM[4'h7][6];
        useV0AsMaskToken_res_103 = _RANDOM[4'h7][7];
        useV0AsMaskToken_res_104 = _RANDOM[4'h7][8];
        useV0AsMaskToken_res_105 = _RANDOM[4'h7][9];
        useV0AsMaskToken_res_106 = _RANDOM[4'h7][10];
        useV0AsMaskToken_res_107 = _RANDOM[4'h7][11];
        useV0AsMaskToken_res_108 = _RANDOM[4'h7][12];
        useV0AsMaskToken_res_109 = _RANDOM[4'h7][13];
        useV0AsMaskToken_res_110 = _RANDOM[4'h7][14];
        useV0AsMaskToken_res_111 = _RANDOM[4'h7][15];
        useV0AsMaskToken_res_112 = _RANDOM[4'h7][16];
        useV0AsMaskToken_res_113 = _RANDOM[4'h7][17];
        useV0AsMaskToken_res_114 = _RANDOM[4'h7][18];
        useV0AsMaskToken_res_115 = _RANDOM[4'h7][19];
        useV0AsMaskToken_res_116 = _RANDOM[4'h7][20];
        useV0AsMaskToken_res_117 = _RANDOM[4'h7][21];
        useV0AsMaskToken_res_118 = _RANDOM[4'h7][22];
        useV0AsMaskToken_res_119 = _RANDOM[4'h7][23];
        useV0AsMaskToken_res_120 = _RANDOM[4'h7][24];
        useV0AsMaskToken_res_121 = _RANDOM[4'h7][25];
        useV0AsMaskToken_res_122 = _RANDOM[4'h7][26];
        useV0AsMaskToken_res_123 = _RANDOM[4'h7][27];
        useV0AsMaskToken_res_124 = _RANDOM[4'h7][28];
        useV0AsMaskToken_res_125 = _RANDOM[4'h7][29];
        useV0AsMaskToken_res_126 = _RANDOM[4'h7][30];
        useV0AsMaskToken_res_127 = _RANDOM[4'h7][31];
        maskUnitWriteV0 = _RANDOM[4'h8][0];
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  assign issueAllow = ~v0Conflict;
  assign v0WriteValid = _v0WriteValid_output;
endmodule

