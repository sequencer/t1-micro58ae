
// Include register initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for register randomization.

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_
module MaskUnit(
  input         clock,
                reset,
                instReq_valid,
  input  [2:0]  instReq_bits_instructionIndex,
  input         instReq_bits_decodeResult_specialSlot,
  input  [4:0]  instReq_bits_decodeResult_topUop,
  input         instReq_bits_decodeResult_popCount,
                instReq_bits_decodeResult_ffo,
                instReq_bits_decodeResult_average,
                instReq_bits_decodeResult_reverse,
                instReq_bits_decodeResult_dontNeedExecuteInLane,
                instReq_bits_decodeResult_scheduler,
                instReq_bits_decodeResult_sReadVD,
                instReq_bits_decodeResult_vtype,
                instReq_bits_decodeResult_sWrite,
                instReq_bits_decodeResult_crossRead,
                instReq_bits_decodeResult_crossWrite,
                instReq_bits_decodeResult_maskUnit,
                instReq_bits_decodeResult_special,
                instReq_bits_decodeResult_saturate,
                instReq_bits_decodeResult_vwmacc,
                instReq_bits_decodeResult_readOnly,
                instReq_bits_decodeResult_maskSource,
                instReq_bits_decodeResult_maskDestination,
                instReq_bits_decodeResult_maskLogic,
  input  [3:0]  instReq_bits_decodeResult_uop,
  input         instReq_bits_decodeResult_iota,
                instReq_bits_decodeResult_mv,
                instReq_bits_decodeResult_extend,
                instReq_bits_decodeResult_unOrderWrite,
                instReq_bits_decodeResult_compress,
                instReq_bits_decodeResult_gather16,
                instReq_bits_decodeResult_gather,
                instReq_bits_decodeResult_slid,
                instReq_bits_decodeResult_targetRd,
                instReq_bits_decodeResult_widenReduce,
                instReq_bits_decodeResult_red,
                instReq_bits_decodeResult_nr,
                instReq_bits_decodeResult_itype,
                instReq_bits_decodeResult_unsigned1,
                instReq_bits_decodeResult_unsigned0,
                instReq_bits_decodeResult_other,
                instReq_bits_decodeResult_multiCycle,
                instReq_bits_decodeResult_divider,
                instReq_bits_decodeResult_multiplier,
                instReq_bits_decodeResult_shift,
                instReq_bits_decodeResult_adder,
                instReq_bits_decodeResult_logic,
  input  [31:0] instReq_bits_readFromScala,
  input  [1:0]  instReq_bits_sew,
  input  [2:0]  instReq_bits_vlmul,
  input         instReq_bits_maskType,
  input  [2:0]  instReq_bits_vxrm,
  input  [4:0]  instReq_bits_vs2,
                instReq_bits_vs1,
                instReq_bits_vd,
  input  [8:0]  instReq_bits_vl,
  input         exeReq_0_valid,
  input  [31:0] exeReq_0_bits_source1,
                exeReq_0_bits_source2,
  input  [2:0]  exeReq_0_bits_index,
  input         exeReq_0_bits_ffo,
                exeReq_1_valid,
  input  [31:0] exeReq_1_bits_source1,
                exeReq_1_bits_source2,
  input  [2:0]  exeReq_1_bits_index,
  input         exeReq_1_bits_ffo,
                exeReq_2_valid,
  input  [31:0] exeReq_2_bits_source1,
                exeReq_2_bits_source2,
  input  [2:0]  exeReq_2_bits_index,
  input         exeReq_2_bits_ffo,
                exeReq_3_valid,
  input  [31:0] exeReq_3_bits_source1,
                exeReq_3_bits_source2,
  input  [2:0]  exeReq_3_bits_index,
  input         exeReq_3_bits_ffo,
                exeResp_0_ready,
  output        exeResp_0_valid,
  output [4:0]  exeResp_0_bits_vd,
  output        exeResp_0_bits_offset,
  output [3:0]  exeResp_0_bits_mask,
  output [31:0] exeResp_0_bits_data,
  output [2:0]  exeResp_0_bits_instructionIndex,
  input         exeResp_1_ready,
  output        exeResp_1_valid,
  output [4:0]  exeResp_1_bits_vd,
  output        exeResp_1_bits_offset,
  output [3:0]  exeResp_1_bits_mask,
  output [31:0] exeResp_1_bits_data,
  output [2:0]  exeResp_1_bits_instructionIndex,
  input         exeResp_2_ready,
  output        exeResp_2_valid,
  output [4:0]  exeResp_2_bits_vd,
  output        exeResp_2_bits_offset,
  output [3:0]  exeResp_2_bits_mask,
  output [31:0] exeResp_2_bits_data,
  output [2:0]  exeResp_2_bits_instructionIndex,
  input         exeResp_3_ready,
  output        exeResp_3_valid,
  output [4:0]  exeResp_3_bits_vd,
  output        exeResp_3_bits_offset,
  output [3:0]  exeResp_3_bits_mask,
  output [31:0] exeResp_3_bits_data,
  output [2:0]  exeResp_3_bits_instructionIndex,
  input         writeRelease_0,
                writeRelease_1,
                writeRelease_2,
                writeRelease_3,
  output        tokenIO_0_maskRequestRelease,
                tokenIO_1_maskRequestRelease,
                tokenIO_2_maskRequestRelease,
                tokenIO_3_maskRequestRelease,
  input         readChannel_0_ready,
  output        readChannel_0_valid,
  output [4:0]  readChannel_0_bits_vs,
  output        readChannel_0_bits_offset,
  output [2:0]  readChannel_0_bits_instructionIndex,
  input         readChannel_1_ready,
  output        readChannel_1_valid,
  output [4:0]  readChannel_1_bits_vs,
  output        readChannel_1_bits_offset,
  output [2:0]  readChannel_1_bits_instructionIndex,
  input         readChannel_2_ready,
  output        readChannel_2_valid,
  output [4:0]  readChannel_2_bits_vs,
  output        readChannel_2_bits_offset,
  output [2:0]  readChannel_2_bits_instructionIndex,
  input         readChannel_3_ready,
  output        readChannel_3_valid,
  output [4:0]  readChannel_3_bits_vs,
  output        readChannel_3_bits_offset,
  output [2:0]  readChannel_3_bits_instructionIndex,
  input         readResult_0_valid,
  input  [31:0] readResult_0_bits,
  input         readResult_1_valid,
  input  [31:0] readResult_1_bits,
  input         readResult_2_valid,
  input  [31:0] readResult_2_bits,
  input         readResult_3_valid,
  input  [31:0] readResult_3_bits,
  output [7:0]  lastReport,
  output [31:0] laneMaskInput_0,
                laneMaskInput_1,
                laneMaskInput_2,
                laneMaskInput_3,
  input  [2:0]  laneMaskSelect_0,
                laneMaskSelect_1,
                laneMaskSelect_2,
                laneMaskSelect_3,
  input  [1:0]  laneMaskSewSelect_0,
                laneMaskSewSelect_1,
                laneMaskSewSelect_2,
                laneMaskSewSelect_3,
  input         v0UpdateVec_0_valid,
  input  [31:0] v0UpdateVec_0_bits_data,
  input         v0UpdateVec_0_bits_offset,
  input  [3:0]  v0UpdateVec_0_bits_mask,
  input         v0UpdateVec_1_valid,
  input  [31:0] v0UpdateVec_1_bits_data,
  input         v0UpdateVec_1_bits_offset,
  input  [3:0]  v0UpdateVec_1_bits_mask,
  input         v0UpdateVec_2_valid,
  input  [31:0] v0UpdateVec_2_bits_data,
  input         v0UpdateVec_2_bits_offset,
  input  [3:0]  v0UpdateVec_2_bits_mask,
  input         v0UpdateVec_3_valid,
  input  [31:0] v0UpdateVec_3_bits_data,
  input         v0UpdateVec_3_bits_offset,
  input  [3:0]  v0UpdateVec_3_bits_mask,
  output [31:0] writeRDData,
  input         gatherData_ready,
  output        gatherData_valid,
  output [31:0] gatherData_bits,
  input         gatherRead
);

  wire              readCrossBar_input_3_valid;
  wire              readCrossBar_input_2_valid;
  wire              readCrossBar_input_1_valid;
  wire              readCrossBar_input_0_valid;
  wire              _writeQueue_fifo_3_empty;
  wire              _writeQueue_fifo_3_full;
  wire              _writeQueue_fifo_3_error;
  wire [49:0]       _writeQueue_fifo_3_data_out;
  wire              _writeQueue_fifo_2_empty;
  wire              _writeQueue_fifo_2_full;
  wire              _writeQueue_fifo_2_error;
  wire [49:0]       _writeQueue_fifo_2_data_out;
  wire              _writeQueue_fifo_1_empty;
  wire              _writeQueue_fifo_1_full;
  wire              _writeQueue_fifo_1_error;
  wire [49:0]       _writeQueue_fifo_1_data_out;
  wire              _writeQueue_fifo_empty;
  wire              _writeQueue_fifo_full;
  wire              _writeQueue_fifo_error;
  wire [49:0]       _writeQueue_fifo_data_out;
  wire [127:0]      _extendUnit_out;
  wire              _reduceUnit_in_ready;
  wire              _reduceUnit_out_valid;
  wire [31:0]       _reduceUnit_out_bits_data;
  wire [3:0]        _reduceUnit_out_bits_mask;
  wire              _compressUnit_out_compressValid;
  wire [31:0]       _compressUnit_writeData;
  wire              _compressUnit_stageValid;
  wire              _readData_readDataQueue_fifo_3_empty;
  wire              _readData_readDataQueue_fifo_3_full;
  wire              _readData_readDataQueue_fifo_3_error;
  wire [31:0]       _readData_readDataQueue_fifo_3_data_out;
  wire              _readData_readDataQueue_fifo_2_empty;
  wire              _readData_readDataQueue_fifo_2_full;
  wire              _readData_readDataQueue_fifo_2_error;
  wire [31:0]       _readData_readDataQueue_fifo_2_data_out;
  wire              _readData_readDataQueue_fifo_1_empty;
  wire              _readData_readDataQueue_fifo_1_full;
  wire              _readData_readDataQueue_fifo_1_error;
  wire [31:0]       _readData_readDataQueue_fifo_1_data_out;
  wire              _readData_readDataQueue_fifo_empty;
  wire              _readData_readDataQueue_fifo_full;
  wire              _readData_readDataQueue_fifo_error;
  wire [31:0]       _readData_readDataQueue_fifo_data_out;
  wire              _readMessageQueue_fifo_3_empty;
  wire              _readMessageQueue_fifo_3_full;
  wire              _readMessageQueue_fifo_3_error;
  wire [5:0]        _readMessageQueue_fifo_3_data_out;
  wire              _readMessageQueue_fifo_2_empty;
  wire              _readMessageQueue_fifo_2_full;
  wire              _readMessageQueue_fifo_2_error;
  wire [5:0]        _readMessageQueue_fifo_2_data_out;
  wire              _readMessageQueue_fifo_1_empty;
  wire              _readMessageQueue_fifo_1_full;
  wire              _readMessageQueue_fifo_1_error;
  wire [5:0]        _readMessageQueue_fifo_1_data_out;
  wire              _readMessageQueue_fifo_empty;
  wire              _readMessageQueue_fifo_full;
  wire              _readMessageQueue_fifo_error;
  wire [5:0]        _readMessageQueue_fifo_data_out;
  wire              _reorderQueueVec_fifo_3_empty;
  wire              _reorderQueueVec_fifo_3_full;
  wire              _reorderQueueVec_fifo_3_error;
  wire [35:0]       _reorderQueueVec_fifo_3_data_out;
  wire              _reorderQueueVec_fifo_2_empty;
  wire              _reorderQueueVec_fifo_2_full;
  wire              _reorderQueueVec_fifo_2_error;
  wire [35:0]       _reorderQueueVec_fifo_2_data_out;
  wire              _reorderQueueVec_fifo_1_empty;
  wire              _reorderQueueVec_fifo_1_full;
  wire              _reorderQueueVec_fifo_1_error;
  wire [35:0]       _reorderQueueVec_fifo_1_data_out;
  wire              _reorderQueueVec_fifo_empty;
  wire              _reorderQueueVec_fifo_full;
  wire              _reorderQueueVec_fifo_error;
  wire [35:0]       _reorderQueueVec_fifo_data_out;
  wire              _compressUnitResultQueue_fifo_empty;
  wire              _compressUnitResultQueue_fifo_full;
  wire              _compressUnitResultQueue_fifo_error;
  wire [153:0]      _compressUnitResultQueue_fifo_data_out;
  wire              _readWaitQueue_fifo_empty;
  wire              _readWaitQueue_fifo_full;
  wire              _readWaitQueue_fifo_error;
  wire [19:0]       _readWaitQueue_fifo_data_out;
  wire              _readCrossBar_input_0_ready;
  wire              _readCrossBar_input_1_ready;
  wire              _readCrossBar_input_2_ready;
  wire              _readCrossBar_input_3_ready;
  wire              _readCrossBar_output_0_valid;
  wire [4:0]        _readCrossBar_output_0_bits_vs;
  wire              _readCrossBar_output_0_bits_offset;
  wire [1:0]        _readCrossBar_output_0_bits_writeIndex;
  wire              _readCrossBar_output_1_valid;
  wire [4:0]        _readCrossBar_output_1_bits_vs;
  wire              _readCrossBar_output_1_bits_offset;
  wire [1:0]        _readCrossBar_output_1_bits_writeIndex;
  wire              _readCrossBar_output_2_valid;
  wire [4:0]        _readCrossBar_output_2_bits_vs;
  wire              _readCrossBar_output_2_bits_offset;
  wire [1:0]        _readCrossBar_output_2_bits_writeIndex;
  wire              _readCrossBar_output_3_valid;
  wire [4:0]        _readCrossBar_output_3_bits_vs;
  wire              _readCrossBar_output_3_bits_offset;
  wire [1:0]        _readCrossBar_output_3_bits_writeIndex;
  wire              _accessCountQueue_fifo_empty;
  wire              _accessCountQueue_fifo_full;
  wire              _accessCountQueue_fifo_error;
  wire [11:0]       _accessCountQueue_fifo_data_out;
  wire              _slideAddressGen_indexDeq_valid;
  wire [3:0]        _slideAddressGen_indexDeq_bits_needRead;
  wire [3:0]        _slideAddressGen_indexDeq_bits_elementValid;
  wire [3:0]        _slideAddressGen_indexDeq_bits_replaceVs1;
  wire [3:0]        _slideAddressGen_indexDeq_bits_readOffset;
  wire [1:0]        _slideAddressGen_indexDeq_bits_accessLane_0;
  wire [1:0]        _slideAddressGen_indexDeq_bits_accessLane_1;
  wire [1:0]        _slideAddressGen_indexDeq_bits_accessLane_2;
  wire [1:0]        _slideAddressGen_indexDeq_bits_accessLane_3;
  wire [2:0]        _slideAddressGen_indexDeq_bits_vsGrowth_0;
  wire [2:0]        _slideAddressGen_indexDeq_bits_vsGrowth_1;
  wire [2:0]        _slideAddressGen_indexDeq_bits_vsGrowth_2;
  wire [2:0]        _slideAddressGen_indexDeq_bits_vsGrowth_3;
  wire [6:0]        _slideAddressGen_indexDeq_bits_executeGroup;
  wire [7:0]        _slideAddressGen_indexDeq_bits_readDataOffset;
  wire              _slideAddressGen_indexDeq_bits_last;
  wire [6:0]        _slideAddressGen_slideGroupOut;
  wire              _exeRequestQueue_queue_fifo_3_empty;
  wire              _exeRequestQueue_queue_fifo_3_full;
  wire              _exeRequestQueue_queue_fifo_3_error;
  wire [67:0]       _exeRequestQueue_queue_fifo_3_data_out;
  wire              _exeRequestQueue_queue_fifo_2_empty;
  wire              _exeRequestQueue_queue_fifo_2_full;
  wire              _exeRequestQueue_queue_fifo_2_error;
  wire [67:0]       _exeRequestQueue_queue_fifo_2_data_out;
  wire              _exeRequestQueue_queue_fifo_1_empty;
  wire              _exeRequestQueue_queue_fifo_1_full;
  wire              _exeRequestQueue_queue_fifo_1_error;
  wire [67:0]       _exeRequestQueue_queue_fifo_1_data_out;
  wire              _exeRequestQueue_queue_fifo_empty;
  wire              _exeRequestQueue_queue_fifo_full;
  wire              _exeRequestQueue_queue_fifo_error;
  wire [67:0]       _exeRequestQueue_queue_fifo_data_out;
  wire              _maskedWrite_in_0_ready;
  wire              _maskedWrite_in_1_ready;
  wire              _maskedWrite_in_2_ready;
  wire              _maskedWrite_in_3_ready;
  wire              _maskedWrite_out_0_valid;
  wire              _maskedWrite_out_0_bits_ffoByOther;
  wire [31:0]       _maskedWrite_out_0_bits_writeData_data;
  wire [3:0]        _maskedWrite_out_0_bits_writeData_mask;
  wire [4:0]        _maskedWrite_out_0_bits_writeData_groupCounter;
  wire              _maskedWrite_out_1_valid;
  wire              _maskedWrite_out_1_bits_ffoByOther;
  wire [31:0]       _maskedWrite_out_1_bits_writeData_data;
  wire [3:0]        _maskedWrite_out_1_bits_writeData_mask;
  wire [4:0]        _maskedWrite_out_1_bits_writeData_groupCounter;
  wire              _maskedWrite_out_2_valid;
  wire              _maskedWrite_out_2_bits_ffoByOther;
  wire [31:0]       _maskedWrite_out_2_bits_writeData_data;
  wire [3:0]        _maskedWrite_out_2_bits_writeData_mask;
  wire [4:0]        _maskedWrite_out_2_bits_writeData_groupCounter;
  wire              _maskedWrite_out_3_valid;
  wire              _maskedWrite_out_3_bits_ffoByOther;
  wire [31:0]       _maskedWrite_out_3_bits_writeData_data;
  wire [3:0]        _maskedWrite_out_3_bits_writeData_mask;
  wire [4:0]        _maskedWrite_out_3_bits_writeData_groupCounter;
  wire              _maskedWrite_readChannel_0_valid;
  wire [4:0]        _maskedWrite_readChannel_0_bits_vs;
  wire              _maskedWrite_readChannel_0_bits_offset;
  wire              _maskedWrite_readChannel_1_valid;
  wire [4:0]        _maskedWrite_readChannel_1_bits_vs;
  wire              _maskedWrite_readChannel_1_bits_offset;
  wire              _maskedWrite_readChannel_2_valid;
  wire [4:0]        _maskedWrite_readChannel_2_bits_vs;
  wire              _maskedWrite_readChannel_2_bits_offset;
  wire              _maskedWrite_readChannel_3_valid;
  wire [4:0]        _maskedWrite_readChannel_3_bits_vs;
  wire              _maskedWrite_readChannel_3_bits_offset;
  wire              _maskedWrite_stageClear;
  wire              writeQueue_3_almostFull;
  wire              writeQueue_3_almostEmpty;
  wire              writeQueue_2_almostFull;
  wire              writeQueue_2_almostEmpty;
  wire              writeQueue_1_almostFull;
  wire              writeQueue_1_almostEmpty;
  wire              writeQueue_0_almostFull;
  wire              writeQueue_0_almostEmpty;
  wire              readData_readDataQueue_3_almostFull;
  wire              readData_readDataQueue_3_almostEmpty;
  wire              readData_readDataQueue_2_almostFull;
  wire              readData_readDataQueue_2_almostEmpty;
  wire              readData_readDataQueue_1_almostFull;
  wire              readData_readDataQueue_1_almostEmpty;
  wire              readData_readDataQueue_almostFull;
  wire              readData_readDataQueue_almostEmpty;
  wire              readMessageQueue_3_almostFull;
  wire              readMessageQueue_3_almostEmpty;
  wire              readMessageQueue_2_almostFull;
  wire              readMessageQueue_2_almostEmpty;
  wire              readMessageQueue_1_almostFull;
  wire              readMessageQueue_1_almostEmpty;
  wire              readMessageQueue_almostFull;
  wire              readMessageQueue_almostEmpty;
  wire              reorderQueueVec_3_almostFull;
  wire              reorderQueueVec_3_almostEmpty;
  wire              reorderQueueVec_2_almostFull;
  wire              reorderQueueVec_2_almostEmpty;
  wire              reorderQueueVec_1_almostFull;
  wire              reorderQueueVec_1_almostEmpty;
  wire              reorderQueueVec_0_almostFull;
  wire              reorderQueueVec_0_almostEmpty;
  wire              compressUnitResultQueue_almostFull;
  wire              compressUnitResultQueue_almostEmpty;
  wire              readWaitQueue_almostFull;
  wire              readWaitQueue_almostEmpty;
  wire              accessCountQueue_almostFull;
  wire              accessCountQueue_almostEmpty;
  wire              exeRequestQueue_3_almostFull;
  wire              exeRequestQueue_3_almostEmpty;
  wire              exeRequestQueue_2_almostFull;
  wire              exeRequestQueue_2_almostEmpty;
  wire              exeRequestQueue_1_almostFull;
  wire              exeRequestQueue_1_almostEmpty;
  wire              exeRequestQueue_0_almostFull;
  wire              exeRequestQueue_0_almostEmpty;
  wire [31:0]       reorderQueueVec_3_deq_bits_data;
  wire [31:0]       reorderQueueVec_2_deq_bits_data;
  wire [31:0]       reorderQueueVec_1_deq_bits_data;
  wire [31:0]       reorderQueueVec_0_deq_bits_data;
  wire [2:0]        accessCountEnq_3;
  wire [2:0]        accessCountEnq_2;
  wire [2:0]        accessCountEnq_1;
  wire [2:0]        accessCountEnq_0;
  wire              exeResp_0_ready_0 = exeResp_0_ready;
  wire              exeResp_1_ready_0 = exeResp_1_ready;
  wire              exeResp_2_ready_0 = exeResp_2_ready;
  wire              exeResp_3_ready_0 = exeResp_3_ready;
  wire              readChannel_0_ready_0 = readChannel_0_ready;
  wire              readChannel_1_ready_0 = readChannel_1_ready;
  wire              readChannel_2_ready_0 = readChannel_2_ready;
  wire              readChannel_3_ready_0 = readChannel_3_ready;
  wire              gatherData_ready_0 = gatherData_ready;
  wire              exeRequestQueue_0_enq_valid = exeReq_0_valid;
  wire [31:0]       exeRequestQueue_0_enq_bits_source1 = exeReq_0_bits_source1;
  wire [31:0]       exeRequestQueue_0_enq_bits_source2 = exeReq_0_bits_source2;
  wire [2:0]        exeRequestQueue_0_enq_bits_index = exeReq_0_bits_index;
  wire              exeRequestQueue_0_enq_bits_ffo = exeReq_0_bits_ffo;
  wire              exeRequestQueue_1_enq_valid = exeReq_1_valid;
  wire [31:0]       exeRequestQueue_1_enq_bits_source1 = exeReq_1_bits_source1;
  wire [31:0]       exeRequestQueue_1_enq_bits_source2 = exeReq_1_bits_source2;
  wire [2:0]        exeRequestQueue_1_enq_bits_index = exeReq_1_bits_index;
  wire              exeRequestQueue_1_enq_bits_ffo = exeReq_1_bits_ffo;
  wire              exeRequestQueue_2_enq_valid = exeReq_2_valid;
  wire [31:0]       exeRequestQueue_2_enq_bits_source1 = exeReq_2_bits_source1;
  wire [31:0]       exeRequestQueue_2_enq_bits_source2 = exeReq_2_bits_source2;
  wire [2:0]        exeRequestQueue_2_enq_bits_index = exeReq_2_bits_index;
  wire              exeRequestQueue_2_enq_bits_ffo = exeReq_2_bits_ffo;
  wire              exeRequestQueue_3_enq_valid = exeReq_3_valid;
  wire [31:0]       exeRequestQueue_3_enq_bits_source1 = exeReq_3_bits_source1;
  wire [31:0]       exeRequestQueue_3_enq_bits_source2 = exeReq_3_bits_source2;
  wire [2:0]        exeRequestQueue_3_enq_bits_index = exeReq_3_bits_index;
  wire              exeRequestQueue_3_enq_bits_ffo = exeReq_3_bits_ffo;
  wire              reorderQueueVec_0_enq_valid = readResult_0_valid;
  wire              reorderQueueVec_1_enq_valid = readResult_1_valid;
  wire              reorderQueueVec_2_enq_valid = readResult_2_valid;
  wire              reorderQueueVec_3_enq_valid = readResult_3_valid;
  wire              readMessageQueue_deq_ready = readResult_0_valid;
  wire              readMessageQueue_1_deq_ready = readResult_1_valid;
  wire              readMessageQueue_2_deq_ready = readResult_2_valid;
  wire              readMessageQueue_3_deq_ready = readResult_3_valid;
  wire [7:0]        checkVec_checkResult_lo_14 = 8'hFF;
  wire [7:0]        checkVec_checkResult_hi_14 = 8'hFF;
  wire [15:0]       checkVec_2_0 = 16'hFFFF;
  wire [7:0]        checkVec_2_1 = 8'h0;
  wire [1:0]        readVS1Req_requestIndex = 2'h0;
  wire [1:0]        checkVec_checkResultVec_0_1_2 = 2'h0;
  wire [1:0]        checkVec_checkResultVec_1_1_2 = 2'h0;
  wire [1:0]        checkVec_checkResultVec_2_1_2 = 2'h0;
  wire [1:0]        checkVec_checkResultVec_3_1_2 = 2'h0;
  wire [1:0]        selectExecuteReq_0_bits_requestIndex = 2'h0;
  wire [1:0]        selectExecuteReq_1_bits_requestIndex = 2'h1;
  wire [1:0]        selectExecuteReq_3_bits_requestIndex = 2'h3;
  wire [3:0]        checkVec_checkResult_lo_15 = 4'h0;
  wire [3:0]        checkVec_checkResult_hi_15 = 4'h0;
  wire [1:0]        readChannel_0_bits_readSource = 2'h2;
  wire [1:0]        readChannel_1_bits_readSource = 2'h2;
  wire [1:0]        readChannel_2_bits_readSource = 2'h2;
  wire [1:0]        readChannel_3_bits_readSource = 2'h2;
  wire [1:0]        selectExecuteReq_2_bits_requestIndex = 2'h2;
  wire              exeResp_0_bits_last = 1'h0;
  wire              exeResp_1_bits_last = 1'h0;
  wire              exeResp_2_bits_last = 1'h0;
  wire              exeResp_3_bits_last = 1'h0;
  wire              writeRequest_0_ffoByOther = 1'h0;
  wire              writeRequest_1_ffoByOther = 1'h0;
  wire              writeRequest_2_ffoByOther = 1'h0;
  wire              writeRequest_3_ffoByOther = 1'h0;
  wire              writeQueue_0_deq_ready = exeResp_0_ready_0;
  wire              writeQueue_0_deq_valid;
  wire [3:0]        writeQueue_0_deq_bits_writeData_mask;
  wire [31:0]       writeQueue_0_deq_bits_writeData_data;
  wire              writeQueue_1_deq_ready = exeResp_1_ready_0;
  wire              writeQueue_1_deq_valid;
  wire [3:0]        writeQueue_1_deq_bits_writeData_mask;
  wire [31:0]       writeQueue_1_deq_bits_writeData_data;
  wire              writeQueue_2_deq_ready = exeResp_2_ready_0;
  wire              writeQueue_2_deq_valid;
  wire [3:0]        writeQueue_2_deq_bits_writeData_mask;
  wire [31:0]       writeQueue_2_deq_bits_writeData_data;
  wire              writeQueue_3_deq_ready = exeResp_3_ready_0;
  wire              writeQueue_3_deq_valid;
  wire [3:0]        writeQueue_3_deq_bits_writeData_mask;
  wire [31:0]       writeQueue_3_deq_bits_writeData_data;
  wire              gatherResponse;
  reg  [31:0]       v0_0;
  reg  [31:0]       v0_1;
  reg  [31:0]       v0_2;
  reg  [31:0]       v0_3;
  reg  [31:0]       v0_4;
  reg  [31:0]       v0_5;
  reg  [31:0]       v0_6;
  reg  [31:0]       v0_7;
  wire [15:0]       maskExt_lo = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]       maskExt_hi = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]       maskExt = {maskExt_hi, maskExt_lo};
  wire [15:0]       maskExt_lo_1 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_1 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]       maskExt_1 = {maskExt_hi_1, maskExt_lo_1};
  wire [15:0]       maskExt_lo_2 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_2 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]       maskExt_2 = {maskExt_hi_2, maskExt_lo_2};
  wire [15:0]       maskExt_lo_3 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_3 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]       maskExt_3 = {maskExt_hi_3, maskExt_lo_3};
  wire [15:0]       maskExt_lo_4 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_4 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]       maskExt_4 = {maskExt_hi_4, maskExt_lo_4};
  wire [15:0]       maskExt_lo_5 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_5 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]       maskExt_5 = {maskExt_hi_5, maskExt_lo_5};
  wire [15:0]       maskExt_lo_6 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_6 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]       maskExt_6 = {maskExt_hi_6, maskExt_lo_6};
  wire [15:0]       maskExt_lo_7 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_7 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]       maskExt_7 = {maskExt_hi_7, maskExt_lo_7};
  wire [63:0]       _GEN = {v0_1, v0_0};
  wire [63:0]       regroupV0_lo_lo;
  assign regroupV0_lo_lo = _GEN;
  wire [63:0]       regroupV0_lo_lo_5;
  assign regroupV0_lo_lo_5 = _GEN;
  wire [63:0]       regroupV0_lo_lo_10;
  assign regroupV0_lo_lo_10 = _GEN;
  wire [63:0]       slideAddressGen_slideMaskInput_lo_lo;
  assign slideAddressGen_slideMaskInput_lo_lo = _GEN;
  wire [63:0]       selectReadStageMask_lo_lo;
  assign selectReadStageMask_lo_lo = _GEN;
  wire [63:0]       maskSplit_maskSelect_lo_lo;
  assign maskSplit_maskSelect_lo_lo = _GEN;
  wire [63:0]       maskSplit_maskSelect_lo_lo_1;
  assign maskSplit_maskSelect_lo_lo_1 = _GEN;
  wire [63:0]       maskSplit_maskSelect_lo_lo_2;
  assign maskSplit_maskSelect_lo_lo_2 = _GEN;
  wire [63:0]       maskForDestination_lo_lo;
  assign maskForDestination_lo_lo = _GEN;
  wire [63:0]       _GEN_0 = {v0_3, v0_2};
  wire [63:0]       regroupV0_lo_hi;
  assign regroupV0_lo_hi = _GEN_0;
  wire [63:0]       regroupV0_lo_hi_5;
  assign regroupV0_lo_hi_5 = _GEN_0;
  wire [63:0]       regroupV0_lo_hi_10;
  assign regroupV0_lo_hi_10 = _GEN_0;
  wire [63:0]       slideAddressGen_slideMaskInput_lo_hi;
  assign slideAddressGen_slideMaskInput_lo_hi = _GEN_0;
  wire [63:0]       selectReadStageMask_lo_hi;
  assign selectReadStageMask_lo_hi = _GEN_0;
  wire [63:0]       maskSplit_maskSelect_lo_hi;
  assign maskSplit_maskSelect_lo_hi = _GEN_0;
  wire [63:0]       maskSplit_maskSelect_lo_hi_1;
  assign maskSplit_maskSelect_lo_hi_1 = _GEN_0;
  wire [63:0]       maskSplit_maskSelect_lo_hi_2;
  assign maskSplit_maskSelect_lo_hi_2 = _GEN_0;
  wire [63:0]       maskForDestination_lo_hi;
  assign maskForDestination_lo_hi = _GEN_0;
  wire [127:0]      regroupV0_lo = {regroupV0_lo_hi, regroupV0_lo_lo};
  wire [63:0]       _GEN_1 = {v0_5, v0_4};
  wire [63:0]       regroupV0_hi_lo;
  assign regroupV0_hi_lo = _GEN_1;
  wire [63:0]       regroupV0_hi_lo_5;
  assign regroupV0_hi_lo_5 = _GEN_1;
  wire [63:0]       regroupV0_hi_lo_10;
  assign regroupV0_hi_lo_10 = _GEN_1;
  wire [63:0]       slideAddressGen_slideMaskInput_hi_lo;
  assign slideAddressGen_slideMaskInput_hi_lo = _GEN_1;
  wire [63:0]       selectReadStageMask_hi_lo;
  assign selectReadStageMask_hi_lo = _GEN_1;
  wire [63:0]       maskSplit_maskSelect_hi_lo;
  assign maskSplit_maskSelect_hi_lo = _GEN_1;
  wire [63:0]       maskSplit_maskSelect_hi_lo_1;
  assign maskSplit_maskSelect_hi_lo_1 = _GEN_1;
  wire [63:0]       maskSplit_maskSelect_hi_lo_2;
  assign maskSplit_maskSelect_hi_lo_2 = _GEN_1;
  wire [63:0]       maskForDestination_hi_lo;
  assign maskForDestination_hi_lo = _GEN_1;
  wire [63:0]       _GEN_2 = {v0_7, v0_6};
  wire [63:0]       regroupV0_hi_hi;
  assign regroupV0_hi_hi = _GEN_2;
  wire [63:0]       regroupV0_hi_hi_5;
  assign regroupV0_hi_hi_5 = _GEN_2;
  wire [63:0]       regroupV0_hi_hi_10;
  assign regroupV0_hi_hi_10 = _GEN_2;
  wire [63:0]       slideAddressGen_slideMaskInput_hi_hi;
  assign slideAddressGen_slideMaskInput_hi_hi = _GEN_2;
  wire [63:0]       selectReadStageMask_hi_hi;
  assign selectReadStageMask_hi_hi = _GEN_2;
  wire [63:0]       maskSplit_maskSelect_hi_hi;
  assign maskSplit_maskSelect_hi_hi = _GEN_2;
  wire [63:0]       maskSplit_maskSelect_hi_hi_1;
  assign maskSplit_maskSelect_hi_hi_1 = _GEN_2;
  wire [63:0]       maskSplit_maskSelect_hi_hi_2;
  assign maskSplit_maskSelect_hi_hi_2 = _GEN_2;
  wire [63:0]       maskForDestination_hi_hi;
  assign maskForDestination_hi_hi = _GEN_2;
  wire [127:0]      regroupV0_hi = {regroupV0_hi_hi, regroupV0_hi_lo};
  wire [7:0]        regroupV0_lo_lo_lo = {regroupV0_lo[19:16], regroupV0_lo[3:0]};
  wire [7:0]        regroupV0_lo_lo_hi = {regroupV0_lo[51:48], regroupV0_lo[35:32]};
  wire [15:0]       regroupV0_lo_lo_1 = {regroupV0_lo_lo_hi, regroupV0_lo_lo_lo};
  wire [7:0]        regroupV0_lo_hi_lo = {regroupV0_lo[83:80], regroupV0_lo[67:64]};
  wire [7:0]        regroupV0_lo_hi_hi = {regroupV0_lo[115:112], regroupV0_lo[99:96]};
  wire [15:0]       regroupV0_lo_hi_1 = {regroupV0_lo_hi_hi, regroupV0_lo_hi_lo};
  wire [31:0]       regroupV0_lo_1 = {regroupV0_lo_hi_1, regroupV0_lo_lo_1};
  wire [7:0]        regroupV0_hi_lo_lo = {regroupV0_hi[19:16], regroupV0_hi[3:0]};
  wire [7:0]        regroupV0_hi_lo_hi = {regroupV0_hi[51:48], regroupV0_hi[35:32]};
  wire [15:0]       regroupV0_hi_lo_1 = {regroupV0_hi_lo_hi, regroupV0_hi_lo_lo};
  wire [7:0]        regroupV0_hi_hi_lo = {regroupV0_hi[83:80], regroupV0_hi[67:64]};
  wire [7:0]        regroupV0_hi_hi_hi = {regroupV0_hi[115:112], regroupV0_hi[99:96]};
  wire [15:0]       regroupV0_hi_hi_1 = {regroupV0_hi_hi_hi, regroupV0_hi_hi_lo};
  wire [31:0]       regroupV0_hi_1 = {regroupV0_hi_hi_1, regroupV0_hi_lo_1};
  wire [7:0]        regroupV0_lo_lo_lo_1 = {regroupV0_lo[23:20], regroupV0_lo[7:4]};
  wire [7:0]        regroupV0_lo_lo_hi_1 = {regroupV0_lo[55:52], regroupV0_lo[39:36]};
  wire [15:0]       regroupV0_lo_lo_2 = {regroupV0_lo_lo_hi_1, regroupV0_lo_lo_lo_1};
  wire [7:0]        regroupV0_lo_hi_lo_1 = {regroupV0_lo[87:84], regroupV0_lo[71:68]};
  wire [7:0]        regroupV0_lo_hi_hi_1 = {regroupV0_lo[119:116], regroupV0_lo[103:100]};
  wire [15:0]       regroupV0_lo_hi_2 = {regroupV0_lo_hi_hi_1, regroupV0_lo_hi_lo_1};
  wire [31:0]       regroupV0_lo_2 = {regroupV0_lo_hi_2, regroupV0_lo_lo_2};
  wire [7:0]        regroupV0_hi_lo_lo_1 = {regroupV0_hi[23:20], regroupV0_hi[7:4]};
  wire [7:0]        regroupV0_hi_lo_hi_1 = {regroupV0_hi[55:52], regroupV0_hi[39:36]};
  wire [15:0]       regroupV0_hi_lo_2 = {regroupV0_hi_lo_hi_1, regroupV0_hi_lo_lo_1};
  wire [7:0]        regroupV0_hi_hi_lo_1 = {regroupV0_hi[87:84], regroupV0_hi[71:68]};
  wire [7:0]        regroupV0_hi_hi_hi_1 = {regroupV0_hi[119:116], regroupV0_hi[103:100]};
  wire [15:0]       regroupV0_hi_hi_2 = {regroupV0_hi_hi_hi_1, regroupV0_hi_hi_lo_1};
  wire [31:0]       regroupV0_hi_2 = {regroupV0_hi_hi_2, regroupV0_hi_lo_2};
  wire [7:0]        regroupV0_lo_lo_lo_2 = {regroupV0_lo[27:24], regroupV0_lo[11:8]};
  wire [7:0]        regroupV0_lo_lo_hi_2 = {regroupV0_lo[59:56], regroupV0_lo[43:40]};
  wire [15:0]       regroupV0_lo_lo_3 = {regroupV0_lo_lo_hi_2, regroupV0_lo_lo_lo_2};
  wire [7:0]        regroupV0_lo_hi_lo_2 = {regroupV0_lo[91:88], regroupV0_lo[75:72]};
  wire [7:0]        regroupV0_lo_hi_hi_2 = {regroupV0_lo[123:120], regroupV0_lo[107:104]};
  wire [15:0]       regroupV0_lo_hi_3 = {regroupV0_lo_hi_hi_2, regroupV0_lo_hi_lo_2};
  wire [31:0]       regroupV0_lo_3 = {regroupV0_lo_hi_3, regroupV0_lo_lo_3};
  wire [7:0]        regroupV0_hi_lo_lo_2 = {regroupV0_hi[27:24], regroupV0_hi[11:8]};
  wire [7:0]        regroupV0_hi_lo_hi_2 = {regroupV0_hi[59:56], regroupV0_hi[43:40]};
  wire [15:0]       regroupV0_hi_lo_3 = {regroupV0_hi_lo_hi_2, regroupV0_hi_lo_lo_2};
  wire [7:0]        regroupV0_hi_hi_lo_2 = {regroupV0_hi[91:88], regroupV0_hi[75:72]};
  wire [7:0]        regroupV0_hi_hi_hi_2 = {regroupV0_hi[123:120], regroupV0_hi[107:104]};
  wire [15:0]       regroupV0_hi_hi_3 = {regroupV0_hi_hi_hi_2, regroupV0_hi_hi_lo_2};
  wire [31:0]       regroupV0_hi_3 = {regroupV0_hi_hi_3, regroupV0_hi_lo_3};
  wire [7:0]        regroupV0_lo_lo_lo_3 = {regroupV0_lo[31:28], regroupV0_lo[15:12]};
  wire [7:0]        regroupV0_lo_lo_hi_3 = {regroupV0_lo[63:60], regroupV0_lo[47:44]};
  wire [15:0]       regroupV0_lo_lo_4 = {regroupV0_lo_lo_hi_3, regroupV0_lo_lo_lo_3};
  wire [7:0]        regroupV0_lo_hi_lo_3 = {regroupV0_lo[95:92], regroupV0_lo[79:76]};
  wire [7:0]        regroupV0_lo_hi_hi_3 = {regroupV0_lo[127:124], regroupV0_lo[111:108]};
  wire [15:0]       regroupV0_lo_hi_4 = {regroupV0_lo_hi_hi_3, regroupV0_lo_hi_lo_3};
  wire [31:0]       regroupV0_lo_4 = {regroupV0_lo_hi_4, regroupV0_lo_lo_4};
  wire [7:0]        regroupV0_hi_lo_lo_3 = {regroupV0_hi[31:28], regroupV0_hi[15:12]};
  wire [7:0]        regroupV0_hi_lo_hi_3 = {regroupV0_hi[63:60], regroupV0_hi[47:44]};
  wire [15:0]       regroupV0_hi_lo_4 = {regroupV0_hi_lo_hi_3, regroupV0_hi_lo_lo_3};
  wire [7:0]        regroupV0_hi_hi_lo_3 = {regroupV0_hi[95:92], regroupV0_hi[79:76]};
  wire [7:0]        regroupV0_hi_hi_hi_3 = {regroupV0_hi[127:124], regroupV0_hi[111:108]};
  wire [15:0]       regroupV0_hi_hi_4 = {regroupV0_hi_hi_hi_3, regroupV0_hi_hi_lo_3};
  wire [31:0]       regroupV0_hi_4 = {regroupV0_hi_hi_4, regroupV0_hi_lo_4};
  wire [127:0]      regroupV0_lo_5 = {regroupV0_hi_2, regroupV0_lo_2, regroupV0_hi_1, regroupV0_lo_1};
  wire [127:0]      regroupV0_hi_5 = {regroupV0_hi_4, regroupV0_lo_4, regroupV0_hi_3, regroupV0_lo_3};
  wire [255:0]      regroupV0_0 = {regroupV0_hi_5, regroupV0_lo_5};
  wire [127:0]      regroupV0_lo_6 = {regroupV0_lo_hi_5, regroupV0_lo_lo_5};
  wire [127:0]      regroupV0_hi_6 = {regroupV0_hi_hi_5, regroupV0_hi_lo_5};
  wire [3:0]        regroupV0_lo_lo_lo_lo = {regroupV0_lo_6[9:8], regroupV0_lo_6[1:0]};
  wire [3:0]        regroupV0_lo_lo_lo_hi = {regroupV0_lo_6[25:24], regroupV0_lo_6[17:16]};
  wire [7:0]        regroupV0_lo_lo_lo_4 = {regroupV0_lo_lo_lo_hi, regroupV0_lo_lo_lo_lo};
  wire [3:0]        regroupV0_lo_lo_hi_lo = {regroupV0_lo_6[41:40], regroupV0_lo_6[33:32]};
  wire [3:0]        regroupV0_lo_lo_hi_hi = {regroupV0_lo_6[57:56], regroupV0_lo_6[49:48]};
  wire [7:0]        regroupV0_lo_lo_hi_4 = {regroupV0_lo_lo_hi_hi, regroupV0_lo_lo_hi_lo};
  wire [15:0]       regroupV0_lo_lo_6 = {regroupV0_lo_lo_hi_4, regroupV0_lo_lo_lo_4};
  wire [3:0]        regroupV0_lo_hi_lo_lo = {regroupV0_lo_6[73:72], regroupV0_lo_6[65:64]};
  wire [3:0]        regroupV0_lo_hi_lo_hi = {regroupV0_lo_6[89:88], regroupV0_lo_6[81:80]};
  wire [7:0]        regroupV0_lo_hi_lo_4 = {regroupV0_lo_hi_lo_hi, regroupV0_lo_hi_lo_lo};
  wire [3:0]        regroupV0_lo_hi_hi_lo = {regroupV0_lo_6[105:104], regroupV0_lo_6[97:96]};
  wire [3:0]        regroupV0_lo_hi_hi_hi = {regroupV0_lo_6[121:120], regroupV0_lo_6[113:112]};
  wire [7:0]        regroupV0_lo_hi_hi_4 = {regroupV0_lo_hi_hi_hi, regroupV0_lo_hi_hi_lo};
  wire [15:0]       regroupV0_lo_hi_6 = {regroupV0_lo_hi_hi_4, regroupV0_lo_hi_lo_4};
  wire [31:0]       regroupV0_lo_7 = {regroupV0_lo_hi_6, regroupV0_lo_lo_6};
  wire [3:0]        regroupV0_hi_lo_lo_lo = {regroupV0_hi_6[9:8], regroupV0_hi_6[1:0]};
  wire [3:0]        regroupV0_hi_lo_lo_hi = {regroupV0_hi_6[25:24], regroupV0_hi_6[17:16]};
  wire [7:0]        regroupV0_hi_lo_lo_4 = {regroupV0_hi_lo_lo_hi, regroupV0_hi_lo_lo_lo};
  wire [3:0]        regroupV0_hi_lo_hi_lo = {regroupV0_hi_6[41:40], regroupV0_hi_6[33:32]};
  wire [3:0]        regroupV0_hi_lo_hi_hi = {regroupV0_hi_6[57:56], regroupV0_hi_6[49:48]};
  wire [7:0]        regroupV0_hi_lo_hi_4 = {regroupV0_hi_lo_hi_hi, regroupV0_hi_lo_hi_lo};
  wire [15:0]       regroupV0_hi_lo_6 = {regroupV0_hi_lo_hi_4, regroupV0_hi_lo_lo_4};
  wire [3:0]        regroupV0_hi_hi_lo_lo = {regroupV0_hi_6[73:72], regroupV0_hi_6[65:64]};
  wire [3:0]        regroupV0_hi_hi_lo_hi = {regroupV0_hi_6[89:88], regroupV0_hi_6[81:80]};
  wire [7:0]        regroupV0_hi_hi_lo_4 = {regroupV0_hi_hi_lo_hi, regroupV0_hi_hi_lo_lo};
  wire [3:0]        regroupV0_hi_hi_hi_lo = {regroupV0_hi_6[105:104], regroupV0_hi_6[97:96]};
  wire [3:0]        regroupV0_hi_hi_hi_hi = {regroupV0_hi_6[121:120], regroupV0_hi_6[113:112]};
  wire [7:0]        regroupV0_hi_hi_hi_4 = {regroupV0_hi_hi_hi_hi, regroupV0_hi_hi_hi_lo};
  wire [15:0]       regroupV0_hi_hi_6 = {regroupV0_hi_hi_hi_4, regroupV0_hi_hi_lo_4};
  wire [31:0]       regroupV0_hi_7 = {regroupV0_hi_hi_6, regroupV0_hi_lo_6};
  wire [3:0]        regroupV0_lo_lo_lo_lo_1 = {regroupV0_lo_6[11:10], regroupV0_lo_6[3:2]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_1 = {regroupV0_lo_6[27:26], regroupV0_lo_6[19:18]};
  wire [7:0]        regroupV0_lo_lo_lo_5 = {regroupV0_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_1};
  wire [3:0]        regroupV0_lo_lo_hi_lo_1 = {regroupV0_lo_6[43:42], regroupV0_lo_6[35:34]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_1 = {regroupV0_lo_6[59:58], regroupV0_lo_6[51:50]};
  wire [7:0]        regroupV0_lo_lo_hi_5 = {regroupV0_lo_lo_hi_hi_1, regroupV0_lo_lo_hi_lo_1};
  wire [15:0]       regroupV0_lo_lo_7 = {regroupV0_lo_lo_hi_5, regroupV0_lo_lo_lo_5};
  wire [3:0]        regroupV0_lo_hi_lo_lo_1 = {regroupV0_lo_6[75:74], regroupV0_lo_6[67:66]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_1 = {regroupV0_lo_6[91:90], regroupV0_lo_6[83:82]};
  wire [7:0]        regroupV0_lo_hi_lo_5 = {regroupV0_lo_hi_lo_hi_1, regroupV0_lo_hi_lo_lo_1};
  wire [3:0]        regroupV0_lo_hi_hi_lo_1 = {regroupV0_lo_6[107:106], regroupV0_lo_6[99:98]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_1 = {regroupV0_lo_6[123:122], regroupV0_lo_6[115:114]};
  wire [7:0]        regroupV0_lo_hi_hi_5 = {regroupV0_lo_hi_hi_hi_1, regroupV0_lo_hi_hi_lo_1};
  wire [15:0]       regroupV0_lo_hi_7 = {regroupV0_lo_hi_hi_5, regroupV0_lo_hi_lo_5};
  wire [31:0]       regroupV0_lo_8 = {regroupV0_lo_hi_7, regroupV0_lo_lo_7};
  wire [3:0]        regroupV0_hi_lo_lo_lo_1 = {regroupV0_hi_6[11:10], regroupV0_hi_6[3:2]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_1 = {regroupV0_hi_6[27:26], regroupV0_hi_6[19:18]};
  wire [7:0]        regroupV0_hi_lo_lo_5 = {regroupV0_hi_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_1};
  wire [3:0]        regroupV0_hi_lo_hi_lo_1 = {regroupV0_hi_6[43:42], regroupV0_hi_6[35:34]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_1 = {regroupV0_hi_6[59:58], regroupV0_hi_6[51:50]};
  wire [7:0]        regroupV0_hi_lo_hi_5 = {regroupV0_hi_lo_hi_hi_1, regroupV0_hi_lo_hi_lo_1};
  wire [15:0]       regroupV0_hi_lo_7 = {regroupV0_hi_lo_hi_5, regroupV0_hi_lo_lo_5};
  wire [3:0]        regroupV0_hi_hi_lo_lo_1 = {regroupV0_hi_6[75:74], regroupV0_hi_6[67:66]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_1 = {regroupV0_hi_6[91:90], regroupV0_hi_6[83:82]};
  wire [7:0]        regroupV0_hi_hi_lo_5 = {regroupV0_hi_hi_lo_hi_1, regroupV0_hi_hi_lo_lo_1};
  wire [3:0]        regroupV0_hi_hi_hi_lo_1 = {regroupV0_hi_6[107:106], regroupV0_hi_6[99:98]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_1 = {regroupV0_hi_6[123:122], regroupV0_hi_6[115:114]};
  wire [7:0]        regroupV0_hi_hi_hi_5 = {regroupV0_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_lo_1};
  wire [15:0]       regroupV0_hi_hi_7 = {regroupV0_hi_hi_hi_5, regroupV0_hi_hi_lo_5};
  wire [31:0]       regroupV0_hi_8 = {regroupV0_hi_hi_7, regroupV0_hi_lo_7};
  wire [3:0]        regroupV0_lo_lo_lo_lo_2 = {regroupV0_lo_6[13:12], regroupV0_lo_6[5:4]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_2 = {regroupV0_lo_6[29:28], regroupV0_lo_6[21:20]};
  wire [7:0]        regroupV0_lo_lo_lo_6 = {regroupV0_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_2};
  wire [3:0]        regroupV0_lo_lo_hi_lo_2 = {regroupV0_lo_6[45:44], regroupV0_lo_6[37:36]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_2 = {regroupV0_lo_6[61:60], regroupV0_lo_6[53:52]};
  wire [7:0]        regroupV0_lo_lo_hi_6 = {regroupV0_lo_lo_hi_hi_2, regroupV0_lo_lo_hi_lo_2};
  wire [15:0]       regroupV0_lo_lo_8 = {regroupV0_lo_lo_hi_6, regroupV0_lo_lo_lo_6};
  wire [3:0]        regroupV0_lo_hi_lo_lo_2 = {regroupV0_lo_6[77:76], regroupV0_lo_6[69:68]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_2 = {regroupV0_lo_6[93:92], regroupV0_lo_6[85:84]};
  wire [7:0]        regroupV0_lo_hi_lo_6 = {regroupV0_lo_hi_lo_hi_2, regroupV0_lo_hi_lo_lo_2};
  wire [3:0]        regroupV0_lo_hi_hi_lo_2 = {regroupV0_lo_6[109:108], regroupV0_lo_6[101:100]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_2 = {regroupV0_lo_6[125:124], regroupV0_lo_6[117:116]};
  wire [7:0]        regroupV0_lo_hi_hi_6 = {regroupV0_lo_hi_hi_hi_2, regroupV0_lo_hi_hi_lo_2};
  wire [15:0]       regroupV0_lo_hi_8 = {regroupV0_lo_hi_hi_6, regroupV0_lo_hi_lo_6};
  wire [31:0]       regroupV0_lo_9 = {regroupV0_lo_hi_8, regroupV0_lo_lo_8};
  wire [3:0]        regroupV0_hi_lo_lo_lo_2 = {regroupV0_hi_6[13:12], regroupV0_hi_6[5:4]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_2 = {regroupV0_hi_6[29:28], regroupV0_hi_6[21:20]};
  wire [7:0]        regroupV0_hi_lo_lo_6 = {regroupV0_hi_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_2};
  wire [3:0]        regroupV0_hi_lo_hi_lo_2 = {regroupV0_hi_6[45:44], regroupV0_hi_6[37:36]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_2 = {regroupV0_hi_6[61:60], regroupV0_hi_6[53:52]};
  wire [7:0]        regroupV0_hi_lo_hi_6 = {regroupV0_hi_lo_hi_hi_2, regroupV0_hi_lo_hi_lo_2};
  wire [15:0]       regroupV0_hi_lo_8 = {regroupV0_hi_lo_hi_6, regroupV0_hi_lo_lo_6};
  wire [3:0]        regroupV0_hi_hi_lo_lo_2 = {regroupV0_hi_6[77:76], regroupV0_hi_6[69:68]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_2 = {regroupV0_hi_6[93:92], regroupV0_hi_6[85:84]};
  wire [7:0]        regroupV0_hi_hi_lo_6 = {regroupV0_hi_hi_lo_hi_2, regroupV0_hi_hi_lo_lo_2};
  wire [3:0]        regroupV0_hi_hi_hi_lo_2 = {regroupV0_hi_6[109:108], regroupV0_hi_6[101:100]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_2 = {regroupV0_hi_6[125:124], regroupV0_hi_6[117:116]};
  wire [7:0]        regroupV0_hi_hi_hi_6 = {regroupV0_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_lo_2};
  wire [15:0]       regroupV0_hi_hi_8 = {regroupV0_hi_hi_hi_6, regroupV0_hi_hi_lo_6};
  wire [31:0]       regroupV0_hi_9 = {regroupV0_hi_hi_8, regroupV0_hi_lo_8};
  wire [3:0]        regroupV0_lo_lo_lo_lo_3 = {regroupV0_lo_6[15:14], regroupV0_lo_6[7:6]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_3 = {regroupV0_lo_6[31:30], regroupV0_lo_6[23:22]};
  wire [7:0]        regroupV0_lo_lo_lo_7 = {regroupV0_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_3};
  wire [3:0]        regroupV0_lo_lo_hi_lo_3 = {regroupV0_lo_6[47:46], regroupV0_lo_6[39:38]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_3 = {regroupV0_lo_6[63:62], regroupV0_lo_6[55:54]};
  wire [7:0]        regroupV0_lo_lo_hi_7 = {regroupV0_lo_lo_hi_hi_3, regroupV0_lo_lo_hi_lo_3};
  wire [15:0]       regroupV0_lo_lo_9 = {regroupV0_lo_lo_hi_7, regroupV0_lo_lo_lo_7};
  wire [3:0]        regroupV0_lo_hi_lo_lo_3 = {regroupV0_lo_6[79:78], regroupV0_lo_6[71:70]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_3 = {regroupV0_lo_6[95:94], regroupV0_lo_6[87:86]};
  wire [7:0]        regroupV0_lo_hi_lo_7 = {regroupV0_lo_hi_lo_hi_3, regroupV0_lo_hi_lo_lo_3};
  wire [3:0]        regroupV0_lo_hi_hi_lo_3 = {regroupV0_lo_6[111:110], regroupV0_lo_6[103:102]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_3 = {regroupV0_lo_6[127:126], regroupV0_lo_6[119:118]};
  wire [7:0]        regroupV0_lo_hi_hi_7 = {regroupV0_lo_hi_hi_hi_3, regroupV0_lo_hi_hi_lo_3};
  wire [15:0]       regroupV0_lo_hi_9 = {regroupV0_lo_hi_hi_7, regroupV0_lo_hi_lo_7};
  wire [31:0]       regroupV0_lo_10 = {regroupV0_lo_hi_9, regroupV0_lo_lo_9};
  wire [3:0]        regroupV0_hi_lo_lo_lo_3 = {regroupV0_hi_6[15:14], regroupV0_hi_6[7:6]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_3 = {regroupV0_hi_6[31:30], regroupV0_hi_6[23:22]};
  wire [7:0]        regroupV0_hi_lo_lo_7 = {regroupV0_hi_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_3};
  wire [3:0]        regroupV0_hi_lo_hi_lo_3 = {regroupV0_hi_6[47:46], regroupV0_hi_6[39:38]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_3 = {regroupV0_hi_6[63:62], regroupV0_hi_6[55:54]};
  wire [7:0]        regroupV0_hi_lo_hi_7 = {regroupV0_hi_lo_hi_hi_3, regroupV0_hi_lo_hi_lo_3};
  wire [15:0]       regroupV0_hi_lo_9 = {regroupV0_hi_lo_hi_7, regroupV0_hi_lo_lo_7};
  wire [3:0]        regroupV0_hi_hi_lo_lo_3 = {regroupV0_hi_6[79:78], regroupV0_hi_6[71:70]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_3 = {regroupV0_hi_6[95:94], regroupV0_hi_6[87:86]};
  wire [7:0]        regroupV0_hi_hi_lo_7 = {regroupV0_hi_hi_lo_hi_3, regroupV0_hi_hi_lo_lo_3};
  wire [3:0]        regroupV0_hi_hi_hi_lo_3 = {regroupV0_hi_6[111:110], regroupV0_hi_6[103:102]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_3 = {regroupV0_hi_6[127:126], regroupV0_hi_6[119:118]};
  wire [7:0]        regroupV0_hi_hi_hi_7 = {regroupV0_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_lo_3};
  wire [15:0]       regroupV0_hi_hi_9 = {regroupV0_hi_hi_hi_7, regroupV0_hi_hi_lo_7};
  wire [31:0]       regroupV0_hi_10 = {regroupV0_hi_hi_9, regroupV0_hi_lo_9};
  wire [127:0]      regroupV0_lo_11 = {regroupV0_hi_8, regroupV0_lo_8, regroupV0_hi_7, regroupV0_lo_7};
  wire [127:0]      regroupV0_hi_11 = {regroupV0_hi_10, regroupV0_lo_10, regroupV0_hi_9, regroupV0_lo_9};
  wire [255:0]      regroupV0_1 = {regroupV0_hi_11, regroupV0_lo_11};
  wire [127:0]      regroupV0_lo_12 = {regroupV0_lo_hi_10, regroupV0_lo_lo_10};
  wire [127:0]      regroupV0_hi_12 = {regroupV0_hi_hi_10, regroupV0_hi_lo_10};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo = {regroupV0_lo_12[4], regroupV0_lo_12[0]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi = {regroupV0_lo_12[12], regroupV0_lo_12[8]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_4 = {regroupV0_lo_lo_lo_lo_hi, regroupV0_lo_lo_lo_lo_lo};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo = {regroupV0_lo_12[20], regroupV0_lo_12[16]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi = {regroupV0_lo_12[28], regroupV0_lo_12[24]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_4 = {regroupV0_lo_lo_lo_hi_hi, regroupV0_lo_lo_lo_hi_lo};
  wire [7:0]        regroupV0_lo_lo_lo_8 = {regroupV0_lo_lo_lo_hi_4, regroupV0_lo_lo_lo_lo_4};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo = {regroupV0_lo_12[36], regroupV0_lo_12[32]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi = {regroupV0_lo_12[44], regroupV0_lo_12[40]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_4 = {regroupV0_lo_lo_hi_lo_hi, regroupV0_lo_lo_hi_lo_lo};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo = {regroupV0_lo_12[52], regroupV0_lo_12[48]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi = {regroupV0_lo_12[60], regroupV0_lo_12[56]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_4 = {regroupV0_lo_lo_hi_hi_hi, regroupV0_lo_lo_hi_hi_lo};
  wire [7:0]        regroupV0_lo_lo_hi_8 = {regroupV0_lo_lo_hi_hi_4, regroupV0_lo_lo_hi_lo_4};
  wire [15:0]       regroupV0_lo_lo_11 = {regroupV0_lo_lo_hi_8, regroupV0_lo_lo_lo_8};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo = {regroupV0_lo_12[68], regroupV0_lo_12[64]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi = {regroupV0_lo_12[76], regroupV0_lo_12[72]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_4 = {regroupV0_lo_hi_lo_lo_hi, regroupV0_lo_hi_lo_lo_lo};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo = {regroupV0_lo_12[84], regroupV0_lo_12[80]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi = {regroupV0_lo_12[92], regroupV0_lo_12[88]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_4 = {regroupV0_lo_hi_lo_hi_hi, regroupV0_lo_hi_lo_hi_lo};
  wire [7:0]        regroupV0_lo_hi_lo_8 = {regroupV0_lo_hi_lo_hi_4, regroupV0_lo_hi_lo_lo_4};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo = {regroupV0_lo_12[100], regroupV0_lo_12[96]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi = {regroupV0_lo_12[108], regroupV0_lo_12[104]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_4 = {regroupV0_lo_hi_hi_lo_hi, regroupV0_lo_hi_hi_lo_lo};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo = {regroupV0_lo_12[116], regroupV0_lo_12[112]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi = {regroupV0_lo_12[124], regroupV0_lo_12[120]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_4 = {regroupV0_lo_hi_hi_hi_hi, regroupV0_lo_hi_hi_hi_lo};
  wire [7:0]        regroupV0_lo_hi_hi_8 = {regroupV0_lo_hi_hi_hi_4, regroupV0_lo_hi_hi_lo_4};
  wire [15:0]       regroupV0_lo_hi_11 = {regroupV0_lo_hi_hi_8, regroupV0_lo_hi_lo_8};
  wire [31:0]       regroupV0_lo_13 = {regroupV0_lo_hi_11, regroupV0_lo_lo_11};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo = {regroupV0_hi_12[4], regroupV0_hi_12[0]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi = {regroupV0_hi_12[12], regroupV0_hi_12[8]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_4 = {regroupV0_hi_lo_lo_lo_hi, regroupV0_hi_lo_lo_lo_lo};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo = {regroupV0_hi_12[20], regroupV0_hi_12[16]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi = {regroupV0_hi_12[28], regroupV0_hi_12[24]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_4 = {regroupV0_hi_lo_lo_hi_hi, regroupV0_hi_lo_lo_hi_lo};
  wire [7:0]        regroupV0_hi_lo_lo_8 = {regroupV0_hi_lo_lo_hi_4, regroupV0_hi_lo_lo_lo_4};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo = {regroupV0_hi_12[36], regroupV0_hi_12[32]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi = {regroupV0_hi_12[44], regroupV0_hi_12[40]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_4 = {regroupV0_hi_lo_hi_lo_hi, regroupV0_hi_lo_hi_lo_lo};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo = {regroupV0_hi_12[52], regroupV0_hi_12[48]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi = {regroupV0_hi_12[60], regroupV0_hi_12[56]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_4 = {regroupV0_hi_lo_hi_hi_hi, regroupV0_hi_lo_hi_hi_lo};
  wire [7:0]        regroupV0_hi_lo_hi_8 = {regroupV0_hi_lo_hi_hi_4, regroupV0_hi_lo_hi_lo_4};
  wire [15:0]       regroupV0_hi_lo_11 = {regroupV0_hi_lo_hi_8, regroupV0_hi_lo_lo_8};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo = {regroupV0_hi_12[68], regroupV0_hi_12[64]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi = {regroupV0_hi_12[76], regroupV0_hi_12[72]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_4 = {regroupV0_hi_hi_lo_lo_hi, regroupV0_hi_hi_lo_lo_lo};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo = {regroupV0_hi_12[84], regroupV0_hi_12[80]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi = {regroupV0_hi_12[92], regroupV0_hi_12[88]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_4 = {regroupV0_hi_hi_lo_hi_hi, regroupV0_hi_hi_lo_hi_lo};
  wire [7:0]        regroupV0_hi_hi_lo_8 = {regroupV0_hi_hi_lo_hi_4, regroupV0_hi_hi_lo_lo_4};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo = {regroupV0_hi_12[100], regroupV0_hi_12[96]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi = {regroupV0_hi_12[108], regroupV0_hi_12[104]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_4 = {regroupV0_hi_hi_hi_lo_hi, regroupV0_hi_hi_hi_lo_lo};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo = {regroupV0_hi_12[116], regroupV0_hi_12[112]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi = {regroupV0_hi_12[124], regroupV0_hi_12[120]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_4 = {regroupV0_hi_hi_hi_hi_hi, regroupV0_hi_hi_hi_hi_lo};
  wire [7:0]        regroupV0_hi_hi_hi_8 = {regroupV0_hi_hi_hi_hi_4, regroupV0_hi_hi_hi_lo_4};
  wire [15:0]       regroupV0_hi_hi_11 = {regroupV0_hi_hi_hi_8, regroupV0_hi_hi_lo_8};
  wire [31:0]       regroupV0_hi_13 = {regroupV0_hi_hi_11, regroupV0_hi_lo_11};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_1 = {regroupV0_lo_12[5], regroupV0_lo_12[1]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_1 = {regroupV0_lo_12[13], regroupV0_lo_12[9]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_5 = {regroupV0_lo_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_lo_1};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_1 = {regroupV0_lo_12[21], regroupV0_lo_12[17]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_1 = {regroupV0_lo_12[29], regroupV0_lo_12[25]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_5 = {regroupV0_lo_lo_lo_hi_hi_1, regroupV0_lo_lo_lo_hi_lo_1};
  wire [7:0]        regroupV0_lo_lo_lo_9 = {regroupV0_lo_lo_lo_hi_5, regroupV0_lo_lo_lo_lo_5};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_1 = {regroupV0_lo_12[37], regroupV0_lo_12[33]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_1 = {regroupV0_lo_12[45], regroupV0_lo_12[41]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_5 = {regroupV0_lo_lo_hi_lo_hi_1, regroupV0_lo_lo_hi_lo_lo_1};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_1 = {regroupV0_lo_12[53], regroupV0_lo_12[49]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_1 = {regroupV0_lo_12[61], regroupV0_lo_12[57]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_5 = {regroupV0_lo_lo_hi_hi_hi_1, regroupV0_lo_lo_hi_hi_lo_1};
  wire [7:0]        regroupV0_lo_lo_hi_9 = {regroupV0_lo_lo_hi_hi_5, regroupV0_lo_lo_hi_lo_5};
  wire [15:0]       regroupV0_lo_lo_12 = {regroupV0_lo_lo_hi_9, regroupV0_lo_lo_lo_9};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_1 = {regroupV0_lo_12[69], regroupV0_lo_12[65]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_1 = {regroupV0_lo_12[77], regroupV0_lo_12[73]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_5 = {regroupV0_lo_hi_lo_lo_hi_1, regroupV0_lo_hi_lo_lo_lo_1};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_1 = {regroupV0_lo_12[85], regroupV0_lo_12[81]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_1 = {regroupV0_lo_12[93], regroupV0_lo_12[89]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_5 = {regroupV0_lo_hi_lo_hi_hi_1, regroupV0_lo_hi_lo_hi_lo_1};
  wire [7:0]        regroupV0_lo_hi_lo_9 = {regroupV0_lo_hi_lo_hi_5, regroupV0_lo_hi_lo_lo_5};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_1 = {regroupV0_lo_12[101], regroupV0_lo_12[97]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_1 = {regroupV0_lo_12[109], regroupV0_lo_12[105]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_5 = {regroupV0_lo_hi_hi_lo_hi_1, regroupV0_lo_hi_hi_lo_lo_1};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_1 = {regroupV0_lo_12[117], regroupV0_lo_12[113]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_1 = {regroupV0_lo_12[125], regroupV0_lo_12[121]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_5 = {regroupV0_lo_hi_hi_hi_hi_1, regroupV0_lo_hi_hi_hi_lo_1};
  wire [7:0]        regroupV0_lo_hi_hi_9 = {regroupV0_lo_hi_hi_hi_5, regroupV0_lo_hi_hi_lo_5};
  wire [15:0]       regroupV0_lo_hi_12 = {regroupV0_lo_hi_hi_9, regroupV0_lo_hi_lo_9};
  wire [31:0]       regroupV0_lo_14 = {regroupV0_lo_hi_12, regroupV0_lo_lo_12};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_1 = {regroupV0_hi_12[5], regroupV0_hi_12[1]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_1 = {regroupV0_hi_12[13], regroupV0_hi_12[9]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_5 = {regroupV0_hi_lo_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_lo_1};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_1 = {regroupV0_hi_12[21], regroupV0_hi_12[17]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_1 = {regroupV0_hi_12[29], regroupV0_hi_12[25]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_5 = {regroupV0_hi_lo_lo_hi_hi_1, regroupV0_hi_lo_lo_hi_lo_1};
  wire [7:0]        regroupV0_hi_lo_lo_9 = {regroupV0_hi_lo_lo_hi_5, regroupV0_hi_lo_lo_lo_5};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_1 = {regroupV0_hi_12[37], regroupV0_hi_12[33]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_1 = {regroupV0_hi_12[45], regroupV0_hi_12[41]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_5 = {regroupV0_hi_lo_hi_lo_hi_1, regroupV0_hi_lo_hi_lo_lo_1};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_1 = {regroupV0_hi_12[53], regroupV0_hi_12[49]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_1 = {regroupV0_hi_12[61], regroupV0_hi_12[57]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_5 = {regroupV0_hi_lo_hi_hi_hi_1, regroupV0_hi_lo_hi_hi_lo_1};
  wire [7:0]        regroupV0_hi_lo_hi_9 = {regroupV0_hi_lo_hi_hi_5, regroupV0_hi_lo_hi_lo_5};
  wire [15:0]       regroupV0_hi_lo_12 = {regroupV0_hi_lo_hi_9, regroupV0_hi_lo_lo_9};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_1 = {regroupV0_hi_12[69], regroupV0_hi_12[65]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_1 = {regroupV0_hi_12[77], regroupV0_hi_12[73]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_5 = {regroupV0_hi_hi_lo_lo_hi_1, regroupV0_hi_hi_lo_lo_lo_1};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_1 = {regroupV0_hi_12[85], regroupV0_hi_12[81]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_1 = {regroupV0_hi_12[93], regroupV0_hi_12[89]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_5 = {regroupV0_hi_hi_lo_hi_hi_1, regroupV0_hi_hi_lo_hi_lo_1};
  wire [7:0]        regroupV0_hi_hi_lo_9 = {regroupV0_hi_hi_lo_hi_5, regroupV0_hi_hi_lo_lo_5};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_1 = {regroupV0_hi_12[101], regroupV0_hi_12[97]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_1 = {regroupV0_hi_12[109], regroupV0_hi_12[105]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_5 = {regroupV0_hi_hi_hi_lo_hi_1, regroupV0_hi_hi_hi_lo_lo_1};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_1 = {regroupV0_hi_12[117], regroupV0_hi_12[113]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_1 = {regroupV0_hi_12[125], regroupV0_hi_12[121]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_5 = {regroupV0_hi_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_hi_lo_1};
  wire [7:0]        regroupV0_hi_hi_hi_9 = {regroupV0_hi_hi_hi_hi_5, regroupV0_hi_hi_hi_lo_5};
  wire [15:0]       regroupV0_hi_hi_12 = {regroupV0_hi_hi_hi_9, regroupV0_hi_hi_lo_9};
  wire [31:0]       regroupV0_hi_14 = {regroupV0_hi_hi_12, regroupV0_hi_lo_12};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_2 = {regroupV0_lo_12[6], regroupV0_lo_12[2]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_2 = {regroupV0_lo_12[14], regroupV0_lo_12[10]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_6 = {regroupV0_lo_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_lo_2};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_2 = {regroupV0_lo_12[22], regroupV0_lo_12[18]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_2 = {regroupV0_lo_12[30], regroupV0_lo_12[26]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_6 = {regroupV0_lo_lo_lo_hi_hi_2, regroupV0_lo_lo_lo_hi_lo_2};
  wire [7:0]        regroupV0_lo_lo_lo_10 = {regroupV0_lo_lo_lo_hi_6, regroupV0_lo_lo_lo_lo_6};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_2 = {regroupV0_lo_12[38], regroupV0_lo_12[34]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_2 = {regroupV0_lo_12[46], regroupV0_lo_12[42]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_6 = {regroupV0_lo_lo_hi_lo_hi_2, regroupV0_lo_lo_hi_lo_lo_2};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_2 = {regroupV0_lo_12[54], regroupV0_lo_12[50]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_2 = {regroupV0_lo_12[62], regroupV0_lo_12[58]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_6 = {regroupV0_lo_lo_hi_hi_hi_2, regroupV0_lo_lo_hi_hi_lo_2};
  wire [7:0]        regroupV0_lo_lo_hi_10 = {regroupV0_lo_lo_hi_hi_6, regroupV0_lo_lo_hi_lo_6};
  wire [15:0]       regroupV0_lo_lo_13 = {regroupV0_lo_lo_hi_10, regroupV0_lo_lo_lo_10};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_2 = {regroupV0_lo_12[70], regroupV0_lo_12[66]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_2 = {regroupV0_lo_12[78], regroupV0_lo_12[74]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_6 = {regroupV0_lo_hi_lo_lo_hi_2, regroupV0_lo_hi_lo_lo_lo_2};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_2 = {regroupV0_lo_12[86], regroupV0_lo_12[82]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_2 = {regroupV0_lo_12[94], regroupV0_lo_12[90]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_6 = {regroupV0_lo_hi_lo_hi_hi_2, regroupV0_lo_hi_lo_hi_lo_2};
  wire [7:0]        regroupV0_lo_hi_lo_10 = {regroupV0_lo_hi_lo_hi_6, regroupV0_lo_hi_lo_lo_6};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_2 = {regroupV0_lo_12[102], regroupV0_lo_12[98]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_2 = {regroupV0_lo_12[110], regroupV0_lo_12[106]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_6 = {regroupV0_lo_hi_hi_lo_hi_2, regroupV0_lo_hi_hi_lo_lo_2};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_2 = {regroupV0_lo_12[118], regroupV0_lo_12[114]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_2 = {regroupV0_lo_12[126], regroupV0_lo_12[122]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_6 = {regroupV0_lo_hi_hi_hi_hi_2, regroupV0_lo_hi_hi_hi_lo_2};
  wire [7:0]        regroupV0_lo_hi_hi_10 = {regroupV0_lo_hi_hi_hi_6, regroupV0_lo_hi_hi_lo_6};
  wire [15:0]       regroupV0_lo_hi_13 = {regroupV0_lo_hi_hi_10, regroupV0_lo_hi_lo_10};
  wire [31:0]       regroupV0_lo_15 = {regroupV0_lo_hi_13, regroupV0_lo_lo_13};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_2 = {regroupV0_hi_12[6], regroupV0_hi_12[2]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_2 = {regroupV0_hi_12[14], regroupV0_hi_12[10]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_6 = {regroupV0_hi_lo_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_lo_2};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_2 = {regroupV0_hi_12[22], regroupV0_hi_12[18]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_2 = {regroupV0_hi_12[30], regroupV0_hi_12[26]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_6 = {regroupV0_hi_lo_lo_hi_hi_2, regroupV0_hi_lo_lo_hi_lo_2};
  wire [7:0]        regroupV0_hi_lo_lo_10 = {regroupV0_hi_lo_lo_hi_6, regroupV0_hi_lo_lo_lo_6};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_2 = {regroupV0_hi_12[38], regroupV0_hi_12[34]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_2 = {regroupV0_hi_12[46], regroupV0_hi_12[42]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_6 = {regroupV0_hi_lo_hi_lo_hi_2, regroupV0_hi_lo_hi_lo_lo_2};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_2 = {regroupV0_hi_12[54], regroupV0_hi_12[50]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_2 = {regroupV0_hi_12[62], regroupV0_hi_12[58]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_6 = {regroupV0_hi_lo_hi_hi_hi_2, regroupV0_hi_lo_hi_hi_lo_2};
  wire [7:0]        regroupV0_hi_lo_hi_10 = {regroupV0_hi_lo_hi_hi_6, regroupV0_hi_lo_hi_lo_6};
  wire [15:0]       regroupV0_hi_lo_13 = {regroupV0_hi_lo_hi_10, regroupV0_hi_lo_lo_10};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_2 = {regroupV0_hi_12[70], regroupV0_hi_12[66]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_2 = {regroupV0_hi_12[78], regroupV0_hi_12[74]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_6 = {regroupV0_hi_hi_lo_lo_hi_2, regroupV0_hi_hi_lo_lo_lo_2};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_2 = {regroupV0_hi_12[86], regroupV0_hi_12[82]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_2 = {regroupV0_hi_12[94], regroupV0_hi_12[90]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_6 = {regroupV0_hi_hi_lo_hi_hi_2, regroupV0_hi_hi_lo_hi_lo_2};
  wire [7:0]        regroupV0_hi_hi_lo_10 = {regroupV0_hi_hi_lo_hi_6, regroupV0_hi_hi_lo_lo_6};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_2 = {regroupV0_hi_12[102], regroupV0_hi_12[98]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_2 = {regroupV0_hi_12[110], regroupV0_hi_12[106]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_6 = {regroupV0_hi_hi_hi_lo_hi_2, regroupV0_hi_hi_hi_lo_lo_2};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_2 = {regroupV0_hi_12[118], regroupV0_hi_12[114]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_2 = {regroupV0_hi_12[126], regroupV0_hi_12[122]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_6 = {regroupV0_hi_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_hi_lo_2};
  wire [7:0]        regroupV0_hi_hi_hi_10 = {regroupV0_hi_hi_hi_hi_6, regroupV0_hi_hi_hi_lo_6};
  wire [15:0]       regroupV0_hi_hi_13 = {regroupV0_hi_hi_hi_10, regroupV0_hi_hi_lo_10};
  wire [31:0]       regroupV0_hi_15 = {regroupV0_hi_hi_13, regroupV0_hi_lo_13};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_3 = {regroupV0_lo_12[7], regroupV0_lo_12[3]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_3 = {regroupV0_lo_12[15], regroupV0_lo_12[11]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_7 = {regroupV0_lo_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_lo_3};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_3 = {regroupV0_lo_12[23], regroupV0_lo_12[19]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_3 = {regroupV0_lo_12[31], regroupV0_lo_12[27]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_7 = {regroupV0_lo_lo_lo_hi_hi_3, regroupV0_lo_lo_lo_hi_lo_3};
  wire [7:0]        regroupV0_lo_lo_lo_11 = {regroupV0_lo_lo_lo_hi_7, regroupV0_lo_lo_lo_lo_7};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_3 = {regroupV0_lo_12[39], regroupV0_lo_12[35]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_3 = {regroupV0_lo_12[47], regroupV0_lo_12[43]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_7 = {regroupV0_lo_lo_hi_lo_hi_3, regroupV0_lo_lo_hi_lo_lo_3};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_3 = {regroupV0_lo_12[55], regroupV0_lo_12[51]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_3 = {regroupV0_lo_12[63], regroupV0_lo_12[59]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_7 = {regroupV0_lo_lo_hi_hi_hi_3, regroupV0_lo_lo_hi_hi_lo_3};
  wire [7:0]        regroupV0_lo_lo_hi_11 = {regroupV0_lo_lo_hi_hi_7, regroupV0_lo_lo_hi_lo_7};
  wire [15:0]       regroupV0_lo_lo_14 = {regroupV0_lo_lo_hi_11, regroupV0_lo_lo_lo_11};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_3 = {regroupV0_lo_12[71], regroupV0_lo_12[67]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_3 = {regroupV0_lo_12[79], regroupV0_lo_12[75]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_7 = {regroupV0_lo_hi_lo_lo_hi_3, regroupV0_lo_hi_lo_lo_lo_3};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_3 = {regroupV0_lo_12[87], regroupV0_lo_12[83]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_3 = {regroupV0_lo_12[95], regroupV0_lo_12[91]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_7 = {regroupV0_lo_hi_lo_hi_hi_3, regroupV0_lo_hi_lo_hi_lo_3};
  wire [7:0]        regroupV0_lo_hi_lo_11 = {regroupV0_lo_hi_lo_hi_7, regroupV0_lo_hi_lo_lo_7};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_3 = {regroupV0_lo_12[103], regroupV0_lo_12[99]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_3 = {regroupV0_lo_12[111], regroupV0_lo_12[107]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_7 = {regroupV0_lo_hi_hi_lo_hi_3, regroupV0_lo_hi_hi_lo_lo_3};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_3 = {regroupV0_lo_12[119], regroupV0_lo_12[115]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_3 = {regroupV0_lo_12[127], regroupV0_lo_12[123]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_7 = {regroupV0_lo_hi_hi_hi_hi_3, regroupV0_lo_hi_hi_hi_lo_3};
  wire [7:0]        regroupV0_lo_hi_hi_11 = {regroupV0_lo_hi_hi_hi_7, regroupV0_lo_hi_hi_lo_7};
  wire [15:0]       regroupV0_lo_hi_14 = {regroupV0_lo_hi_hi_11, regroupV0_lo_hi_lo_11};
  wire [31:0]       regroupV0_lo_16 = {regroupV0_lo_hi_14, regroupV0_lo_lo_14};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_3 = {regroupV0_hi_12[7], regroupV0_hi_12[3]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_3 = {regroupV0_hi_12[15], regroupV0_hi_12[11]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_7 = {regroupV0_hi_lo_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_lo_3};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_3 = {regroupV0_hi_12[23], regroupV0_hi_12[19]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_3 = {regroupV0_hi_12[31], regroupV0_hi_12[27]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_7 = {regroupV0_hi_lo_lo_hi_hi_3, regroupV0_hi_lo_lo_hi_lo_3};
  wire [7:0]        regroupV0_hi_lo_lo_11 = {regroupV0_hi_lo_lo_hi_7, regroupV0_hi_lo_lo_lo_7};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_3 = {regroupV0_hi_12[39], regroupV0_hi_12[35]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_3 = {regroupV0_hi_12[47], regroupV0_hi_12[43]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_7 = {regroupV0_hi_lo_hi_lo_hi_3, regroupV0_hi_lo_hi_lo_lo_3};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_3 = {regroupV0_hi_12[55], regroupV0_hi_12[51]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_3 = {regroupV0_hi_12[63], regroupV0_hi_12[59]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_7 = {regroupV0_hi_lo_hi_hi_hi_3, regroupV0_hi_lo_hi_hi_lo_3};
  wire [7:0]        regroupV0_hi_lo_hi_11 = {regroupV0_hi_lo_hi_hi_7, regroupV0_hi_lo_hi_lo_7};
  wire [15:0]       regroupV0_hi_lo_14 = {regroupV0_hi_lo_hi_11, regroupV0_hi_lo_lo_11};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_3 = {regroupV0_hi_12[71], regroupV0_hi_12[67]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_3 = {regroupV0_hi_12[79], regroupV0_hi_12[75]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_7 = {regroupV0_hi_hi_lo_lo_hi_3, regroupV0_hi_hi_lo_lo_lo_3};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_3 = {regroupV0_hi_12[87], regroupV0_hi_12[83]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_3 = {regroupV0_hi_12[95], regroupV0_hi_12[91]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_7 = {regroupV0_hi_hi_lo_hi_hi_3, regroupV0_hi_hi_lo_hi_lo_3};
  wire [7:0]        regroupV0_hi_hi_lo_11 = {regroupV0_hi_hi_lo_hi_7, regroupV0_hi_hi_lo_lo_7};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_3 = {regroupV0_hi_12[103], regroupV0_hi_12[99]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_3 = {regroupV0_hi_12[111], regroupV0_hi_12[107]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_7 = {regroupV0_hi_hi_hi_lo_hi_3, regroupV0_hi_hi_hi_lo_lo_3};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_3 = {regroupV0_hi_12[119], regroupV0_hi_12[115]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_3 = {regroupV0_hi_12[127], regroupV0_hi_12[123]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_7 = {regroupV0_hi_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_hi_lo_3};
  wire [7:0]        regroupV0_hi_hi_hi_11 = {regroupV0_hi_hi_hi_hi_7, regroupV0_hi_hi_hi_lo_7};
  wire [15:0]       regroupV0_hi_hi_14 = {regroupV0_hi_hi_hi_11, regroupV0_hi_hi_lo_11};
  wire [31:0]       regroupV0_hi_16 = {regroupV0_hi_hi_14, regroupV0_hi_lo_14};
  wire [127:0]      regroupV0_lo_17 = {regroupV0_hi_14, regroupV0_lo_14, regroupV0_hi_13, regroupV0_lo_13};
  wire [127:0]      regroupV0_hi_17 = {regroupV0_hi_16, regroupV0_lo_16, regroupV0_hi_15, regroupV0_lo_15};
  wire [255:0]      regroupV0_2 = {regroupV0_hi_17, regroupV0_lo_17};
  wire [3:0]        _v0SelectBySew_T = 4'h1 << laneMaskSewSelect_0;
  wire [63:0]       v0SelectBySew = (_v0SelectBySew_T[0] ? regroupV0_0[63:0] : 64'h0) | (_v0SelectBySew_T[1] ? regroupV0_1[63:0] : 64'h0) | (_v0SelectBySew_T[2] ? regroupV0_2[63:0] : 64'h0);
  wire [3:0]        _v0SelectBySew_T_9 = 4'h1 << laneMaskSewSelect_1;
  wire [63:0]       v0SelectBySew_1 = (_v0SelectBySew_T_9[0] ? regroupV0_0[127:64] : 64'h0) | (_v0SelectBySew_T_9[1] ? regroupV0_1[127:64] : 64'h0) | (_v0SelectBySew_T_9[2] ? regroupV0_2[127:64] : 64'h0);
  wire [3:0]        _v0SelectBySew_T_18 = 4'h1 << laneMaskSewSelect_2;
  wire [63:0]       v0SelectBySew_2 = (_v0SelectBySew_T_18[0] ? regroupV0_0[191:128] : 64'h0) | (_v0SelectBySew_T_18[1] ? regroupV0_1[191:128] : 64'h0) | (_v0SelectBySew_T_18[2] ? regroupV0_2[191:128] : 64'h0);
  wire [3:0]        _v0SelectBySew_T_27 = 4'h1 << laneMaskSewSelect_3;
  wire [63:0]       v0SelectBySew_3 = (_v0SelectBySew_T_27[0] ? regroupV0_0[255:192] : 64'h0) | (_v0SelectBySew_T_27[1] ? regroupV0_1[255:192] : 64'h0) | (_v0SelectBySew_T_27[2] ? regroupV0_2[255:192] : 64'h0);
  wire [3:0]        intLMULInput = 4'h1 << instReq_bits_vlmul[1:0];
  wire [10:0]       _dataPosition_T_1 = {3'h0, instReq_bits_readFromScala[7:0]} << instReq_bits_sew;
  wire [7:0]        dataPosition = _dataPosition_T_1[7:0];
  wire [3:0]        _sewOHInput_T = 4'h1 << instReq_bits_sew;
  wire [2:0]        sewOHInput = _sewOHInput_T[2:0];
  wire [1:0]        dataOffset = {dataPosition[1] & (|(sewOHInput[1:0])), dataPosition[0] & sewOHInput[0]};
  wire [1:0]        accessLane = dataPosition[3:2];
  wire [3:0]        dataGroup = dataPosition[7:4];
  wire              offset = dataGroup[0];
  wire [2:0]        accessRegGrowth = dataGroup[3:1];
  wire [2:0]        reallyGrowth = accessRegGrowth;
  wire [2:0]        decimalProportion = {offset, accessLane};
  wire [2:0]        decimal = decimalProportion;
  wire              notNeedRead = |{instReq_bits_vlmul[2] & decimal >= intLMULInput[3:1] | ~(instReq_bits_vlmul[2]) & {1'h0, accessRegGrowth} >= intLMULInput, instReq_bits_readFromScala[31:8]};
  reg  [1:0]        gatherReadState;
  wire              gatherSRead = gatherReadState == 2'h1;
  wire              gatherWaiteRead = gatherReadState == 2'h2;
  assign gatherResponse = &gatherReadState;
  wire              gatherData_valid_0 = gatherResponse;
  reg  [1:0]        gatherDatOffset;
  reg  [1:0]        gatherLane;
  reg               gatherOffset;
  reg  [2:0]        gatherGrowth;
  reg  [2:0]        instReg_instructionIndex;
  wire [2:0]        exeResp_0_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        exeResp_1_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        exeResp_2_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        exeResp_3_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        readChannel_0_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        readChannel_1_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        readChannel_2_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        readChannel_3_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        writeRequest_0_index = instReg_instructionIndex;
  wire [2:0]        writeRequest_1_index = instReg_instructionIndex;
  wire [2:0]        writeRequest_2_index = instReg_instructionIndex;
  wire [2:0]        writeRequest_3_index = instReg_instructionIndex;
  wire [2:0]        writeQueue_0_enq_bits_index = instReg_instructionIndex;
  wire [2:0]        writeQueue_1_enq_bits_index = instReg_instructionIndex;
  wire [2:0]        writeQueue_2_enq_bits_index = instReg_instructionIndex;
  wire [2:0]        writeQueue_3_enq_bits_index = instReg_instructionIndex;
  reg               instReg_decodeResult_specialSlot;
  reg  [4:0]        instReg_decodeResult_topUop;
  reg               instReg_decodeResult_popCount;
  reg               instReg_decodeResult_ffo;
  reg               instReg_decodeResult_average;
  reg               instReg_decodeResult_reverse;
  reg               instReg_decodeResult_dontNeedExecuteInLane;
  reg               instReg_decodeResult_scheduler;
  reg               instReg_decodeResult_sReadVD;
  reg               instReg_decodeResult_vtype;
  reg               instReg_decodeResult_sWrite;
  reg               instReg_decodeResult_crossRead;
  reg               instReg_decodeResult_crossWrite;
  reg               instReg_decodeResult_maskUnit;
  reg               instReg_decodeResult_special;
  reg               instReg_decodeResult_saturate;
  reg               instReg_decodeResult_vwmacc;
  reg               instReg_decodeResult_readOnly;
  reg               instReg_decodeResult_maskSource;
  reg               instReg_decodeResult_maskDestination;
  reg               instReg_decodeResult_maskLogic;
  reg  [3:0]        instReg_decodeResult_uop;
  reg               instReg_decodeResult_iota;
  reg               instReg_decodeResult_mv;
  reg               instReg_decodeResult_extend;
  reg               instReg_decodeResult_unOrderWrite;
  reg               instReg_decodeResult_compress;
  reg               instReg_decodeResult_gather16;
  reg               instReg_decodeResult_gather;
  reg               instReg_decodeResult_slid;
  reg               instReg_decodeResult_targetRd;
  reg               instReg_decodeResult_widenReduce;
  reg               instReg_decodeResult_red;
  reg               instReg_decodeResult_nr;
  reg               instReg_decodeResult_itype;
  reg               instReg_decodeResult_unsigned1;
  reg               instReg_decodeResult_unsigned0;
  reg               instReg_decodeResult_other;
  reg               instReg_decodeResult_multiCycle;
  reg               instReg_decodeResult_divider;
  reg               instReg_decodeResult_multiplier;
  reg               instReg_decodeResult_shift;
  reg               instReg_decodeResult_adder;
  reg               instReg_decodeResult_logic;
  reg  [31:0]       instReg_readFromScala;
  reg  [1:0]        instReg_sew;
  reg  [2:0]        instReg_vlmul;
  reg               instReg_maskType;
  reg  [2:0]        instReg_vxrm;
  reg  [4:0]        instReg_vs2;
  reg  [4:0]        instReg_vs1;
  reg  [4:0]        instReg_vd;
  wire [4:0]        writeRequest_0_writeData_vd = instReg_vd;
  wire [4:0]        writeRequest_1_writeData_vd = instReg_vd;
  wire [4:0]        writeRequest_2_writeData_vd = instReg_vd;
  wire [4:0]        writeRequest_3_writeData_vd = instReg_vd;
  reg  [8:0]        instReg_vl;
  wire [8:0]        reduceLastDataNeed_byteForVl = instReg_vl;
  wire              enqMvRD = instReq_bits_decodeResult_topUop == 5'hB;
  reg               instVlValid;
  wire              gatherRequestFire = gatherReadState == 2'h0 & gatherRead & ~instVlValid;
  wire              viotaReq = instReq_bits_decodeResult_topUop == 5'h8;
  reg               readVS1Reg_dataValid;
  reg               readVS1Reg_requestSend;
  reg               readVS1Reg_sendToExecution;
  reg  [31:0]       readVS1Reg_data;
  reg  [3:0]        readVS1Reg_readIndex;
  wire [3:0]        _sew1H_T = 4'h1 << instReg_sew;
  wire [2:0]        sew1H = _sew1H_T[2:0];
  wire [3:0]        unitType = 4'h1 << instReg_decodeResult_topUop[4:3];
  wire [3:0]        subType = 4'h1 << instReg_decodeResult_topUop[2:1];
  wire              readType = unitType[0];
  wire              gather16 = instReg_decodeResult_topUop == 5'h5;
  wire              maskDestinationType = instReg_decodeResult_topUop == 5'h18;
  wire              compress = instReg_decodeResult_topUop[4:1] == 4'h4;
  wire              viota = instReg_decodeResult_topUop == 5'h8;
  wire              mv = instReg_decodeResult_topUop[4:1] == 4'h5;
  wire              mvRd = instReg_decodeResult_topUop == 5'hB;
  wire              mvVd = instReg_decodeResult_topUop == 5'hA;
  wire              orderReduce = {instReg_decodeResult_topUop[4:2], instReg_decodeResult_topUop[0]} == 4'hB;
  wire              ffo = instReg_decodeResult_topUop[4:1] == 4'h7;
  wire              extendType = unitType[3] & (subType[2] | subType[1]);
  wire              readValid = readType & instVlValid;
  wire              noSource = mv | viota;
  wire              allGroupExecute = maskDestinationType | unitType[2] | compress | ffo;
  wire              useDefaultSew = readType & ~gather16;
  wire [1:0]        _dataSplitSew_T_11 = useDefaultSew ? instReg_sew : 2'h0;
  wire [1:0]        dataSplitSew = {_dataSplitSew_T_11[1], _dataSplitSew_T_11[0] | unitType[3] & subType[1] | gather16} | {allGroupExecute, 1'h0};
  wire              sourceDataUseDefaultSew = ~(unitType[3] | gather16);
  wire [1:0]        _sourceDataEEW_T_6 = (sourceDataUseDefaultSew ? instReg_sew : 2'h0) | (unitType[3] ? instReg_sew >> subType[2:1] : 2'h0);
  wire [1:0]        sourceDataEEW = {_sourceDataEEW_T_6[1], _sourceDataEEW_T_6[0] | gather16};
  wire [3:0]        executeIndexGrowth = 4'h1 << dataSplitSew;
  wire [1:0]        lastExecuteIndex = {2{executeIndexGrowth[0]}} | {executeIndexGrowth[1], 1'h0};
  wire [3:0]        _sourceDataEEW1H_T = 4'h1 << sourceDataEEW;
  wire [2:0]        sourceDataEEW1H = _sourceDataEEW1H_T[2:0];
  wire [7:0]        lastElementIndex = instReg_vl[7:0] - {7'h0, |instReg_vl};
  wire [7:0]        processingVl_lastByteIndex = lastElementIndex;
  wire              maskFormatSource = ffo | maskDestinationType;
  wire [3:0]        processingVl_lastGroupRemaining = processingVl_lastByteIndex[3:0];
  wire [3:0]        processingVl_0_1 = processingVl_lastByteIndex[7:4];
  wire [1:0]        processingVl_lastLaneIndex = processingVl_lastGroupRemaining[3:2];
  wire [3:0]        _processingVl_lastGroupDataNeed_T = 4'h1 << processingVl_lastLaneIndex;
  wire [2:0]        _GEN_3 = _processingVl_lastGroupDataNeed_T[2:0] | _processingVl_lastGroupDataNeed_T[3:1];
  wire [3:0]        processingVl_0_2 = {_processingVl_lastGroupDataNeed_T[3], _GEN_3[2], _GEN_3[1:0] | {_processingVl_lastGroupDataNeed_T[3], _GEN_3[2]}};
  wire [8:0]        processingVl_lastByteIndex_1 = {lastElementIndex, 1'h0};
  wire [3:0]        processingVl_lastGroupRemaining_1 = processingVl_lastByteIndex_1[3:0];
  wire [4:0]        processingVl_1_1 = processingVl_lastByteIndex_1[8:4];
  wire [1:0]        processingVl_lastLaneIndex_1 = processingVl_lastGroupRemaining_1[3:2];
  wire [3:0]        _processingVl_lastGroupDataNeed_T_5 = 4'h1 << processingVl_lastLaneIndex_1;
  wire [2:0]        _GEN_4 = _processingVl_lastGroupDataNeed_T_5[2:0] | _processingVl_lastGroupDataNeed_T_5[3:1];
  wire [3:0]        processingVl_1_2 = {_processingVl_lastGroupDataNeed_T_5[3], _GEN_4[2], _GEN_4[1:0] | {_processingVl_lastGroupDataNeed_T_5[3], _GEN_4[2]}};
  wire [9:0]        processingVl_lastByteIndex_2 = {lastElementIndex, 2'h0};
  wire [3:0]        processingVl_lastGroupRemaining_2 = processingVl_lastByteIndex_2[3:0];
  wire [5:0]        processingVl_2_1 = processingVl_lastByteIndex_2[9:4];
  wire [1:0]        processingVl_lastLaneIndex_2 = processingVl_lastGroupRemaining_2[3:2];
  wire [3:0]        _processingVl_lastGroupDataNeed_T_10 = 4'h1 << processingVl_lastLaneIndex_2;
  wire [2:0]        _GEN_5 = _processingVl_lastGroupDataNeed_T_10[2:0] | _processingVl_lastGroupDataNeed_T_10[3:1];
  wire [3:0]        processingVl_2_2 = {_processingVl_lastGroupDataNeed_T_10[3], _GEN_5[2], _GEN_5[1:0] | {_processingVl_lastGroupDataNeed_T_10[3], _GEN_5[2]}};
  wire [6:0]        processingMaskVl_lastGroupRemaining = lastElementIndex[6:0];
  wire [6:0]        elementTailForMaskDestination = lastElementIndex[6:0];
  wire              processingMaskVl_lastGroupMisAlign = |processingMaskVl_lastGroupRemaining;
  wire              processingMaskVl_0_1 = lastElementIndex[7];
  wire [1:0]        processingMaskVl_lastLaneIndex = processingMaskVl_lastGroupRemaining[6:5] - {1'h0, processingMaskVl_lastGroupRemaining[4:0] == 5'h0};
  wire [3:0]        _processingMaskVl_dataNeedForPL_T = 4'h1 << processingMaskVl_lastLaneIndex;
  wire [2:0]        _GEN_6 = _processingMaskVl_dataNeedForPL_T[2:0] | _processingMaskVl_dataNeedForPL_T[3:1];
  wire [3:0]        processingMaskVl_dataNeedForPL = {_processingMaskVl_dataNeedForPL_T[3], _GEN_6[2], _GEN_6[1:0] | {_processingMaskVl_dataNeedForPL_T[3], _GEN_6[2]}};
  wire              processingMaskVl_dataNeedForNPL_misAlign = |(processingMaskVl_lastGroupRemaining[1:0]);
  wire [5:0]        processingMaskVl_dataNeedForNPL_datapathSize = {1'h0, processingMaskVl_lastGroupRemaining[6:2]} + {5'h0, processingMaskVl_dataNeedForNPL_misAlign};
  wire              processingMaskVl_dataNeedForNPL_allNeed = |(processingMaskVl_dataNeedForNPL_datapathSize[5:2]);
  wire [1:0]        processingMaskVl_dataNeedForNPL_lastLaneIndex = processingMaskVl_dataNeedForNPL_datapathSize[1:0];
  wire [3:0]        _processingMaskVl_dataNeedForNPL_dataNeed_T = 4'h1 << processingMaskVl_dataNeedForNPL_lastLaneIndex;
  wire [3:0]        _processingMaskVl_dataNeedForNPL_dataNeed_T_3 = _processingMaskVl_dataNeedForNPL_dataNeed_T | {_processingMaskVl_dataNeedForNPL_dataNeed_T[2:0], 1'h0};
  wire [3:0]        processingMaskVl_dataNeedForNPL_dataNeed = ~(_processingMaskVl_dataNeedForNPL_dataNeed_T_3 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_3[1:0], 2'h0}) | {4{processingMaskVl_dataNeedForNPL_allNeed}};
  wire              processingMaskVl_dataNeedForNPL_misAlign_1 = processingMaskVl_lastGroupRemaining[0];
  wire [6:0]        processingMaskVl_dataNeedForNPL_datapathSize_1 = {1'h0, processingMaskVl_lastGroupRemaining[6:1]} + {6'h0, processingMaskVl_dataNeedForNPL_misAlign_1};
  wire              processingMaskVl_dataNeedForNPL_allNeed_1 = |(processingMaskVl_dataNeedForNPL_datapathSize_1[6:2]);
  wire [1:0]        processingMaskVl_dataNeedForNPL_lastLaneIndex_1 = processingMaskVl_dataNeedForNPL_datapathSize_1[1:0];
  wire [3:0]        _processingMaskVl_dataNeedForNPL_dataNeed_T_10 = 4'h1 << processingMaskVl_dataNeedForNPL_lastLaneIndex_1;
  wire [3:0]        _processingMaskVl_dataNeedForNPL_dataNeed_T_13 = _processingMaskVl_dataNeedForNPL_dataNeed_T_10 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_10[2:0], 1'h0};
  wire [3:0]        processingMaskVl_dataNeedForNPL_dataNeed_1 = ~(_processingMaskVl_dataNeedForNPL_dataNeed_T_13 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_13[1:0], 2'h0}) | {4{processingMaskVl_dataNeedForNPL_allNeed_1}};
  wire [7:0]        processingMaskVl_dataNeedForNPL_datapathSize_2 = {1'h0, processingMaskVl_lastGroupRemaining};
  wire              processingMaskVl_dataNeedForNPL_allNeed_2 = |(processingMaskVl_dataNeedForNPL_datapathSize_2[7:2]);
  wire [1:0]        processingMaskVl_dataNeedForNPL_lastLaneIndex_2 = processingMaskVl_dataNeedForNPL_datapathSize_2[1:0];
  wire [3:0]        _processingMaskVl_dataNeedForNPL_dataNeed_T_20 = 4'h1 << processingMaskVl_dataNeedForNPL_lastLaneIndex_2;
  wire [3:0]        _processingMaskVl_dataNeedForNPL_dataNeed_T_23 = _processingMaskVl_dataNeedForNPL_dataNeed_T_20 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_20[2:0], 1'h0};
  wire [3:0]        processingMaskVl_dataNeedForNPL_dataNeed_2 = ~(_processingMaskVl_dataNeedForNPL_dataNeed_T_23 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_23[1:0], 2'h0}) | {4{processingMaskVl_dataNeedForNPL_allNeed_2}};
  wire [3:0]        processingMaskVl_dataNeedForNPL =
    (sew1H[0] ? processingMaskVl_dataNeedForNPL_dataNeed : 4'h0) | (sew1H[1] ? processingMaskVl_dataNeedForNPL_dataNeed_1 : 4'h0) | (sew1H[2] ? processingMaskVl_dataNeedForNPL_dataNeed_2 : 4'h0);
  wire [3:0]        processingMaskVl_0_2 = ffo ? processingMaskVl_dataNeedForPL : processingMaskVl_dataNeedForNPL;
  wire              reduceLastDataNeed_vlMSB = |(reduceLastDataNeed_byteForVl[8:4]);
  wire [3:0]        reduceLastDataNeed_vlLSB = instReg_vl[3:0];
  wire [3:0]        reduceLastDataNeed_vlLSB_1 = instReg_vl[3:0];
  wire [3:0]        reduceLastDataNeed_vlLSB_2 = instReg_vl[3:0];
  wire [1:0]        reduceLastDataNeed_lsbDSize = reduceLastDataNeed_vlLSB[3:2] - {1'h0, reduceLastDataNeed_vlLSB[1:0] == 2'h0};
  wire [3:0]        _reduceLastDataNeed_T = 4'h1 << reduceLastDataNeed_lsbDSize;
  wire [2:0]        _GEN_7 = _reduceLastDataNeed_T[2:0] | _reduceLastDataNeed_T[3:1];
  wire [9:0]        reduceLastDataNeed_byteForVl_1 = {instReg_vl, 1'h0};
  wire              reduceLastDataNeed_vlMSB_1 = |(reduceLastDataNeed_byteForVl_1[9:4]);
  wire [1:0]        reduceLastDataNeed_lsbDSize_1 = reduceLastDataNeed_vlLSB_1[3:2] - {1'h0, reduceLastDataNeed_vlLSB_1[1:0] == 2'h0};
  wire [3:0]        _reduceLastDataNeed_T_8 = 4'h1 << reduceLastDataNeed_lsbDSize_1;
  wire [2:0]        _GEN_8 = _reduceLastDataNeed_T_8[2:0] | _reduceLastDataNeed_T_8[3:1];
  wire [10:0]       reduceLastDataNeed_byteForVl_2 = {instReg_vl, 2'h0};
  wire              reduceLastDataNeed_vlMSB_2 = |(reduceLastDataNeed_byteForVl_2[10:4]);
  wire [1:0]        reduceLastDataNeed_lsbDSize_2 = reduceLastDataNeed_vlLSB_2[3:2] - {1'h0, reduceLastDataNeed_vlLSB_2[1:0] == 2'h0};
  wire [3:0]        _reduceLastDataNeed_T_16 = 4'h1 << reduceLastDataNeed_lsbDSize_2;
  wire [2:0]        _GEN_9 = _reduceLastDataNeed_T_16[2:0] | _reduceLastDataNeed_T_16[3:1];
  wire [3:0]        reduceLastDataNeed =
    (sew1H[0] ? {_reduceLastDataNeed_T[3], _GEN_7[2], _GEN_7[1:0] | {_reduceLastDataNeed_T[3], _GEN_7[2]}} | {4{reduceLastDataNeed_vlMSB}} : 4'h0)
    | (sew1H[1] ? {_reduceLastDataNeed_T_8[3], _GEN_8[2], _GEN_8[1:0] | {_reduceLastDataNeed_T_8[3], _GEN_8[2]}} | {4{reduceLastDataNeed_vlMSB_1}} : 4'h0)
    | (sew1H[2] ? {_reduceLastDataNeed_T_16[3], _GEN_9[2], _GEN_9[1:0] | {_reduceLastDataNeed_T_16[3], _GEN_9[2]}} | {4{reduceLastDataNeed_vlMSB_2}} : 4'h0);
  wire [1:0]        dataSourceSew = unitType[3] ? instReg_sew - instReg_decodeResult_topUop[2:1] : gather16 ? 2'h1 : instReg_sew;
  wire [3:0]        _dataSourceSew1H_T = 4'h1 << dataSourceSew;
  wire [2:0]        dataSourceSew1H = _dataSourceSew1H_T[2:0];
  wire              unorderReduce = ~orderReduce & unitType[2];
  wire              normalFormat = ~maskFormatSource & ~unorderReduce & ~mv;
  wire [5:0]        lastGroupForInstruction =
    {1'h0, {1'h0, {3'h0, maskFormatSource & processingMaskVl_0_1} | (normalFormat & dataSourceSew1H[0] ? processingVl_0_1 : 4'h0)} | (normalFormat & dataSourceSew1H[1] ? processingVl_1_1 : 5'h0)}
    | (normalFormat & dataSourceSew1H[2] ? processingVl_2_1 : 6'h0);
  wire [2:0]        popDataNeed_dataPathGroups = lastElementIndex[7:5];
  wire [1:0]        popDataNeed_lastLaneIndex = popDataNeed_dataPathGroups[1:0];
  wire              popDataNeed_lagerThanDLen = popDataNeed_dataPathGroups[2];
  wire [3:0]        _popDataNeed_T = 4'h1 << popDataNeed_lastLaneIndex;
  wire [2:0]        _GEN_10 = _popDataNeed_T[2:0] | _popDataNeed_T[3:1];
  wire [3:0]        popDataNeed = {_popDataNeed_T[3], _GEN_10[2], _GEN_10[1:0] | {_popDataNeed_T[3], _GEN_10[2]}} | {4{popDataNeed_lagerThanDLen}};
  wire [3:0]        lastGroupDataNeed =
    (unorderReduce & instReg_decodeResult_popCount ? popDataNeed : 4'h0) | (unorderReduce & ~instReg_decodeResult_popCount ? reduceLastDataNeed : 4'h0) | (maskFormatSource ? processingMaskVl_0_2 : 4'h0)
    | (normalFormat & dataSourceSew1H[0] ? processingVl_0_2 : 4'h0) | (normalFormat & dataSourceSew1H[1] ? processingVl_1_2 : 4'h0) | (normalFormat & dataSourceSew1H[2] ? processingVl_2_2 : 4'h0);
  wire [3:0]        exeRequestQueue_queue_dataIn_lo = {exeRequestQueue_0_enq_bits_index, exeRequestQueue_0_enq_bits_ffo};
  wire [63:0]       exeRequestQueue_queue_dataIn_hi = {exeRequestQueue_0_enq_bits_source1, exeRequestQueue_0_enq_bits_source2};
  wire [67:0]       exeRequestQueue_queue_dataIn = {exeRequestQueue_queue_dataIn_hi, exeRequestQueue_queue_dataIn_lo};
  wire              exeRequestQueue_queue_dataOut_ffo = _exeRequestQueue_queue_fifo_data_out[0];
  wire [2:0]        exeRequestQueue_queue_dataOut_index = _exeRequestQueue_queue_fifo_data_out[3:1];
  wire [31:0]       exeRequestQueue_queue_dataOut_source2 = _exeRequestQueue_queue_fifo_data_out[35:4];
  wire [31:0]       exeRequestQueue_queue_dataOut_source1 = _exeRequestQueue_queue_fifo_data_out[67:36];
  wire              exeRequestQueue_0_enq_ready = ~_exeRequestQueue_queue_fifo_full;
  wire              exeRequestQueue_0_deq_ready;
  wire              exeRequestQueue_0_deq_valid = ~_exeRequestQueue_queue_fifo_empty | exeRequestQueue_0_enq_valid;
  wire [31:0]       exeRequestQueue_0_deq_bits_source1 = _exeRequestQueue_queue_fifo_empty ? exeRequestQueue_0_enq_bits_source1 : exeRequestQueue_queue_dataOut_source1;
  wire [31:0]       exeRequestQueue_0_deq_bits_source2 = _exeRequestQueue_queue_fifo_empty ? exeRequestQueue_0_enq_bits_source2 : exeRequestQueue_queue_dataOut_source2;
  wire [2:0]        exeRequestQueue_0_deq_bits_index = _exeRequestQueue_queue_fifo_empty ? exeRequestQueue_0_enq_bits_index : exeRequestQueue_queue_dataOut_index;
  wire              exeRequestQueue_0_deq_bits_ffo = _exeRequestQueue_queue_fifo_empty ? exeRequestQueue_0_enq_bits_ffo : exeRequestQueue_queue_dataOut_ffo;
  wire              tokenIO_0_maskRequestRelease_0 = exeRequestQueue_0_deq_ready & exeRequestQueue_0_deq_valid;
  wire [3:0]        exeRequestQueue_queue_dataIn_lo_1 = {exeRequestQueue_1_enq_bits_index, exeRequestQueue_1_enq_bits_ffo};
  wire [63:0]       exeRequestQueue_queue_dataIn_hi_1 = {exeRequestQueue_1_enq_bits_source1, exeRequestQueue_1_enq_bits_source2};
  wire [67:0]       exeRequestQueue_queue_dataIn_1 = {exeRequestQueue_queue_dataIn_hi_1, exeRequestQueue_queue_dataIn_lo_1};
  wire              exeRequestQueue_queue_dataOut_1_ffo = _exeRequestQueue_queue_fifo_1_data_out[0];
  wire [2:0]        exeRequestQueue_queue_dataOut_1_index = _exeRequestQueue_queue_fifo_1_data_out[3:1];
  wire [31:0]       exeRequestQueue_queue_dataOut_1_source2 = _exeRequestQueue_queue_fifo_1_data_out[35:4];
  wire [31:0]       exeRequestQueue_queue_dataOut_1_source1 = _exeRequestQueue_queue_fifo_1_data_out[67:36];
  wire              exeRequestQueue_1_enq_ready = ~_exeRequestQueue_queue_fifo_1_full;
  wire              exeRequestQueue_1_deq_ready;
  wire              exeRequestQueue_1_deq_valid = ~_exeRequestQueue_queue_fifo_1_empty | exeRequestQueue_1_enq_valid;
  wire [31:0]       exeRequestQueue_1_deq_bits_source1 = _exeRequestQueue_queue_fifo_1_empty ? exeRequestQueue_1_enq_bits_source1 : exeRequestQueue_queue_dataOut_1_source1;
  wire [31:0]       exeRequestQueue_1_deq_bits_source2 = _exeRequestQueue_queue_fifo_1_empty ? exeRequestQueue_1_enq_bits_source2 : exeRequestQueue_queue_dataOut_1_source2;
  wire [2:0]        exeRequestQueue_1_deq_bits_index = _exeRequestQueue_queue_fifo_1_empty ? exeRequestQueue_1_enq_bits_index : exeRequestQueue_queue_dataOut_1_index;
  wire              exeRequestQueue_1_deq_bits_ffo = _exeRequestQueue_queue_fifo_1_empty ? exeRequestQueue_1_enq_bits_ffo : exeRequestQueue_queue_dataOut_1_ffo;
  wire              tokenIO_1_maskRequestRelease_0 = exeRequestQueue_1_deq_ready & exeRequestQueue_1_deq_valid;
  wire [3:0]        exeRequestQueue_queue_dataIn_lo_2 = {exeRequestQueue_2_enq_bits_index, exeRequestQueue_2_enq_bits_ffo};
  wire [63:0]       exeRequestQueue_queue_dataIn_hi_2 = {exeRequestQueue_2_enq_bits_source1, exeRequestQueue_2_enq_bits_source2};
  wire [67:0]       exeRequestQueue_queue_dataIn_2 = {exeRequestQueue_queue_dataIn_hi_2, exeRequestQueue_queue_dataIn_lo_2};
  wire              exeRequestQueue_queue_dataOut_2_ffo = _exeRequestQueue_queue_fifo_2_data_out[0];
  wire [2:0]        exeRequestQueue_queue_dataOut_2_index = _exeRequestQueue_queue_fifo_2_data_out[3:1];
  wire [31:0]       exeRequestQueue_queue_dataOut_2_source2 = _exeRequestQueue_queue_fifo_2_data_out[35:4];
  wire [31:0]       exeRequestQueue_queue_dataOut_2_source1 = _exeRequestQueue_queue_fifo_2_data_out[67:36];
  wire              exeRequestQueue_2_enq_ready = ~_exeRequestQueue_queue_fifo_2_full;
  wire              exeRequestQueue_2_deq_ready;
  wire              exeRequestQueue_2_deq_valid = ~_exeRequestQueue_queue_fifo_2_empty | exeRequestQueue_2_enq_valid;
  wire [31:0]       exeRequestQueue_2_deq_bits_source1 = _exeRequestQueue_queue_fifo_2_empty ? exeRequestQueue_2_enq_bits_source1 : exeRequestQueue_queue_dataOut_2_source1;
  wire [31:0]       exeRequestQueue_2_deq_bits_source2 = _exeRequestQueue_queue_fifo_2_empty ? exeRequestQueue_2_enq_bits_source2 : exeRequestQueue_queue_dataOut_2_source2;
  wire [2:0]        exeRequestQueue_2_deq_bits_index = _exeRequestQueue_queue_fifo_2_empty ? exeRequestQueue_2_enq_bits_index : exeRequestQueue_queue_dataOut_2_index;
  wire              exeRequestQueue_2_deq_bits_ffo = _exeRequestQueue_queue_fifo_2_empty ? exeRequestQueue_2_enq_bits_ffo : exeRequestQueue_queue_dataOut_2_ffo;
  wire              tokenIO_2_maskRequestRelease_0 = exeRequestQueue_2_deq_ready & exeRequestQueue_2_deq_valid;
  wire [3:0]        exeRequestQueue_queue_dataIn_lo_3 = {exeRequestQueue_3_enq_bits_index, exeRequestQueue_3_enq_bits_ffo};
  wire [63:0]       exeRequestQueue_queue_dataIn_hi_3 = {exeRequestQueue_3_enq_bits_source1, exeRequestQueue_3_enq_bits_source2};
  wire [67:0]       exeRequestQueue_queue_dataIn_3 = {exeRequestQueue_queue_dataIn_hi_3, exeRequestQueue_queue_dataIn_lo_3};
  wire              exeRequestQueue_queue_dataOut_3_ffo = _exeRequestQueue_queue_fifo_3_data_out[0];
  wire [2:0]        exeRequestQueue_queue_dataOut_3_index = _exeRequestQueue_queue_fifo_3_data_out[3:1];
  wire [31:0]       exeRequestQueue_queue_dataOut_3_source2 = _exeRequestQueue_queue_fifo_3_data_out[35:4];
  wire [31:0]       exeRequestQueue_queue_dataOut_3_source1 = _exeRequestQueue_queue_fifo_3_data_out[67:36];
  wire              exeRequestQueue_3_enq_ready = ~_exeRequestQueue_queue_fifo_3_full;
  wire              exeRequestQueue_3_deq_ready;
  wire              exeRequestQueue_3_deq_valid = ~_exeRequestQueue_queue_fifo_3_empty | exeRequestQueue_3_enq_valid;
  wire [31:0]       exeRequestQueue_3_deq_bits_source1 = _exeRequestQueue_queue_fifo_3_empty ? exeRequestQueue_3_enq_bits_source1 : exeRequestQueue_queue_dataOut_3_source1;
  wire [31:0]       exeRequestQueue_3_deq_bits_source2 = _exeRequestQueue_queue_fifo_3_empty ? exeRequestQueue_3_enq_bits_source2 : exeRequestQueue_queue_dataOut_3_source2;
  wire [2:0]        exeRequestQueue_3_deq_bits_index = _exeRequestQueue_queue_fifo_3_empty ? exeRequestQueue_3_enq_bits_index : exeRequestQueue_queue_dataOut_3_index;
  wire              exeRequestQueue_3_deq_bits_ffo = _exeRequestQueue_queue_fifo_3_empty ? exeRequestQueue_3_enq_bits_ffo : exeRequestQueue_queue_dataOut_3_ffo;
  wire              tokenIO_3_maskRequestRelease_0 = exeRequestQueue_3_deq_ready & exeRequestQueue_3_deq_valid;
  reg               exeReqReg_0_valid;
  reg  [31:0]       exeReqReg_0_bits_source1;
  reg  [31:0]       exeReqReg_0_bits_source2;
  reg  [2:0]        exeReqReg_0_bits_index;
  reg               exeReqReg_0_bits_ffo;
  reg               exeReqReg_1_valid;
  reg  [31:0]       exeReqReg_1_bits_source1;
  reg  [31:0]       exeReqReg_1_bits_source2;
  reg  [2:0]        exeReqReg_1_bits_index;
  reg               exeReqReg_1_bits_ffo;
  reg               exeReqReg_2_valid;
  reg  [31:0]       exeReqReg_2_bits_source1;
  reg  [31:0]       exeReqReg_2_bits_source2;
  reg  [2:0]        exeReqReg_2_bits_index;
  reg               exeReqReg_2_bits_ffo;
  reg               exeReqReg_3_valid;
  reg  [31:0]       exeReqReg_3_bits_source1;
  reg  [31:0]       exeReqReg_3_bits_source2;
  reg  [2:0]        exeReqReg_3_bits_index;
  reg               exeReqReg_3_bits_ffo;
  reg  [4:0]        requestCounter;
  wire [5:0]        _GEN_11 = {1'h0, requestCounter};
  wire              counterValid = _GEN_11 <= lastGroupForInstruction;
  wire              lastGroup = _GEN_11 == lastGroupForInstruction | ~orderReduce & unitType[2] | mv;
  wire [127:0]      slideAddressGen_slideMaskInput_lo = {slideAddressGen_slideMaskInput_lo_hi, slideAddressGen_slideMaskInput_lo_lo};
  wire [127:0]      slideAddressGen_slideMaskInput_hi = {slideAddressGen_slideMaskInput_hi_hi, slideAddressGen_slideMaskInput_hi_lo};
  wire [63:0][3:0]  _GEN_12 =
    {{slideAddressGen_slideMaskInput_hi[127:124]},
     {slideAddressGen_slideMaskInput_hi[123:120]},
     {slideAddressGen_slideMaskInput_hi[119:116]},
     {slideAddressGen_slideMaskInput_hi[115:112]},
     {slideAddressGen_slideMaskInput_hi[111:108]},
     {slideAddressGen_slideMaskInput_hi[107:104]},
     {slideAddressGen_slideMaskInput_hi[103:100]},
     {slideAddressGen_slideMaskInput_hi[99:96]},
     {slideAddressGen_slideMaskInput_hi[95:92]},
     {slideAddressGen_slideMaskInput_hi[91:88]},
     {slideAddressGen_slideMaskInput_hi[87:84]},
     {slideAddressGen_slideMaskInput_hi[83:80]},
     {slideAddressGen_slideMaskInput_hi[79:76]},
     {slideAddressGen_slideMaskInput_hi[75:72]},
     {slideAddressGen_slideMaskInput_hi[71:68]},
     {slideAddressGen_slideMaskInput_hi[67:64]},
     {slideAddressGen_slideMaskInput_hi[63:60]},
     {slideAddressGen_slideMaskInput_hi[59:56]},
     {slideAddressGen_slideMaskInput_hi[55:52]},
     {slideAddressGen_slideMaskInput_hi[51:48]},
     {slideAddressGen_slideMaskInput_hi[47:44]},
     {slideAddressGen_slideMaskInput_hi[43:40]},
     {slideAddressGen_slideMaskInput_hi[39:36]},
     {slideAddressGen_slideMaskInput_hi[35:32]},
     {slideAddressGen_slideMaskInput_hi[31:28]},
     {slideAddressGen_slideMaskInput_hi[27:24]},
     {slideAddressGen_slideMaskInput_hi[23:20]},
     {slideAddressGen_slideMaskInput_hi[19:16]},
     {slideAddressGen_slideMaskInput_hi[15:12]},
     {slideAddressGen_slideMaskInput_hi[11:8]},
     {slideAddressGen_slideMaskInput_hi[7:4]},
     {slideAddressGen_slideMaskInput_hi[3:0]},
     {slideAddressGen_slideMaskInput_lo[127:124]},
     {slideAddressGen_slideMaskInput_lo[123:120]},
     {slideAddressGen_slideMaskInput_lo[119:116]},
     {slideAddressGen_slideMaskInput_lo[115:112]},
     {slideAddressGen_slideMaskInput_lo[111:108]},
     {slideAddressGen_slideMaskInput_lo[107:104]},
     {slideAddressGen_slideMaskInput_lo[103:100]},
     {slideAddressGen_slideMaskInput_lo[99:96]},
     {slideAddressGen_slideMaskInput_lo[95:92]},
     {slideAddressGen_slideMaskInput_lo[91:88]},
     {slideAddressGen_slideMaskInput_lo[87:84]},
     {slideAddressGen_slideMaskInput_lo[83:80]},
     {slideAddressGen_slideMaskInput_lo[79:76]},
     {slideAddressGen_slideMaskInput_lo[75:72]},
     {slideAddressGen_slideMaskInput_lo[71:68]},
     {slideAddressGen_slideMaskInput_lo[67:64]},
     {slideAddressGen_slideMaskInput_lo[63:60]},
     {slideAddressGen_slideMaskInput_lo[59:56]},
     {slideAddressGen_slideMaskInput_lo[55:52]},
     {slideAddressGen_slideMaskInput_lo[51:48]},
     {slideAddressGen_slideMaskInput_lo[47:44]},
     {slideAddressGen_slideMaskInput_lo[43:40]},
     {slideAddressGen_slideMaskInput_lo[39:36]},
     {slideAddressGen_slideMaskInput_lo[35:32]},
     {slideAddressGen_slideMaskInput_lo[31:28]},
     {slideAddressGen_slideMaskInput_lo[27:24]},
     {slideAddressGen_slideMaskInput_lo[23:20]},
     {slideAddressGen_slideMaskInput_lo[19:16]},
     {slideAddressGen_slideMaskInput_lo[15:12]},
     {slideAddressGen_slideMaskInput_lo[11:8]},
     {slideAddressGen_slideMaskInput_lo[7:4]},
     {slideAddressGen_slideMaskInput_lo[3:0]}};
  wire              lastExecuteGroupDeq;
  wire              viotaCounterAdd;
  wire              groupCounterAdd = noSource ? viotaCounterAdd : lastExecuteGroupDeq;
  wire [3:0]        groupDataNeed = lastGroup ? lastGroupDataNeed : 4'hF;
  reg  [1:0]        executeIndex;
  reg  [3:0]        readIssueStageState_groupReadState;
  reg  [3:0]        readIssueStageState_needRead;
  wire [3:0]        readWaitQueue_enq_bits_needRead = readIssueStageState_needRead;
  reg  [3:0]        readIssueStageState_elementValid;
  wire [3:0]        readWaitQueue_enq_bits_sourceValid = readIssueStageState_elementValid;
  reg  [3:0]        readIssueStageState_replaceVs1;
  wire [3:0]        readWaitQueue_enq_bits_replaceVs1 = readIssueStageState_replaceVs1;
  reg  [3:0]        readIssueStageState_readOffset;
  reg  [1:0]        readIssueStageState_accessLane_0;
  reg  [1:0]        readIssueStageState_accessLane_1;
  wire [1:0]        selectExecuteReq_1_bits_readLane = readIssueStageState_accessLane_1;
  reg  [1:0]        readIssueStageState_accessLane_2;
  wire [1:0]        selectExecuteReq_2_bits_readLane = readIssueStageState_accessLane_2;
  reg  [1:0]        readIssueStageState_accessLane_3;
  wire [1:0]        selectExecuteReq_3_bits_readLane = readIssueStageState_accessLane_3;
  reg  [2:0]        readIssueStageState_vsGrowth_0;
  reg  [2:0]        readIssueStageState_vsGrowth_1;
  reg  [2:0]        readIssueStageState_vsGrowth_2;
  reg  [2:0]        readIssueStageState_vsGrowth_3;
  reg  [6:0]        readIssueStageState_executeGroup;
  wire [6:0]        readWaitQueue_enq_bits_executeGroup = readIssueStageState_executeGroup;
  reg  [7:0]        readIssueStageState_readDataOffset;
  reg               readIssueStageState_last;
  wire              readWaitQueue_enq_bits_last = readIssueStageState_last;
  reg               readIssueStageValid;
  wire [2:0]        accessCountQueue_enq_bits_0 = accessCountEnq_0;
  wire [2:0]        accessCountQueue_enq_bits_1 = accessCountEnq_1;
  wire [2:0]        accessCountQueue_enq_bits_2 = accessCountEnq_2;
  wire [2:0]        accessCountQueue_enq_bits_3 = accessCountEnq_3;
  wire              readIssueStageEnq;
  wire              accessCountQueue_deq_valid;
  assign accessCountQueue_deq_valid = ~_accessCountQueue_fifo_empty;
  wire [2:0]        accessCountQueue_dataOut_0;
  wire [2:0]        accessCountQueue_dataOut_1;
  wire [2:0]        accessCountQueue_dataOut_2;
  wire [2:0]        accessCountQueue_dataOut_3;
  wire [5:0]        accessCountQueue_dataIn_lo = {accessCountQueue_enq_bits_1, accessCountQueue_enq_bits_0};
  wire [5:0]        accessCountQueue_dataIn_hi = {accessCountQueue_enq_bits_3, accessCountQueue_enq_bits_2};
  wire [11:0]       accessCountQueue_dataIn = {accessCountQueue_dataIn_hi, accessCountQueue_dataIn_lo};
  assign accessCountQueue_dataOut_0 = _accessCountQueue_fifo_data_out[2:0];
  assign accessCountQueue_dataOut_1 = _accessCountQueue_fifo_data_out[5:3];
  assign accessCountQueue_dataOut_2 = _accessCountQueue_fifo_data_out[8:6];
  assign accessCountQueue_dataOut_3 = _accessCountQueue_fifo_data_out[11:9];
  wire [2:0]        accessCountQueue_deq_bits_0 = accessCountQueue_dataOut_0;
  wire [2:0]        accessCountQueue_deq_bits_1 = accessCountQueue_dataOut_1;
  wire [2:0]        accessCountQueue_deq_bits_2 = accessCountQueue_dataOut_2;
  wire [2:0]        accessCountQueue_deq_bits_3 = accessCountQueue_dataOut_3;
  wire              accessCountQueue_enq_ready = ~_accessCountQueue_fifo_full;
  wire              accessCountQueue_enq_valid;
  wire              accessCountQueue_deq_ready;
  wire [6:0]        _extendGroupCount_T_1 = {requestCounter, executeIndex};
  wire [6:0]        _executeGroup_T_8 = executeIndexGrowth[0] ? _extendGroupCount_T_1 : 7'h0;
  wire [5:0]        _GEN_13 = _executeGroup_T_8[5:0] | (executeIndexGrowth[1] ? {requestCounter, executeIndex[1]} : 6'h0);
  wire [6:0]        executeGroup = {_executeGroup_T_8[6], _GEN_13[5], _GEN_13[4:0] | (executeIndexGrowth[2] ? requestCounter : 5'h0)};
  wire              vlMisAlign;
  assign vlMisAlign = |(instReg_vl[1:0]);
  wire [6:0]        lastexecuteGroup = instReg_vl[8:2] - {6'h0, ~vlMisAlign};
  wire              isVlBoundary = executeGroup == lastexecuteGroup;
  wire              validExecuteGroup = executeGroup <= lastexecuteGroup;
  wire [3:0]        _maskSplit_vlBoundaryCorrection_T_37 = 4'h1 << instReg_vl[1:0];
  wire [3:0]        _vlBoundaryCorrection_T_5 = _maskSplit_vlBoundaryCorrection_T_37 | {_maskSplit_vlBoundaryCorrection_T_37[2:0], 1'h0};
  wire [3:0]        vlBoundaryCorrection = ~({4{vlMisAlign & isVlBoundary}} & (_vlBoundaryCorrection_T_5 | {_vlBoundaryCorrection_T_5[1:0], 2'h0})) & {4{validExecuteGroup}};
  wire [127:0]      selectReadStageMask_lo = {selectReadStageMask_lo_hi, selectReadStageMask_lo_lo};
  wire [127:0]      selectReadStageMask_hi = {selectReadStageMask_hi_hi, selectReadStageMask_hi_lo};
  wire [63:0][3:0]  _GEN_14 =
    {{selectReadStageMask_hi[127:124]},
     {selectReadStageMask_hi[123:120]},
     {selectReadStageMask_hi[119:116]},
     {selectReadStageMask_hi[115:112]},
     {selectReadStageMask_hi[111:108]},
     {selectReadStageMask_hi[107:104]},
     {selectReadStageMask_hi[103:100]},
     {selectReadStageMask_hi[99:96]},
     {selectReadStageMask_hi[95:92]},
     {selectReadStageMask_hi[91:88]},
     {selectReadStageMask_hi[87:84]},
     {selectReadStageMask_hi[83:80]},
     {selectReadStageMask_hi[79:76]},
     {selectReadStageMask_hi[75:72]},
     {selectReadStageMask_hi[71:68]},
     {selectReadStageMask_hi[67:64]},
     {selectReadStageMask_hi[63:60]},
     {selectReadStageMask_hi[59:56]},
     {selectReadStageMask_hi[55:52]},
     {selectReadStageMask_hi[51:48]},
     {selectReadStageMask_hi[47:44]},
     {selectReadStageMask_hi[43:40]},
     {selectReadStageMask_hi[39:36]},
     {selectReadStageMask_hi[35:32]},
     {selectReadStageMask_hi[31:28]},
     {selectReadStageMask_hi[27:24]},
     {selectReadStageMask_hi[23:20]},
     {selectReadStageMask_hi[19:16]},
     {selectReadStageMask_hi[15:12]},
     {selectReadStageMask_hi[11:8]},
     {selectReadStageMask_hi[7:4]},
     {selectReadStageMask_hi[3:0]},
     {selectReadStageMask_lo[127:124]},
     {selectReadStageMask_lo[123:120]},
     {selectReadStageMask_lo[119:116]},
     {selectReadStageMask_lo[115:112]},
     {selectReadStageMask_lo[111:108]},
     {selectReadStageMask_lo[107:104]},
     {selectReadStageMask_lo[103:100]},
     {selectReadStageMask_lo[99:96]},
     {selectReadStageMask_lo[95:92]},
     {selectReadStageMask_lo[91:88]},
     {selectReadStageMask_lo[87:84]},
     {selectReadStageMask_lo[83:80]},
     {selectReadStageMask_lo[79:76]},
     {selectReadStageMask_lo[75:72]},
     {selectReadStageMask_lo[71:68]},
     {selectReadStageMask_lo[67:64]},
     {selectReadStageMask_lo[63:60]},
     {selectReadStageMask_lo[59:56]},
     {selectReadStageMask_lo[55:52]},
     {selectReadStageMask_lo[51:48]},
     {selectReadStageMask_lo[47:44]},
     {selectReadStageMask_lo[43:40]},
     {selectReadStageMask_lo[39:36]},
     {selectReadStageMask_lo[35:32]},
     {selectReadStageMask_lo[31:28]},
     {selectReadStageMask_lo[27:24]},
     {selectReadStageMask_lo[23:20]},
     {selectReadStageMask_lo[19:16]},
     {selectReadStageMask_lo[15:12]},
     {selectReadStageMask_lo[11:8]},
     {selectReadStageMask_lo[7:4]},
     {selectReadStageMask_lo[3:0]}};
  wire [3:0]        readMaskCorrection = (instReg_maskType ? _GEN_14[executeGroup[5:0]] : 4'hF) & vlBoundaryCorrection;
  wire [127:0]      maskSplit_maskSelect_lo = {maskSplit_maskSelect_lo_hi, maskSplit_maskSelect_lo_lo};
  wire [127:0]      maskSplit_maskSelect_hi = {maskSplit_maskSelect_hi_hi, maskSplit_maskSelect_hi_lo};
  wire [4:0]        executeGroupCounter;
  wire              maskSplit_vlMisAlign = |(instReg_vl[3:0]);
  wire [4:0]        maskSplit_lastexecuteGroup = instReg_vl[8:4] - {4'h0, ~maskSplit_vlMisAlign};
  wire              maskSplit_isVlBoundary = executeGroupCounter == maskSplit_lastexecuteGroup;
  wire              maskSplit_validExecuteGroup = executeGroupCounter <= maskSplit_lastexecuteGroup;
  wire [15:0]       _maskSplit_vlBoundaryCorrection_T_2 = 16'h1 << instReg_vl[3:0];
  wire [15:0]       _maskSplit_vlBoundaryCorrection_T_5 = _maskSplit_vlBoundaryCorrection_T_2 | {_maskSplit_vlBoundaryCorrection_T_2[14:0], 1'h0};
  wire [15:0]       _maskSplit_vlBoundaryCorrection_T_8 = _maskSplit_vlBoundaryCorrection_T_5 | {_maskSplit_vlBoundaryCorrection_T_5[13:0], 2'h0};
  wire [15:0]       _maskSplit_vlBoundaryCorrection_T_11 = _maskSplit_vlBoundaryCorrection_T_8 | {_maskSplit_vlBoundaryCorrection_T_8[11:0], 4'h0};
  wire [15:0]       maskSplit_vlBoundaryCorrection = ~({16{maskSplit_vlMisAlign & maskSplit_isVlBoundary}} & (_maskSplit_vlBoundaryCorrection_T_11 | {_maskSplit_vlBoundaryCorrection_T_11[7:0], 8'h0})) & {16{maskSplit_validExecuteGroup}};
  wire [15:0][15:0] _GEN_15 =
    {{maskSplit_maskSelect_hi[127:112]},
     {maskSplit_maskSelect_hi[111:96]},
     {maskSplit_maskSelect_hi[95:80]},
     {maskSplit_maskSelect_hi[79:64]},
     {maskSplit_maskSelect_hi[63:48]},
     {maskSplit_maskSelect_hi[47:32]},
     {maskSplit_maskSelect_hi[31:16]},
     {maskSplit_maskSelect_hi[15:0]},
     {maskSplit_maskSelect_lo[127:112]},
     {maskSplit_maskSelect_lo[111:96]},
     {maskSplit_maskSelect_lo[95:80]},
     {maskSplit_maskSelect_lo[79:64]},
     {maskSplit_maskSelect_lo[63:48]},
     {maskSplit_maskSelect_lo[47:32]},
     {maskSplit_maskSelect_lo[31:16]},
     {maskSplit_maskSelect_lo[15:0]}};
  wire [15:0]       maskSplit_0_2 = (instReg_maskType ? _GEN_15[executeGroupCounter[3:0]] : 16'hFFFF) & maskSplit_vlBoundaryCorrection;
  wire [1:0]        maskSplit_byteMask_lo_lo_lo = maskSplit_0_2[1:0];
  wire [1:0]        maskSplit_byteMask_lo_lo_hi = maskSplit_0_2[3:2];
  wire [3:0]        maskSplit_byteMask_lo_lo = {maskSplit_byteMask_lo_lo_hi, maskSplit_byteMask_lo_lo_lo};
  wire [1:0]        maskSplit_byteMask_lo_hi_lo = maskSplit_0_2[5:4];
  wire [1:0]        maskSplit_byteMask_lo_hi_hi = maskSplit_0_2[7:6];
  wire [3:0]        maskSplit_byteMask_lo_hi = {maskSplit_byteMask_lo_hi_hi, maskSplit_byteMask_lo_hi_lo};
  wire [7:0]        maskSplit_byteMask_lo = {maskSplit_byteMask_lo_hi, maskSplit_byteMask_lo_lo};
  wire [1:0]        maskSplit_byteMask_hi_lo_lo = maskSplit_0_2[9:8];
  wire [1:0]        maskSplit_byteMask_hi_lo_hi = maskSplit_0_2[11:10];
  wire [3:0]        maskSplit_byteMask_hi_lo = {maskSplit_byteMask_hi_lo_hi, maskSplit_byteMask_hi_lo_lo};
  wire [1:0]        maskSplit_byteMask_hi_hi_lo = maskSplit_0_2[13:12];
  wire [1:0]        maskSplit_byteMask_hi_hi_hi = maskSplit_0_2[15:14];
  wire [3:0]        maskSplit_byteMask_hi_hi = {maskSplit_byteMask_hi_hi_hi, maskSplit_byteMask_hi_hi_lo};
  wire [7:0]        maskSplit_byteMask_hi = {maskSplit_byteMask_hi_hi, maskSplit_byteMask_hi_lo};
  wire [15:0]       maskSplit_0_1 = {maskSplit_byteMask_hi, maskSplit_byteMask_lo};
  wire [127:0]      maskSplit_maskSelect_lo_1 = {maskSplit_maskSelect_lo_hi_1, maskSplit_maskSelect_lo_lo_1};
  wire [127:0]      maskSplit_maskSelect_hi_1 = {maskSplit_maskSelect_hi_hi_1, maskSplit_maskSelect_hi_lo_1};
  wire              maskSplit_vlMisAlign_1 = |(instReg_vl[2:0]);
  wire [5:0]        maskSplit_lastexecuteGroup_1 = instReg_vl[8:3] - {5'h0, ~maskSplit_vlMisAlign_1};
  wire [5:0]        _GEN_16 = {1'h0, executeGroupCounter};
  wire              maskSplit_isVlBoundary_1 = _GEN_16 == maskSplit_lastexecuteGroup_1;
  wire              maskSplit_validExecuteGroup_1 = _GEN_16 <= maskSplit_lastexecuteGroup_1;
  wire [7:0]        _maskSplit_vlBoundaryCorrection_T_21 = 8'h1 << instReg_vl[2:0];
  wire [7:0]        _maskSplit_vlBoundaryCorrection_T_24 = _maskSplit_vlBoundaryCorrection_T_21 | {_maskSplit_vlBoundaryCorrection_T_21[6:0], 1'h0};
  wire [7:0]        _maskSplit_vlBoundaryCorrection_T_27 = _maskSplit_vlBoundaryCorrection_T_24 | {_maskSplit_vlBoundaryCorrection_T_24[5:0], 2'h0};
  wire [7:0]        maskSplit_vlBoundaryCorrection_1 =
    ~({8{maskSplit_vlMisAlign_1 & maskSplit_isVlBoundary_1}} & (_maskSplit_vlBoundaryCorrection_T_27 | {_maskSplit_vlBoundaryCorrection_T_27[3:0], 4'h0})) & {8{maskSplit_validExecuteGroup_1}};
  wire [31:0][7:0]  _GEN_17 =
    {{maskSplit_maskSelect_hi_1[127:120]},
     {maskSplit_maskSelect_hi_1[119:112]},
     {maskSplit_maskSelect_hi_1[111:104]},
     {maskSplit_maskSelect_hi_1[103:96]},
     {maskSplit_maskSelect_hi_1[95:88]},
     {maskSplit_maskSelect_hi_1[87:80]},
     {maskSplit_maskSelect_hi_1[79:72]},
     {maskSplit_maskSelect_hi_1[71:64]},
     {maskSplit_maskSelect_hi_1[63:56]},
     {maskSplit_maskSelect_hi_1[55:48]},
     {maskSplit_maskSelect_hi_1[47:40]},
     {maskSplit_maskSelect_hi_1[39:32]},
     {maskSplit_maskSelect_hi_1[31:24]},
     {maskSplit_maskSelect_hi_1[23:16]},
     {maskSplit_maskSelect_hi_1[15:8]},
     {maskSplit_maskSelect_hi_1[7:0]},
     {maskSplit_maskSelect_lo_1[127:120]},
     {maskSplit_maskSelect_lo_1[119:112]},
     {maskSplit_maskSelect_lo_1[111:104]},
     {maskSplit_maskSelect_lo_1[103:96]},
     {maskSplit_maskSelect_lo_1[95:88]},
     {maskSplit_maskSelect_lo_1[87:80]},
     {maskSplit_maskSelect_lo_1[79:72]},
     {maskSplit_maskSelect_lo_1[71:64]},
     {maskSplit_maskSelect_lo_1[63:56]},
     {maskSplit_maskSelect_lo_1[55:48]},
     {maskSplit_maskSelect_lo_1[47:40]},
     {maskSplit_maskSelect_lo_1[39:32]},
     {maskSplit_maskSelect_lo_1[31:24]},
     {maskSplit_maskSelect_lo_1[23:16]},
     {maskSplit_maskSelect_lo_1[15:8]},
     {maskSplit_maskSelect_lo_1[7:0]}};
  wire [7:0]        maskSplit_1_2 = (instReg_maskType ? _GEN_17[executeGroupCounter] : 8'hFF) & maskSplit_vlBoundaryCorrection_1;
  wire [3:0]        maskSplit_byteMask_lo_lo_1 = {{2{maskSplit_1_2[1]}}, {2{maskSplit_1_2[0]}}};
  wire [3:0]        maskSplit_byteMask_lo_hi_1 = {{2{maskSplit_1_2[3]}}, {2{maskSplit_1_2[2]}}};
  wire [7:0]        maskSplit_byteMask_lo_1 = {maskSplit_byteMask_lo_hi_1, maskSplit_byteMask_lo_lo_1};
  wire [3:0]        maskSplit_byteMask_hi_lo_1 = {{2{maskSplit_1_2[5]}}, {2{maskSplit_1_2[4]}}};
  wire [3:0]        maskSplit_byteMask_hi_hi_1 = {{2{maskSplit_1_2[7]}}, {2{maskSplit_1_2[6]}}};
  wire [7:0]        maskSplit_byteMask_hi_1 = {maskSplit_byteMask_hi_hi_1, maskSplit_byteMask_hi_lo_1};
  wire [15:0]       maskSplit_1_1 = {maskSplit_byteMask_hi_1, maskSplit_byteMask_lo_1};
  wire [127:0]      maskSplit_maskSelect_lo_2 = {maskSplit_maskSelect_lo_hi_2, maskSplit_maskSelect_lo_lo_2};
  wire [127:0]      maskSplit_maskSelect_hi_2 = {maskSplit_maskSelect_hi_hi_2, maskSplit_maskSelect_hi_lo_2};
  wire              maskSplit_vlMisAlign_2;
  assign maskSplit_vlMisAlign_2 = |(instReg_vl[1:0]);
  wire [6:0]        maskSplit_lastexecuteGroup_2 = instReg_vl[8:2] - {6'h0, ~maskSplit_vlMisAlign_2};
  wire [6:0]        _GEN_18 = {2'h0, executeGroupCounter};
  wire              maskSplit_isVlBoundary_2 = _GEN_18 == maskSplit_lastexecuteGroup_2;
  wire              maskSplit_validExecuteGroup_2 = _GEN_18 <= maskSplit_lastexecuteGroup_2;
  wire [3:0]        _maskSplit_vlBoundaryCorrection_T_40 = _maskSplit_vlBoundaryCorrection_T_37 | {_maskSplit_vlBoundaryCorrection_T_37[2:0], 1'h0};
  wire [3:0]        maskSplit_vlBoundaryCorrection_2 =
    ~({4{maskSplit_vlMisAlign_2 & maskSplit_isVlBoundary_2}} & (_maskSplit_vlBoundaryCorrection_T_40 | {_maskSplit_vlBoundaryCorrection_T_40[1:0], 2'h0})) & {4{maskSplit_validExecuteGroup_2}};
  wire [31:0][3:0]  _GEN_19 =
    {{maskSplit_maskSelect_lo_2[127:124]},
     {maskSplit_maskSelect_lo_2[123:120]},
     {maskSplit_maskSelect_lo_2[119:116]},
     {maskSplit_maskSelect_lo_2[115:112]},
     {maskSplit_maskSelect_lo_2[111:108]},
     {maskSplit_maskSelect_lo_2[107:104]},
     {maskSplit_maskSelect_lo_2[103:100]},
     {maskSplit_maskSelect_lo_2[99:96]},
     {maskSplit_maskSelect_lo_2[95:92]},
     {maskSplit_maskSelect_lo_2[91:88]},
     {maskSplit_maskSelect_lo_2[87:84]},
     {maskSplit_maskSelect_lo_2[83:80]},
     {maskSplit_maskSelect_lo_2[79:76]},
     {maskSplit_maskSelect_lo_2[75:72]},
     {maskSplit_maskSelect_lo_2[71:68]},
     {maskSplit_maskSelect_lo_2[67:64]},
     {maskSplit_maskSelect_lo_2[63:60]},
     {maskSplit_maskSelect_lo_2[59:56]},
     {maskSplit_maskSelect_lo_2[55:52]},
     {maskSplit_maskSelect_lo_2[51:48]},
     {maskSplit_maskSelect_lo_2[47:44]},
     {maskSplit_maskSelect_lo_2[43:40]},
     {maskSplit_maskSelect_lo_2[39:36]},
     {maskSplit_maskSelect_lo_2[35:32]},
     {maskSplit_maskSelect_lo_2[31:28]},
     {maskSplit_maskSelect_lo_2[27:24]},
     {maskSplit_maskSelect_lo_2[23:20]},
     {maskSplit_maskSelect_lo_2[19:16]},
     {maskSplit_maskSelect_lo_2[15:12]},
     {maskSplit_maskSelect_lo_2[11:8]},
     {maskSplit_maskSelect_lo_2[7:4]},
     {maskSplit_maskSelect_lo_2[3:0]}};
  wire [3:0]        maskSplit_2_2 = (instReg_maskType ? _GEN_19[executeGroupCounter] : 4'hF) & maskSplit_vlBoundaryCorrection_2;
  wire [7:0]        maskSplit_byteMask_lo_2 = {{4{maskSplit_2_2[1]}}, {4{maskSplit_2_2[0]}}};
  wire [7:0]        maskSplit_byteMask_hi_2 = {{4{maskSplit_2_2[3]}}, {4{maskSplit_2_2[2]}}};
  wire [15:0]       maskSplit_2_1 = {maskSplit_byteMask_hi_2, maskSplit_byteMask_lo_2};
  wire [15:0]       executeByteMask = (sew1H[0] ? maskSplit_0_1 : 16'h0) | (sew1H[1] ? maskSplit_1_1 : 16'h0) | (sew1H[2] ? maskSplit_2_1 : 16'h0);
  wire [15:0]       _executeElementMask_T_3 = sew1H[0] ? maskSplit_0_2 : 16'h0;
  wire [7:0]        _GEN_20 = _executeElementMask_T_3[7:0] | (sew1H[1] ? maskSplit_1_2 : 8'h0);
  wire [15:0]       executeElementMask = {_executeElementMask_T_3[15:8], _GEN_20[7:4], _GEN_20[3:0] | (sew1H[2] ? maskSplit_2_2 : 4'h0)};
  wire [127:0]      maskForDestination_lo = {maskForDestination_lo_hi, maskForDestination_lo_lo};
  wire [127:0]      maskForDestination_hi = {maskForDestination_hi_hi, maskForDestination_hi_lo};
  wire              vs1Split_vs1SetIndex = requestCounter[0];
  wire [127:0]      _lastGroupMask_T = 128'h1 << elementTailForMaskDestination;
  wire [126:0]      _GEN_21 = _lastGroupMask_T[126:0] | _lastGroupMask_T[127:1];
  wire [125:0]      _GEN_22 = _GEN_21[125:0] | {_lastGroupMask_T[127], _GEN_21[126:2]};
  wire [123:0]      _GEN_23 = _GEN_22[123:0] | {_lastGroupMask_T[127], _GEN_21[126], _GEN_22[125:4]};
  wire [119:0]      _GEN_24 = _GEN_23[119:0] | {_lastGroupMask_T[127], _GEN_21[126], _GEN_22[125:124], _GEN_23[123:8]};
  wire [111:0]      _GEN_25 = _GEN_24[111:0] | {_lastGroupMask_T[127], _GEN_21[126], _GEN_22[125:124], _GEN_23[123:120], _GEN_24[119:16]};
  wire [95:0]       _GEN_26 = _GEN_25[95:0] | {_lastGroupMask_T[127], _GEN_21[126], _GEN_22[125:124], _GEN_23[123:120], _GEN_24[119:112], _GEN_25[111:32]};
  wire [127:0]      lastGroupMask =
    {_lastGroupMask_T[127],
     _GEN_21[126],
     _GEN_22[125:124],
     _GEN_23[123:120],
     _GEN_24[119:112],
     _GEN_25[111:96],
     _GEN_26[95:64],
     _GEN_26[63:0] | {_lastGroupMask_T[127], _GEN_21[126], _GEN_22[125:124], _GEN_23[123:120], _GEN_24[119:112], _GEN_25[111:96], _GEN_26[95:64]}};
  wire [127:0]      currentMaskGroupForDestination =
    (lastGroup ? lastGroupMask : 128'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
    & (instReg_maskType & ~instReg_decodeResult_maskSource ? (vs1Split_vs1SetIndex ? maskForDestination_hi : maskForDestination_lo) : 128'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF);
  wire [63:0]       _GEN_27 = {exeReqReg_1_bits_source1, exeReqReg_0_bits_source1};
  wire [63:0]       groupSourceData_lo;
  assign groupSourceData_lo = _GEN_27;
  wire [63:0]       source1_lo;
  assign source1_lo = _GEN_27;
  wire [63:0]       _GEN_28 = {exeReqReg_3_bits_source1, exeReqReg_2_bits_source1};
  wire [63:0]       groupSourceData_hi;
  assign groupSourceData_hi = _GEN_28;
  wire [63:0]       source1_hi;
  assign source1_hi = _GEN_28;
  wire [127:0]      groupSourceData = {groupSourceData_hi, groupSourceData_lo};
  wire [1:0]        _GEN_29 = {exeReqReg_1_valid, exeReqReg_0_valid};
  wire [1:0]        groupSourceValid_lo;
  assign groupSourceValid_lo = _GEN_29;
  wire [1:0]        view__in_bits_validInput_lo;
  assign view__in_bits_validInput_lo = _GEN_29;
  wire [1:0]        view__in_bits_sourceValid_lo;
  assign view__in_bits_sourceValid_lo = _GEN_29;
  wire [1:0]        _GEN_30 = {exeReqReg_3_valid, exeReqReg_2_valid};
  wire [1:0]        groupSourceValid_hi;
  assign groupSourceValid_hi = _GEN_30;
  wire [1:0]        view__in_bits_validInput_hi;
  assign view__in_bits_validInput_hi = _GEN_30;
  wire [1:0]        view__in_bits_sourceValid_hi;
  assign view__in_bits_sourceValid_hi = _GEN_30;
  wire [3:0]        groupSourceValid = {groupSourceValid_hi, groupSourceValid_lo};
  wire [1:0]        shifterSize = (sourceDataEEW1H[0] ? executeIndex : 2'h0) | (sourceDataEEW1H[1] ? {executeIndex[1], 1'h0} : 2'h0);
  wire [3:0]        _shifterSource_T = 4'h1 << shifterSize;
  wire [127:0]      _shifterSource_T_8 = _shifterSource_T[0] ? groupSourceData : 128'h0;
  wire [95:0]       _GEN_31 = _shifterSource_T_8[95:0] | (_shifterSource_T[1] ? groupSourceData[127:32] : 96'h0);
  wire [63:0]       _GEN_32 = _GEN_31[63:0] | (_shifterSource_T[2] ? groupSourceData[127:64] : 64'h0);
  wire [127:0]      shifterSource = {_shifterSource_T_8[127:96], _GEN_31[95:64], _GEN_32[63:32], _GEN_32[31:0] | (_shifterSource_T[3] ? groupSourceData[127:96] : 32'h0)};
  wire [7:0]        selectValid_lo = {{4{groupSourceValid[1]}}, {4{groupSourceValid[0]}}};
  wire [7:0]        selectValid_hi = {{4{groupSourceValid[3]}}, {4{groupSourceValid[2]}}};
  wire [3:0]        selectValid_lo_1 = {{2{groupSourceValid[1]}}, {2{groupSourceValid[0]}}};
  wire [3:0]        selectValid_hi_1 = {{2{groupSourceValid[3]}}, {2{groupSourceValid[2]}}};
  wire [3:0][3:0]   _GEN_33 = {{selectValid_hi[7:4]}, {selectValid_hi[3:0]}, {selectValid_lo[7:4]}, {selectValid_lo[3:0]}};
  wire [3:0]        selectValid = (sourceDataEEW1H[0] ? _GEN_33[executeIndex] : 4'h0) | (sourceDataEEW1H[1] ? (executeIndex[1] ? selectValid_hi_1 : selectValid_lo_1) : 4'h0) | (sourceDataEEW1H[2] ? groupSourceValid : 4'h0);
  wire [31:0]       source_0 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[7:0] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[15:0] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[31:0] : 32'h0);
  wire [31:0]       source_1 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[15:8] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[31:16] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[63:32] : 32'h0);
  wire [31:0]       source_2 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[23:16] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[47:32] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[95:64] : 32'h0);
  wire [31:0]       source_3 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[31:24] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[63:48] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[127:96] : 32'h0);
  wire [3:0]        _GEN_34 = selectValid & readMaskCorrection;
  wire [3:0]        checkVec_validVec;
  assign checkVec_validVec = _GEN_34;
  wire [3:0]        checkVec_validVec_1;
  assign checkVec_validVec_1 = _GEN_34;
  wire [3:0]        checkVec_validVec_2;
  assign checkVec_validVec_2 = _GEN_34;
  wire              checkVec_checkResultVec_0_6 = checkVec_validVec[0];
  wire [3:0]        _GEN_35 = 4'h1 << instReg_vlmul[1:0];
  wire [3:0]        checkVec_checkResultVec_intLMULInput;
  assign checkVec_checkResultVec_intLMULInput = _GEN_35;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_1;
  assign checkVec_checkResultVec_intLMULInput_1 = _GEN_35;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_2;
  assign checkVec_checkResultVec_intLMULInput_2 = _GEN_35;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_3;
  assign checkVec_checkResultVec_intLMULInput_3 = _GEN_35;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_4;
  assign checkVec_checkResultVec_intLMULInput_4 = _GEN_35;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_5;
  assign checkVec_checkResultVec_intLMULInput_5 = _GEN_35;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_6;
  assign checkVec_checkResultVec_intLMULInput_6 = _GEN_35;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_7;
  assign checkVec_checkResultVec_intLMULInput_7 = _GEN_35;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_8;
  assign checkVec_checkResultVec_intLMULInput_8 = _GEN_35;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_9;
  assign checkVec_checkResultVec_intLMULInput_9 = _GEN_35;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_10;
  assign checkVec_checkResultVec_intLMULInput_10 = _GEN_35;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_11;
  assign checkVec_checkResultVec_intLMULInput_11 = _GEN_35;
  wire [7:0]        checkVec_checkResultVec_dataPosition = source_0[7:0];
  wire [3:0]        checkVec_checkResultVec_0_0 = 4'h1 << checkVec_checkResultVec_dataPosition[1:0];
  wire [1:0]        checkVec_checkResultVec_0_1 = checkVec_checkResultVec_dataPosition[1:0];
  wire [1:0]        checkVec_checkResultVec_0_2 = checkVec_checkResultVec_dataPosition[3:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup = checkVec_checkResultVec_dataPosition[7:4];
  wire              checkVec_checkResultVec_0_3 = checkVec_checkResultVec_dataGroup[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth = checkVec_checkResultVec_dataGroup[3:1];
  wire [2:0]        checkVec_checkResultVec_0_4 = checkVec_checkResultVec_accessRegGrowth;
  wire [2:0]        checkVec_checkResultVec_decimalProportion = {checkVec_checkResultVec_0_3, checkVec_checkResultVec_0_2};
  wire [2:0]        checkVec_checkResultVec_decimal = checkVec_checkResultVec_decimalProportion;
  wire              checkVec_checkResultVec_overlap =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal >= checkVec_checkResultVec_intLMULInput[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth} >= checkVec_checkResultVec_intLMULInput, source_0[31:8]};
  wire              checkVec_checkResultVec_0_5 = checkVec_checkResultVec_overlap | ~checkVec_checkResultVec_0_6;
  wire              checkVec_checkResultVec_1_6 = checkVec_validVec[1];
  wire [7:0]        checkVec_checkResultVec_dataPosition_1 = source_1[7:0];
  wire [3:0]        checkVec_checkResultVec_1_0 = 4'h1 << checkVec_checkResultVec_dataPosition_1[1:0];
  wire [1:0]        checkVec_checkResultVec_1_1 = checkVec_checkResultVec_dataPosition_1[1:0];
  wire [1:0]        checkVec_checkResultVec_1_2 = checkVec_checkResultVec_dataPosition_1[3:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_1 = checkVec_checkResultVec_dataPosition_1[7:4];
  wire              checkVec_checkResultVec_1_3 = checkVec_checkResultVec_dataGroup_1[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_1 = checkVec_checkResultVec_dataGroup_1[3:1];
  wire [2:0]        checkVec_checkResultVec_1_4 = checkVec_checkResultVec_accessRegGrowth_1;
  wire [2:0]        checkVec_checkResultVec_decimalProportion_1 = {checkVec_checkResultVec_1_3, checkVec_checkResultVec_1_2};
  wire [2:0]        checkVec_checkResultVec_decimal_1 = checkVec_checkResultVec_decimalProportion_1;
  wire              checkVec_checkResultVec_overlap_1 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_1 >= checkVec_checkResultVec_intLMULInput_1[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_1} >= checkVec_checkResultVec_intLMULInput_1, source_1[31:8]};
  wire              checkVec_checkResultVec_1_5 = checkVec_checkResultVec_overlap_1 | ~checkVec_checkResultVec_1_6;
  wire              checkVec_checkResultVec_2_6 = checkVec_validVec[2];
  wire [7:0]        checkVec_checkResultVec_dataPosition_2 = source_2[7:0];
  wire [3:0]        checkVec_checkResultVec_2_0 = 4'h1 << checkVec_checkResultVec_dataPosition_2[1:0];
  wire [1:0]        checkVec_checkResultVec_2_1 = checkVec_checkResultVec_dataPosition_2[1:0];
  wire [1:0]        checkVec_checkResultVec_2_2 = checkVec_checkResultVec_dataPosition_2[3:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_2 = checkVec_checkResultVec_dataPosition_2[7:4];
  wire              checkVec_checkResultVec_2_3 = checkVec_checkResultVec_dataGroup_2[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_2 = checkVec_checkResultVec_dataGroup_2[3:1];
  wire [2:0]        checkVec_checkResultVec_2_4 = checkVec_checkResultVec_accessRegGrowth_2;
  wire [2:0]        checkVec_checkResultVec_decimalProportion_2 = {checkVec_checkResultVec_2_3, checkVec_checkResultVec_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_2 = checkVec_checkResultVec_decimalProportion_2;
  wire              checkVec_checkResultVec_overlap_2 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_2 >= checkVec_checkResultVec_intLMULInput_2[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_2} >= checkVec_checkResultVec_intLMULInput_2, source_2[31:8]};
  wire              checkVec_checkResultVec_2_5 = checkVec_checkResultVec_overlap_2 | ~checkVec_checkResultVec_2_6;
  wire              checkVec_checkResultVec_3_6 = checkVec_validVec[3];
  wire [7:0]        checkVec_checkResultVec_dataPosition_3 = source_3[7:0];
  wire [3:0]        checkVec_checkResultVec_3_0 = 4'h1 << checkVec_checkResultVec_dataPosition_3[1:0];
  wire [1:0]        checkVec_checkResultVec_3_1 = checkVec_checkResultVec_dataPosition_3[1:0];
  wire [1:0]        checkVec_checkResultVec_3_2 = checkVec_checkResultVec_dataPosition_3[3:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_3 = checkVec_checkResultVec_dataPosition_3[7:4];
  wire              checkVec_checkResultVec_3_3 = checkVec_checkResultVec_dataGroup_3[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_3 = checkVec_checkResultVec_dataGroup_3[3:1];
  wire [2:0]        checkVec_checkResultVec_3_4 = checkVec_checkResultVec_accessRegGrowth_3;
  wire [2:0]        checkVec_checkResultVec_decimalProportion_3 = {checkVec_checkResultVec_3_3, checkVec_checkResultVec_3_2};
  wire [2:0]        checkVec_checkResultVec_decimal_3 = checkVec_checkResultVec_decimalProportion_3;
  wire              checkVec_checkResultVec_overlap_3 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_3 >= checkVec_checkResultVec_intLMULInput_3[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_3} >= checkVec_checkResultVec_intLMULInput_3, source_3[31:8]};
  wire              checkVec_checkResultVec_3_5 = checkVec_checkResultVec_overlap_3 | ~checkVec_checkResultVec_3_6;
  wire [7:0]        checkVec_checkResult_lo = {checkVec_checkResultVec_1_0, checkVec_checkResultVec_0_0};
  wire [7:0]        checkVec_checkResult_hi = {checkVec_checkResultVec_3_0, checkVec_checkResultVec_2_0};
  wire [15:0]       checkVec_0_0 = {checkVec_checkResult_hi, checkVec_checkResult_lo};
  wire [3:0]        checkVec_checkResult_lo_1 = {checkVec_checkResultVec_1_1, checkVec_checkResultVec_0_1};
  wire [3:0]        checkVec_checkResult_hi_1 = {checkVec_checkResultVec_3_1, checkVec_checkResultVec_2_1};
  wire [7:0]        checkVec_0_1 = {checkVec_checkResult_hi_1, checkVec_checkResult_lo_1};
  wire [3:0]        checkVec_checkResult_lo_2 = {checkVec_checkResultVec_1_2, checkVec_checkResultVec_0_2};
  wire [3:0]        checkVec_checkResult_hi_2 = {checkVec_checkResultVec_3_2, checkVec_checkResultVec_2_2};
  wire [7:0]        checkVec_0_2 = {checkVec_checkResult_hi_2, checkVec_checkResult_lo_2};
  wire [1:0]        checkVec_checkResult_lo_3 = {checkVec_checkResultVec_1_3, checkVec_checkResultVec_0_3};
  wire [1:0]        checkVec_checkResult_hi_3 = {checkVec_checkResultVec_3_3, checkVec_checkResultVec_2_3};
  wire [3:0]        checkVec_0_3 = {checkVec_checkResult_hi_3, checkVec_checkResult_lo_3};
  wire [5:0]        checkVec_checkResult_lo_4 = {checkVec_checkResultVec_1_4, checkVec_checkResultVec_0_4};
  wire [5:0]        checkVec_checkResult_hi_4 = {checkVec_checkResultVec_3_4, checkVec_checkResultVec_2_4};
  wire [11:0]       checkVec_0_4 = {checkVec_checkResult_hi_4, checkVec_checkResult_lo_4};
  wire [1:0]        checkVec_checkResult_lo_5 = {checkVec_checkResultVec_1_5, checkVec_checkResultVec_0_5};
  wire [1:0]        checkVec_checkResult_hi_5 = {checkVec_checkResultVec_3_5, checkVec_checkResultVec_2_5};
  wire [3:0]        checkVec_0_5 = {checkVec_checkResult_hi_5, checkVec_checkResult_lo_5};
  wire [1:0]        checkVec_checkResult_lo_6 = {checkVec_checkResultVec_1_6, checkVec_checkResultVec_0_6};
  wire [1:0]        checkVec_checkResult_hi_6 = {checkVec_checkResultVec_3_6, checkVec_checkResultVec_2_6};
  wire [3:0]        checkVec_0_6 = {checkVec_checkResult_hi_6, checkVec_checkResult_lo_6};
  wire              checkVec_checkResultVec_0_6_1 = checkVec_validVec_1[0];
  wire [7:0]        checkVec_checkResultVec_dataPosition_4 = {source_0[6:0], 1'h0};
  wire [1:0]        _checkVec_checkResultVec_accessMask_T_35 = 2'h1 << checkVec_checkResultVec_dataPosition_4[1];
  wire [3:0]        checkVec_checkResultVec_0_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_35[1]}}, {2{_checkVec_checkResultVec_accessMask_T_35[0]}}};
  wire [1:0]        checkVec_checkResultVec_0_1_1 = {checkVec_checkResultVec_dataPosition_4[1], 1'h0};
  wire [1:0]        checkVec_checkResultVec_0_2_1 = checkVec_checkResultVec_dataPosition_4[3:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_4 = checkVec_checkResultVec_dataPosition_4[7:4];
  wire              checkVec_checkResultVec_0_3_1 = checkVec_checkResultVec_dataGroup_4[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_4 = checkVec_checkResultVec_dataGroup_4[3:1];
  wire [2:0]        checkVec_checkResultVec_0_4_1 = checkVec_checkResultVec_accessRegGrowth_4;
  wire [2:0]        checkVec_checkResultVec_decimalProportion_4 = {checkVec_checkResultVec_0_3_1, checkVec_checkResultVec_0_2_1};
  wire [2:0]        checkVec_checkResultVec_decimal_4 = checkVec_checkResultVec_decimalProportion_4;
  wire              checkVec_checkResultVec_overlap_4 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_4 >= checkVec_checkResultVec_intLMULInput_4[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_4} >= checkVec_checkResultVec_intLMULInput_4, source_0[31:8]};
  wire              checkVec_checkResultVec_0_5_1 = checkVec_checkResultVec_overlap_4 | ~checkVec_checkResultVec_0_6_1;
  wire              checkVec_checkResultVec_1_6_1 = checkVec_validVec_1[1];
  wire [7:0]        checkVec_checkResultVec_dataPosition_5 = {source_1[6:0], 1'h0};
  wire [1:0]        _checkVec_checkResultVec_accessMask_T_43 = 2'h1 << checkVec_checkResultVec_dataPosition_5[1];
  wire [3:0]        checkVec_checkResultVec_1_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_43[1]}}, {2{_checkVec_checkResultVec_accessMask_T_43[0]}}};
  wire [1:0]        checkVec_checkResultVec_1_1_1 = {checkVec_checkResultVec_dataPosition_5[1], 1'h0};
  wire [1:0]        checkVec_checkResultVec_1_2_1 = checkVec_checkResultVec_dataPosition_5[3:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_5 = checkVec_checkResultVec_dataPosition_5[7:4];
  wire              checkVec_checkResultVec_1_3_1 = checkVec_checkResultVec_dataGroup_5[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_5 = checkVec_checkResultVec_dataGroup_5[3:1];
  wire [2:0]        checkVec_checkResultVec_1_4_1 = checkVec_checkResultVec_accessRegGrowth_5;
  wire [2:0]        checkVec_checkResultVec_decimalProportion_5 = {checkVec_checkResultVec_1_3_1, checkVec_checkResultVec_1_2_1};
  wire [2:0]        checkVec_checkResultVec_decimal_5 = checkVec_checkResultVec_decimalProportion_5;
  wire              checkVec_checkResultVec_overlap_5 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_5 >= checkVec_checkResultVec_intLMULInput_5[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_5} >= checkVec_checkResultVec_intLMULInput_5, source_1[31:8]};
  wire              checkVec_checkResultVec_1_5_1 = checkVec_checkResultVec_overlap_5 | ~checkVec_checkResultVec_1_6_1;
  wire              checkVec_checkResultVec_2_6_1 = checkVec_validVec_1[2];
  wire [7:0]        checkVec_checkResultVec_dataPosition_6 = {source_2[6:0], 1'h0};
  wire [1:0]        _checkVec_checkResultVec_accessMask_T_51 = 2'h1 << checkVec_checkResultVec_dataPosition_6[1];
  wire [3:0]        checkVec_checkResultVec_2_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_51[1]}}, {2{_checkVec_checkResultVec_accessMask_T_51[0]}}};
  wire [1:0]        checkVec_checkResultVec_2_1_1 = {checkVec_checkResultVec_dataPosition_6[1], 1'h0};
  wire [1:0]        checkVec_checkResultVec_2_2_1 = checkVec_checkResultVec_dataPosition_6[3:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_6 = checkVec_checkResultVec_dataPosition_6[7:4];
  wire              checkVec_checkResultVec_2_3_1 = checkVec_checkResultVec_dataGroup_6[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_6 = checkVec_checkResultVec_dataGroup_6[3:1];
  wire [2:0]        checkVec_checkResultVec_2_4_1 = checkVec_checkResultVec_accessRegGrowth_6;
  wire [2:0]        checkVec_checkResultVec_decimalProportion_6 = {checkVec_checkResultVec_2_3_1, checkVec_checkResultVec_2_2_1};
  wire [2:0]        checkVec_checkResultVec_decimal_6 = checkVec_checkResultVec_decimalProportion_6;
  wire              checkVec_checkResultVec_overlap_6 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_6 >= checkVec_checkResultVec_intLMULInput_6[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_6} >= checkVec_checkResultVec_intLMULInput_6, source_2[31:8]};
  wire              checkVec_checkResultVec_2_5_1 = checkVec_checkResultVec_overlap_6 | ~checkVec_checkResultVec_2_6_1;
  wire              checkVec_checkResultVec_3_6_1 = checkVec_validVec_1[3];
  wire [7:0]        checkVec_checkResultVec_dataPosition_7 = {source_3[6:0], 1'h0};
  wire [1:0]        _checkVec_checkResultVec_accessMask_T_59 = 2'h1 << checkVec_checkResultVec_dataPosition_7[1];
  wire [3:0]        checkVec_checkResultVec_3_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_59[1]}}, {2{_checkVec_checkResultVec_accessMask_T_59[0]}}};
  wire [1:0]        checkVec_checkResultVec_3_1_1 = {checkVec_checkResultVec_dataPosition_7[1], 1'h0};
  wire [1:0]        checkVec_checkResultVec_3_2_1 = checkVec_checkResultVec_dataPosition_7[3:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_7 = checkVec_checkResultVec_dataPosition_7[7:4];
  wire              checkVec_checkResultVec_3_3_1 = checkVec_checkResultVec_dataGroup_7[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_7 = checkVec_checkResultVec_dataGroup_7[3:1];
  wire [2:0]        checkVec_checkResultVec_3_4_1 = checkVec_checkResultVec_accessRegGrowth_7;
  wire [2:0]        checkVec_checkResultVec_decimalProportion_7 = {checkVec_checkResultVec_3_3_1, checkVec_checkResultVec_3_2_1};
  wire [2:0]        checkVec_checkResultVec_decimal_7 = checkVec_checkResultVec_decimalProportion_7;
  wire              checkVec_checkResultVec_overlap_7 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_7 >= checkVec_checkResultVec_intLMULInput_7[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_7} >= checkVec_checkResultVec_intLMULInput_7, source_3[31:8]};
  wire              checkVec_checkResultVec_3_5_1 = checkVec_checkResultVec_overlap_7 | ~checkVec_checkResultVec_3_6_1;
  wire [7:0]        checkVec_checkResult_lo_7 = {checkVec_checkResultVec_1_0_1, checkVec_checkResultVec_0_0_1};
  wire [7:0]        checkVec_checkResult_hi_7 = {checkVec_checkResultVec_3_0_1, checkVec_checkResultVec_2_0_1};
  wire [15:0]       checkVec_1_0 = {checkVec_checkResult_hi_7, checkVec_checkResult_lo_7};
  wire [3:0]        checkVec_checkResult_lo_8 = {checkVec_checkResultVec_1_1_1, checkVec_checkResultVec_0_1_1};
  wire [3:0]        checkVec_checkResult_hi_8 = {checkVec_checkResultVec_3_1_1, checkVec_checkResultVec_2_1_1};
  wire [7:0]        checkVec_1_1 = {checkVec_checkResult_hi_8, checkVec_checkResult_lo_8};
  wire [3:0]        checkVec_checkResult_lo_9 = {checkVec_checkResultVec_1_2_1, checkVec_checkResultVec_0_2_1};
  wire [3:0]        checkVec_checkResult_hi_9 = {checkVec_checkResultVec_3_2_1, checkVec_checkResultVec_2_2_1};
  wire [7:0]        checkVec_1_2 = {checkVec_checkResult_hi_9, checkVec_checkResult_lo_9};
  wire [1:0]        checkVec_checkResult_lo_10 = {checkVec_checkResultVec_1_3_1, checkVec_checkResultVec_0_3_1};
  wire [1:0]        checkVec_checkResult_hi_10 = {checkVec_checkResultVec_3_3_1, checkVec_checkResultVec_2_3_1};
  wire [3:0]        checkVec_1_3 = {checkVec_checkResult_hi_10, checkVec_checkResult_lo_10};
  wire [5:0]        checkVec_checkResult_lo_11 = {checkVec_checkResultVec_1_4_1, checkVec_checkResultVec_0_4_1};
  wire [5:0]        checkVec_checkResult_hi_11 = {checkVec_checkResultVec_3_4_1, checkVec_checkResultVec_2_4_1};
  wire [11:0]       checkVec_1_4 = {checkVec_checkResult_hi_11, checkVec_checkResult_lo_11};
  wire [1:0]        checkVec_checkResult_lo_12 = {checkVec_checkResultVec_1_5_1, checkVec_checkResultVec_0_5_1};
  wire [1:0]        checkVec_checkResult_hi_12 = {checkVec_checkResultVec_3_5_1, checkVec_checkResultVec_2_5_1};
  wire [3:0]        checkVec_1_5 = {checkVec_checkResult_hi_12, checkVec_checkResult_lo_12};
  wire [1:0]        checkVec_checkResult_lo_13 = {checkVec_checkResultVec_1_6_1, checkVec_checkResultVec_0_6_1};
  wire [1:0]        checkVec_checkResult_hi_13 = {checkVec_checkResultVec_3_6_1, checkVec_checkResultVec_2_6_1};
  wire [3:0]        checkVec_1_6 = {checkVec_checkResult_hi_13, checkVec_checkResult_lo_13};
  wire              checkVec_checkResultVec_0_6_2 = checkVec_validVec_2[0];
  wire [7:0]        checkVec_checkResultVec_dataPosition_8 = {source_0[5:0], 2'h0};
  wire [1:0]        checkVec_checkResultVec_0_2_2 = checkVec_checkResultVec_dataPosition_8[3:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_8 = checkVec_checkResultVec_dataPosition_8[7:4];
  wire              checkVec_checkResultVec_0_3_2 = checkVec_checkResultVec_dataGroup_8[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_8 = checkVec_checkResultVec_dataGroup_8[3:1];
  wire [2:0]        checkVec_checkResultVec_0_4_2 = checkVec_checkResultVec_accessRegGrowth_8;
  wire [2:0]        checkVec_checkResultVec_decimalProportion_8 = {checkVec_checkResultVec_0_3_2, checkVec_checkResultVec_0_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_8 = checkVec_checkResultVec_decimalProportion_8;
  wire              checkVec_checkResultVec_overlap_8 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_8 >= checkVec_checkResultVec_intLMULInput_8[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_8} >= checkVec_checkResultVec_intLMULInput_8, source_0[31:8]};
  wire              checkVec_checkResultVec_0_5_2 = checkVec_checkResultVec_overlap_8 | ~checkVec_checkResultVec_0_6_2;
  wire              checkVec_checkResultVec_1_6_2 = checkVec_validVec_2[1];
  wire [7:0]        checkVec_checkResultVec_dataPosition_9 = {source_1[5:0], 2'h0};
  wire [1:0]        checkVec_checkResultVec_1_2_2 = checkVec_checkResultVec_dataPosition_9[3:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_9 = checkVec_checkResultVec_dataPosition_9[7:4];
  wire              checkVec_checkResultVec_1_3_2 = checkVec_checkResultVec_dataGroup_9[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_9 = checkVec_checkResultVec_dataGroup_9[3:1];
  wire [2:0]        checkVec_checkResultVec_1_4_2 = checkVec_checkResultVec_accessRegGrowth_9;
  wire [2:0]        checkVec_checkResultVec_decimalProportion_9 = {checkVec_checkResultVec_1_3_2, checkVec_checkResultVec_1_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_9 = checkVec_checkResultVec_decimalProportion_9;
  wire              checkVec_checkResultVec_overlap_9 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_9 >= checkVec_checkResultVec_intLMULInput_9[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_9} >= checkVec_checkResultVec_intLMULInput_9, source_1[31:8]};
  wire              checkVec_checkResultVec_1_5_2 = checkVec_checkResultVec_overlap_9 | ~checkVec_checkResultVec_1_6_2;
  wire              checkVec_checkResultVec_2_6_2 = checkVec_validVec_2[2];
  wire [7:0]        checkVec_checkResultVec_dataPosition_10 = {source_2[5:0], 2'h0};
  wire [1:0]        checkVec_checkResultVec_2_2_2 = checkVec_checkResultVec_dataPosition_10[3:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_10 = checkVec_checkResultVec_dataPosition_10[7:4];
  wire              checkVec_checkResultVec_2_3_2 = checkVec_checkResultVec_dataGroup_10[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_10 = checkVec_checkResultVec_dataGroup_10[3:1];
  wire [2:0]        checkVec_checkResultVec_2_4_2 = checkVec_checkResultVec_accessRegGrowth_10;
  wire [2:0]        checkVec_checkResultVec_decimalProportion_10 = {checkVec_checkResultVec_2_3_2, checkVec_checkResultVec_2_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_10 = checkVec_checkResultVec_decimalProportion_10;
  wire              checkVec_checkResultVec_overlap_10 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_10 >= checkVec_checkResultVec_intLMULInput_10[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_10} >= checkVec_checkResultVec_intLMULInput_10,
      source_2[31:8]};
  wire              checkVec_checkResultVec_2_5_2 = checkVec_checkResultVec_overlap_10 | ~checkVec_checkResultVec_2_6_2;
  wire              checkVec_checkResultVec_3_6_2 = checkVec_validVec_2[3];
  wire [7:0]        checkVec_checkResultVec_dataPosition_11 = {source_3[5:0], 2'h0};
  wire [1:0]        checkVec_checkResultVec_3_2_2 = checkVec_checkResultVec_dataPosition_11[3:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_11 = checkVec_checkResultVec_dataPosition_11[7:4];
  wire              checkVec_checkResultVec_3_3_2 = checkVec_checkResultVec_dataGroup_11[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_11 = checkVec_checkResultVec_dataGroup_11[3:1];
  wire [2:0]        checkVec_checkResultVec_3_4_2 = checkVec_checkResultVec_accessRegGrowth_11;
  wire [2:0]        checkVec_checkResultVec_decimalProportion_11 = {checkVec_checkResultVec_3_3_2, checkVec_checkResultVec_3_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_11 = checkVec_checkResultVec_decimalProportion_11;
  wire              checkVec_checkResultVec_overlap_11 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_11 >= checkVec_checkResultVec_intLMULInput_11[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_11} >= checkVec_checkResultVec_intLMULInput_11,
      source_3[31:8]};
  wire              checkVec_checkResultVec_3_5_2 = checkVec_checkResultVec_overlap_11 | ~checkVec_checkResultVec_3_6_2;
  wire [3:0]        checkVec_checkResult_lo_16 = {checkVec_checkResultVec_1_2_2, checkVec_checkResultVec_0_2_2};
  wire [3:0]        checkVec_checkResult_hi_16 = {checkVec_checkResultVec_3_2_2, checkVec_checkResultVec_2_2_2};
  wire [7:0]        checkVec_2_2 = {checkVec_checkResult_hi_16, checkVec_checkResult_lo_16};
  wire [1:0]        checkVec_checkResult_lo_17 = {checkVec_checkResultVec_1_3_2, checkVec_checkResultVec_0_3_2};
  wire [1:0]        checkVec_checkResult_hi_17 = {checkVec_checkResultVec_3_3_2, checkVec_checkResultVec_2_3_2};
  wire [3:0]        checkVec_2_3 = {checkVec_checkResult_hi_17, checkVec_checkResult_lo_17};
  wire [5:0]        checkVec_checkResult_lo_18 = {checkVec_checkResultVec_1_4_2, checkVec_checkResultVec_0_4_2};
  wire [5:0]        checkVec_checkResult_hi_18 = {checkVec_checkResultVec_3_4_2, checkVec_checkResultVec_2_4_2};
  wire [11:0]       checkVec_2_4 = {checkVec_checkResult_hi_18, checkVec_checkResult_lo_18};
  wire [1:0]        checkVec_checkResult_lo_19 = {checkVec_checkResultVec_1_5_2, checkVec_checkResultVec_0_5_2};
  wire [1:0]        checkVec_checkResult_hi_19 = {checkVec_checkResultVec_3_5_2, checkVec_checkResultVec_2_5_2};
  wire [3:0]        checkVec_2_5 = {checkVec_checkResult_hi_19, checkVec_checkResult_lo_19};
  wire [1:0]        checkVec_checkResult_lo_20 = {checkVec_checkResultVec_1_6_2, checkVec_checkResultVec_0_6_2};
  wire [1:0]        checkVec_checkResult_hi_20 = {checkVec_checkResultVec_3_6_2, checkVec_checkResultVec_2_6_2};
  wire [3:0]        checkVec_2_6 = {checkVec_checkResult_hi_20, checkVec_checkResult_lo_20};
  wire [7:0]        dataOffsetSelect = (sew1H[0] ? checkVec_0_1 : 8'h0) | (sew1H[1] ? checkVec_1_1 : 8'h0);
  wire [7:0]        accessLaneSelect = (sew1H[0] ? checkVec_0_2 : 8'h0) | (sew1H[1] ? checkVec_1_2 : 8'h0) | (sew1H[2] ? checkVec_2_2 : 8'h0);
  wire [3:0]        offsetSelect = (sew1H[0] ? checkVec_0_3 : 4'h0) | (sew1H[1] ? checkVec_1_3 : 4'h0) | (sew1H[2] ? checkVec_2_3 : 4'h0);
  wire [11:0]       growthSelect = (sew1H[0] ? checkVec_0_4 : 12'h0) | (sew1H[1] ? checkVec_1_4 : 12'h0) | (sew1H[2] ? checkVec_2_4 : 12'h0);
  wire [3:0]        notReadSelect = (sew1H[0] ? checkVec_0_5 : 4'h0) | (sew1H[1] ? checkVec_1_5 : 4'h0) | (sew1H[2] ? checkVec_2_5 : 4'h0);
  wire [3:0]        elementValidSelect = (sew1H[0] ? checkVec_0_6 : 4'h0) | (sew1H[1] ? checkVec_1_6 : 4'h0) | (sew1H[2] ? checkVec_2_6 : 4'h0);
  wire              readTypeRequestDeq;
  wire              waiteStageEnqReady;
  wire              readWaitQueue_deq_valid;
  assign readWaitQueue_deq_valid = ~_readWaitQueue_fifo_empty;
  wire [6:0]        readWaitQueue_dataOut_executeGroup;
  wire [3:0]        readWaitQueue_dataOut_sourceValid;
  wire [3:0]        readWaitQueue_dataOut_replaceVs1;
  wire [3:0]        readWaitQueue_dataOut_needRead;
  wire              readWaitQueue_dataOut_last;
  wire [4:0]        readWaitQueue_dataIn_lo = {readWaitQueue_enq_bits_needRead, readWaitQueue_enq_bits_last};
  wire [10:0]       readWaitQueue_dataIn_hi_hi = {readWaitQueue_enq_bits_executeGroup, readWaitQueue_enq_bits_sourceValid};
  wire [14:0]       readWaitQueue_dataIn_hi = {readWaitQueue_dataIn_hi_hi, readWaitQueue_enq_bits_replaceVs1};
  wire [19:0]       readWaitQueue_dataIn = {readWaitQueue_dataIn_hi, readWaitQueue_dataIn_lo};
  assign readWaitQueue_dataOut_last = _readWaitQueue_fifo_data_out[0];
  assign readWaitQueue_dataOut_needRead = _readWaitQueue_fifo_data_out[4:1];
  assign readWaitQueue_dataOut_replaceVs1 = _readWaitQueue_fifo_data_out[8:5];
  assign readWaitQueue_dataOut_sourceValid = _readWaitQueue_fifo_data_out[12:9];
  assign readWaitQueue_dataOut_executeGroup = _readWaitQueue_fifo_data_out[19:13];
  wire [6:0]        readWaitQueue_deq_bits_executeGroup = readWaitQueue_dataOut_executeGroup;
  wire [3:0]        readWaitQueue_deq_bits_sourceValid = readWaitQueue_dataOut_sourceValid;
  wire [3:0]        readWaitQueue_deq_bits_replaceVs1 = readWaitQueue_dataOut_replaceVs1;
  wire [3:0]        readWaitQueue_deq_bits_needRead = readWaitQueue_dataOut_needRead;
  wire              readWaitQueue_deq_bits_last = readWaitQueue_dataOut_last;
  wire              readWaitQueue_enq_ready = ~_readWaitQueue_fifo_full;
  wire              readWaitQueue_enq_valid;
  wire              readWaitQueue_deq_ready;
  wire              _GEN_36 = lastExecuteGroupDeq | viota;
  assign exeRequestQueue_0_deq_ready = ~exeReqReg_0_valid | _GEN_36;
  assign exeRequestQueue_1_deq_ready = ~exeReqReg_1_valid | _GEN_36;
  assign exeRequestQueue_2_deq_ready = ~exeReqReg_2_valid | _GEN_36;
  assign exeRequestQueue_3_deq_ready = ~exeReqReg_3_valid | _GEN_36;
  wire              isLastExecuteGroup = executeIndex == lastExecuteIndex;
  wire              allDataValid = (exeReqReg_0_valid | ~(groupDataNeed[0])) & (exeReqReg_1_valid | ~(groupDataNeed[1])) & (exeReqReg_2_valid | ~(groupDataNeed[2])) & (exeReqReg_3_valid | ~(groupDataNeed[3]));
  wire              anyDataValid = exeReqReg_0_valid | exeReqReg_1_valid | exeReqReg_2_valid | exeReqReg_3_valid;
  wire              _GEN_37 = compress | mvRd;
  wire              readVs1Valid = (unitType[2] | _GEN_37) & ~readVS1Reg_requestSend | gatherSRead;
  wire [4:0]        readVS1Req_vs = compress ? instReg_vs1 + {4'h0, readVS1Reg_readIndex[3]} : gatherSRead ? instReg_vs1 + {2'h0, gatherGrowth} : instReg_vs1;
  wire              readVS1Req_offset = compress ? readVS1Reg_readIndex[2] : gatherSRead & gatherOffset;
  wire [1:0]        readVS1Req_readLane = compress ? readVS1Reg_readIndex[1:0] : gatherSRead ? gatherLane : 2'h0;
  wire [1:0]        readVS1Req_dataOffset = compress | ~gatherSRead ? 2'h0 : gatherDatOffset;
  wire              selectExecuteReq_1_bits_offset = readIssueStageState_readOffset[1];
  wire              selectExecuteReq_2_bits_offset = readIssueStageState_readOffset[2];
  wire              selectExecuteReq_3_bits_offset = readIssueStageState_readOffset[3];
  wire [1:0]        selectExecuteReq_1_bits_dataOffset = readIssueStageState_readDataOffset[3:2];
  wire [1:0]        selectExecuteReq_2_bits_dataOffset = readIssueStageState_readDataOffset[5:4];
  wire [1:0]        selectExecuteReq_3_bits_dataOffset = readIssueStageState_readDataOffset[7:6];
  wire              selectExecuteReq_0_valid = readVs1Valid | readIssueStageValid & ~(readIssueStageState_groupReadState[0]) & readIssueStageState_needRead[0] & readType;
  wire [4:0]        selectExecuteReq_0_bits_vs = readVs1Valid ? readVS1Req_vs : instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_0};
  wire              selectExecuteReq_0_bits_offset = readVs1Valid ? readVS1Req_offset : readIssueStageState_readOffset[0];
  wire [1:0]        selectExecuteReq_0_bits_readLane = readVs1Valid ? readVS1Req_readLane : readIssueStageState_accessLane_0;
  wire [1:0]        selectExecuteReq_0_bits_dataOffset = readVs1Valid ? readVS1Req_dataOffset : readIssueStageState_readDataOffset[1:0];
  wire              _tokenCheck_T = _readCrossBar_input_0_ready & readCrossBar_input_0_valid;
  wire              pipeReadFire_0 = ~readVs1Valid & _tokenCheck_T;
  wire [4:0]        selectExecuteReq_1_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_1};
  wire              selectExecuteReq_1_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[1]) & readIssueStageState_needRead[1] & readType;
  wire              pipeReadFire_1 = _readCrossBar_input_1_ready & readCrossBar_input_1_valid;
  wire [4:0]        selectExecuteReq_2_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_2};
  wire              selectExecuteReq_2_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[2]) & readIssueStageState_needRead[2] & readType;
  wire              pipeReadFire_2 = _readCrossBar_input_2_ready & readCrossBar_input_2_valid;
  wire [4:0]        selectExecuteReq_3_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_3};
  wire              selectExecuteReq_3_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[3]) & readIssueStageState_needRead[3] & readType;
  wire              pipeReadFire_3 = _readCrossBar_input_3_ready & readCrossBar_input_3_valid;
  reg  [3:0]        tokenCheck_counter;
  wire [3:0]        tokenCheck_counterChange = _tokenCheck_T ? 4'h1 : 4'hF;
  wire              tokenCheck = ~(tokenCheck_counter[3]);
  assign readCrossBar_input_0_valid = selectExecuteReq_0_valid & tokenCheck;
  reg  [3:0]        tokenCheck_counter_1;
  wire [3:0]        tokenCheck_counterChange_1 = pipeReadFire_1 ? 4'h1 : 4'hF;
  wire              tokenCheck_1 = ~(tokenCheck_counter_1[3]);
  assign readCrossBar_input_1_valid = selectExecuteReq_1_valid & tokenCheck_1;
  reg  [3:0]        tokenCheck_counter_2;
  wire [3:0]        tokenCheck_counterChange_2 = pipeReadFire_2 ? 4'h1 : 4'hF;
  wire              tokenCheck_2 = ~(tokenCheck_counter_2[3]);
  assign readCrossBar_input_2_valid = selectExecuteReq_2_valid & tokenCheck_2;
  reg  [3:0]        tokenCheck_counter_3;
  wire [3:0]        tokenCheck_counterChange_3 = pipeReadFire_3 ? 4'h1 : 4'hF;
  wire              tokenCheck_3 = ~(tokenCheck_counter_3[3]);
  assign readCrossBar_input_3_valid = selectExecuteReq_3_valid & tokenCheck_3;
  wire [1:0]        readFire_lo = {pipeReadFire_1, pipeReadFire_0};
  wire [1:0]        readFire_hi = {pipeReadFire_3, pipeReadFire_2};
  wire [3:0]        readFire = {readFire_hi, readFire_lo};
  wire              anyReadFire = |readFire;
  wire [3:0]        readStateUpdate = readFire | readIssueStageState_groupReadState;
  wire              groupReadFinish = readStateUpdate == readIssueStageState_needRead;
  assign readTypeRequestDeq = anyReadFire & groupReadFinish | readIssueStageValid & readIssueStageState_needRead == 4'h0;
  assign readWaitQueue_enq_valid = readTypeRequestDeq;
  wire [3:0]        compressUnitResultQueue_enq_bits_ffoOutput;
  wire              compressUnitResultQueue_enq_bits_compressValid;
  wire [4:0]        compressUnitResultQueue_dataIn_lo = {compressUnitResultQueue_enq_bits_ffoOutput, compressUnitResultQueue_enq_bits_compressValid};
  wire [127:0]      compressUnitResultQueue_enq_bits_data;
  wire [15:0]       compressUnitResultQueue_enq_bits_mask;
  wire [143:0]      compressUnitResultQueue_dataIn_hi_hi = {compressUnitResultQueue_enq_bits_data, compressUnitResultQueue_enq_bits_mask};
  wire [4:0]        compressUnitResultQueue_enq_bits_groupCounter;
  wire [148:0]      compressUnitResultQueue_dataIn_hi = {compressUnitResultQueue_dataIn_hi_hi, compressUnitResultQueue_enq_bits_groupCounter};
  wire [153:0]      compressUnitResultQueue_dataIn = {compressUnitResultQueue_dataIn_hi, compressUnitResultQueue_dataIn_lo};
  wire              compressUnitResultQueue_dataOut_compressValid = _compressUnitResultQueue_fifo_data_out[0];
  wire [3:0]        compressUnitResultQueue_dataOut_ffoOutput = _compressUnitResultQueue_fifo_data_out[4:1];
  wire [4:0]        compressUnitResultQueue_dataOut_groupCounter = _compressUnitResultQueue_fifo_data_out[9:5];
  wire [15:0]       compressUnitResultQueue_dataOut_mask = _compressUnitResultQueue_fifo_data_out[25:10];
  wire [127:0]      compressUnitResultQueue_dataOut_data = _compressUnitResultQueue_fifo_data_out[153:26];
  wire              compressUnitResultQueue_enq_ready = ~_compressUnitResultQueue_fifo_full;
  wire              compressUnitResultQueue_deq_ready;
  wire              compressUnitResultQueue_enq_valid;
  wire              compressUnitResultQueue_deq_valid = ~_compressUnitResultQueue_fifo_empty | compressUnitResultQueue_enq_valid;
  wire [127:0]      compressUnitResultQueue_deq_bits_data = _compressUnitResultQueue_fifo_empty ? compressUnitResultQueue_enq_bits_data : compressUnitResultQueue_dataOut_data;
  wire [15:0]       compressUnitResultQueue_deq_bits_mask = _compressUnitResultQueue_fifo_empty ? compressUnitResultQueue_enq_bits_mask : compressUnitResultQueue_dataOut_mask;
  wire [4:0]        compressUnitResultQueue_deq_bits_groupCounter = _compressUnitResultQueue_fifo_empty ? compressUnitResultQueue_enq_bits_groupCounter : compressUnitResultQueue_dataOut_groupCounter;
  wire [3:0]        compressUnitResultQueue_deq_bits_ffoOutput = _compressUnitResultQueue_fifo_empty ? compressUnitResultQueue_enq_bits_ffoOutput : compressUnitResultQueue_dataOut_ffoOutput;
  wire              compressUnitResultQueue_deq_bits_compressValid = _compressUnitResultQueue_fifo_empty ? compressUnitResultQueue_enq_bits_compressValid : compressUnitResultQueue_dataOut_compressValid;
  wire              noSourceValid = noSource & counterValid & ((|instReg_vl) | mvRd & ~readVS1Reg_sendToExecution);
  wire              vs1DataValid = readVS1Reg_dataValid | ~(unitType[2] | _GEN_37);
  wire [1:0]        _GEN_38 = {_maskedWrite_in_1_ready, _maskedWrite_in_0_ready};
  wire [1:0]        executeDeqReady_lo;
  assign executeDeqReady_lo = _GEN_38;
  wire [1:0]        compressUnitResultQueue_deq_ready_lo;
  assign compressUnitResultQueue_deq_ready_lo = _GEN_38;
  wire [1:0]        _GEN_39 = {_maskedWrite_in_3_ready, _maskedWrite_in_2_ready};
  wire [1:0]        executeDeqReady_hi;
  assign executeDeqReady_hi = _GEN_39;
  wire [1:0]        compressUnitResultQueue_deq_ready_hi;
  assign compressUnitResultQueue_deq_ready_hi = _GEN_39;
  wire              compressUnitResultQueue_empty;
  wire              executeDeqReady = (&{executeDeqReady_hi, executeDeqReady_lo}) & compressUnitResultQueue_empty;
  wire              otherTypeRequestDeq = (noSource ? noSourceValid : allDataValid) & vs1DataValid & instVlValid & executeDeqReady;
  wire              reorderQueueAllocate;
  wire              _GEN_40 = accessCountQueue_enq_ready & reorderQueueAllocate;
  assign readIssueStageEnq = (allDataValid | _slideAddressGen_indexDeq_valid) & (readTypeRequestDeq | ~readIssueStageValid) & instVlValid & readType & _GEN_40;
  assign accessCountQueue_enq_valid = readIssueStageEnq;
  wire              executeReady;
  wire              requestStageDeq = readType ? readIssueStageEnq : otherTypeRequestDeq & executeReady;
  wire              slideAddressGen_indexDeq_ready = (readTypeRequestDeq | ~readIssueStageValid) & _GEN_40;
  wire              _GEN_41 = slideAddressGen_indexDeq_ready & _slideAddressGen_indexDeq_valid;
  wire              _GEN_42 = readIssueStageEnq & _GEN_41;
  assign accessCountEnq_0 =
    _GEN_42
      ? {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 2'h0 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 2'h0 & _slideAddressGen_indexDeq_bits_needRead[1]}}
        + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 2'h0 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 2'h0 & _slideAddressGen_indexDeq_bits_needRead[3]}}
      : {1'h0, {1'h0, accessLaneSelect[1:0] == 2'h0 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[3:2] == 2'h0 & ~(notReadSelect[1])}}
        + {1'h0, {1'h0, accessLaneSelect[5:4] == 2'h0 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[7:6] == 2'h0 & ~(notReadSelect[3])}};
  assign accessCountEnq_1 =
    _GEN_42
      ? {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 2'h1 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 2'h1 & _slideAddressGen_indexDeq_bits_needRead[1]}}
        + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 2'h1 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 2'h1 & _slideAddressGen_indexDeq_bits_needRead[3]}}
      : {1'h0, {1'h0, accessLaneSelect[1:0] == 2'h1 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[3:2] == 2'h1 & ~(notReadSelect[1])}}
        + {1'h0, {1'h0, accessLaneSelect[5:4] == 2'h1 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[7:6] == 2'h1 & ~(notReadSelect[3])}};
  assign accessCountEnq_2 =
    _GEN_42
      ? {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 2'h2 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 2'h2 & _slideAddressGen_indexDeq_bits_needRead[1]}}
        + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 2'h2 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 2'h2 & _slideAddressGen_indexDeq_bits_needRead[3]}}
      : {1'h0, {1'h0, accessLaneSelect[1:0] == 2'h2 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[3:2] == 2'h2 & ~(notReadSelect[1])}}
        + {1'h0, {1'h0, accessLaneSelect[5:4] == 2'h2 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[7:6] == 2'h2 & ~(notReadSelect[3])}};
  assign accessCountEnq_3 =
    _GEN_42
      ? {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_0) & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_1) & _slideAddressGen_indexDeq_bits_needRead[1]}}
        + {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_2) & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_3) & _slideAddressGen_indexDeq_bits_needRead[3]}}
      : {1'h0, {1'h0, (&(accessLaneSelect[1:0])) & ~(notReadSelect[0])} + {1'h0, (&(accessLaneSelect[3:2])) & ~(notReadSelect[1])}}
        + {1'h0, {1'h0, (&(accessLaneSelect[5:4])) & ~(notReadSelect[2])} + {1'h0, (&(accessLaneSelect[7:6])) & ~(notReadSelect[3])}};
  assign lastExecuteGroupDeq = requestStageDeq & isLastExecuteGroup;
  wire [3:0]        readMessageQueue_deq_bits_readSource;
  wire              deqAllocate;
  wire              reorderQueueVec_0_deq_valid;
  assign reorderQueueVec_0_deq_valid = ~_reorderQueueVec_fifo_empty;
  wire [31:0]       reorderQueueVec_dataOut_data;
  wire [3:0]        reorderQueueVec_dataOut_write1H;
  wire [31:0]       dataAfterReorderCheck_0 = reorderQueueVec_0_deq_bits_data;
  wire [31:0]       reorderQueueVec_0_enq_bits_data;
  wire [3:0]        reorderQueueVec_0_enq_bits_write1H;
  wire [35:0]       reorderQueueVec_dataIn = {reorderQueueVec_0_enq_bits_data, reorderQueueVec_0_enq_bits_write1H};
  assign reorderQueueVec_dataOut_write1H = _reorderQueueVec_fifo_data_out[3:0];
  assign reorderQueueVec_dataOut_data = _reorderQueueVec_fifo_data_out[35:4];
  assign reorderQueueVec_0_deq_bits_data = reorderQueueVec_dataOut_data;
  wire [3:0]        reorderQueueVec_0_deq_bits_write1H = reorderQueueVec_dataOut_write1H;
  wire              reorderQueueVec_0_enq_ready = ~_reorderQueueVec_fifo_full;
  wire              reorderQueueVec_0_deq_ready;
  wire [3:0]        readMessageQueue_1_deq_bits_readSource;
  wire              deqAllocate_1;
  wire              reorderQueueVec_1_deq_valid;
  assign reorderQueueVec_1_deq_valid = ~_reorderQueueVec_fifo_1_empty;
  wire [31:0]       reorderQueueVec_dataOut_1_data;
  wire [3:0]        reorderQueueVec_dataOut_1_write1H;
  wire [31:0]       dataAfterReorderCheck_1 = reorderQueueVec_1_deq_bits_data;
  wire [31:0]       reorderQueueVec_1_enq_bits_data;
  wire [3:0]        reorderQueueVec_1_enq_bits_write1H;
  wire [35:0]       reorderQueueVec_dataIn_1 = {reorderQueueVec_1_enq_bits_data, reorderQueueVec_1_enq_bits_write1H};
  assign reorderQueueVec_dataOut_1_write1H = _reorderQueueVec_fifo_1_data_out[3:0];
  assign reorderQueueVec_dataOut_1_data = _reorderQueueVec_fifo_1_data_out[35:4];
  assign reorderQueueVec_1_deq_bits_data = reorderQueueVec_dataOut_1_data;
  wire [3:0]        reorderQueueVec_1_deq_bits_write1H = reorderQueueVec_dataOut_1_write1H;
  wire              reorderQueueVec_1_enq_ready = ~_reorderQueueVec_fifo_1_full;
  wire              reorderQueueVec_1_deq_ready;
  wire [3:0]        readMessageQueue_2_deq_bits_readSource;
  wire              deqAllocate_2;
  wire              reorderQueueVec_2_deq_valid;
  assign reorderQueueVec_2_deq_valid = ~_reorderQueueVec_fifo_2_empty;
  wire [31:0]       reorderQueueVec_dataOut_2_data;
  wire [3:0]        reorderQueueVec_dataOut_2_write1H;
  wire [31:0]       dataAfterReorderCheck_2 = reorderQueueVec_2_deq_bits_data;
  wire [31:0]       reorderQueueVec_2_enq_bits_data;
  wire [3:0]        reorderQueueVec_2_enq_bits_write1H;
  wire [35:0]       reorderQueueVec_dataIn_2 = {reorderQueueVec_2_enq_bits_data, reorderQueueVec_2_enq_bits_write1H};
  assign reorderQueueVec_dataOut_2_write1H = _reorderQueueVec_fifo_2_data_out[3:0];
  assign reorderQueueVec_dataOut_2_data = _reorderQueueVec_fifo_2_data_out[35:4];
  assign reorderQueueVec_2_deq_bits_data = reorderQueueVec_dataOut_2_data;
  wire [3:0]        reorderQueueVec_2_deq_bits_write1H = reorderQueueVec_dataOut_2_write1H;
  wire              reorderQueueVec_2_enq_ready = ~_reorderQueueVec_fifo_2_full;
  wire              reorderQueueVec_2_deq_ready;
  wire [3:0]        readMessageQueue_3_deq_bits_readSource;
  wire              deqAllocate_3;
  wire              reorderQueueVec_3_deq_valid;
  assign reorderQueueVec_3_deq_valid = ~_reorderQueueVec_fifo_3_empty;
  wire [31:0]       reorderQueueVec_dataOut_3_data;
  wire [3:0]        reorderQueueVec_dataOut_3_write1H;
  wire [31:0]       dataAfterReorderCheck_3 = reorderQueueVec_3_deq_bits_data;
  wire [31:0]       reorderQueueVec_3_enq_bits_data;
  wire [3:0]        reorderQueueVec_3_enq_bits_write1H;
  wire [35:0]       reorderQueueVec_dataIn_3 = {reorderQueueVec_3_enq_bits_data, reorderQueueVec_3_enq_bits_write1H};
  assign reorderQueueVec_dataOut_3_write1H = _reorderQueueVec_fifo_3_data_out[3:0];
  assign reorderQueueVec_dataOut_3_data = _reorderQueueVec_fifo_3_data_out[35:4];
  assign reorderQueueVec_3_deq_bits_data = reorderQueueVec_dataOut_3_data;
  wire [3:0]        reorderQueueVec_3_deq_bits_write1H = reorderQueueVec_dataOut_3_write1H;
  wire              reorderQueueVec_3_enq_ready = ~_reorderQueueVec_fifo_3_full;
  wire              reorderQueueVec_3_deq_ready;
  reg  [3:0]        reorderQueueAllocate_counter;
  reg  [3:0]        reorderQueueAllocate_counterWillUpdate;
  wire              _write1HPipe_0_T = reorderQueueVec_0_deq_ready & reorderQueueVec_0_deq_valid;
  wire              reorderQueueAllocate_release = _write1HPipe_0_T & readValid;
  wire [2:0]        reorderQueueAllocate_allocate = readIssueStageEnq ? accessCountEnq_0 : 3'h0;
  wire [3:0]        reorderQueueAllocate_counterUpdate = reorderQueueAllocate_counter + {1'h0, reorderQueueAllocate_allocate} - {3'h0, reorderQueueAllocate_release};
  reg  [3:0]        reorderQueueAllocate_counter_1;
  reg  [3:0]        reorderQueueAllocate_counterWillUpdate_1;
  wire              _write1HPipe_1_T = reorderQueueVec_1_deq_ready & reorderQueueVec_1_deq_valid;
  wire              reorderQueueAllocate_release_1 = _write1HPipe_1_T & readValid;
  wire [2:0]        reorderQueueAllocate_allocate_1 = readIssueStageEnq ? accessCountEnq_1 : 3'h0;
  wire [3:0]        reorderQueueAllocate_counterUpdate_1 = reorderQueueAllocate_counter_1 + {1'h0, reorderQueueAllocate_allocate_1} - {3'h0, reorderQueueAllocate_release_1};
  reg  [3:0]        reorderQueueAllocate_counter_2;
  reg  [3:0]        reorderQueueAllocate_counterWillUpdate_2;
  wire              _write1HPipe_2_T = reorderQueueVec_2_deq_ready & reorderQueueVec_2_deq_valid;
  wire              reorderQueueAllocate_release_2 = _write1HPipe_2_T & readValid;
  wire [2:0]        reorderQueueAllocate_allocate_2 = readIssueStageEnq ? accessCountEnq_2 : 3'h0;
  wire [3:0]        reorderQueueAllocate_counterUpdate_2 = reorderQueueAllocate_counter_2 + {1'h0, reorderQueueAllocate_allocate_2} - {3'h0, reorderQueueAllocate_release_2};
  reg  [3:0]        reorderQueueAllocate_counter_3;
  reg  [3:0]        reorderQueueAllocate_counterWillUpdate_3;
  wire              _write1HPipe_3_T = reorderQueueVec_3_deq_ready & reorderQueueVec_3_deq_valid;
  wire              reorderQueueAllocate_release_3 = _write1HPipe_3_T & readValid;
  wire [2:0]        reorderQueueAllocate_allocate_3 = readIssueStageEnq ? accessCountEnq_3 : 3'h0;
  wire [3:0]        reorderQueueAllocate_counterUpdate_3 = reorderQueueAllocate_counter_3 + {1'h0, reorderQueueAllocate_allocate_3} - {3'h0, reorderQueueAllocate_release_3};
  assign reorderQueueAllocate = ~(reorderQueueAllocate_counterWillUpdate[3]) & ~(reorderQueueAllocate_counterWillUpdate_1[3]) & ~(reorderQueueAllocate_counterWillUpdate_2[3]) & ~(reorderQueueAllocate_counterWillUpdate_3[3]);
  reg               reorderStageValid;
  reg  [2:0]        reorderStageState_0;
  reg  [2:0]        reorderStageState_1;
  reg  [2:0]        reorderStageState_2;
  reg  [2:0]        reorderStageState_3;
  reg  [2:0]        reorderStageNeed_0;
  reg  [2:0]        reorderStageNeed_1;
  reg  [2:0]        reorderStageNeed_2;
  reg  [2:0]        reorderStageNeed_3;
  wire              stateCheck = reorderStageState_0 == reorderStageNeed_0 & reorderStageState_1 == reorderStageNeed_1 & reorderStageState_2 == reorderStageNeed_2 & reorderStageState_3 == reorderStageNeed_3;
  assign accessCountQueue_deq_ready = ~reorderStageValid | stateCheck;
  wire              reorderStageEnqFire = accessCountQueue_deq_ready & accessCountQueue_deq_valid;
  wire              reorderStageDeqFire = stateCheck & reorderStageValid;
  wire [3:0]        sourceLane;
  wire              readMessageQueue_deq_valid;
  assign readMessageQueue_deq_valid = ~_readMessageQueue_fifo_empty;
  wire [3:0]        readMessageQueue_dataOut_readSource;
  assign reorderQueueVec_0_enq_bits_write1H = readMessageQueue_deq_bits_readSource;
  wire [1:0]        readMessageQueue_dataOut_dataOffset;
  wire [3:0]        readMessageQueue_enq_bits_readSource;
  wire [1:0]        readMessageQueue_enq_bits_dataOffset;
  wire [5:0]        readMessageQueue_dataIn = {readMessageQueue_enq_bits_readSource, readMessageQueue_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_dataOffset = _readMessageQueue_fifo_data_out[1:0];
  assign readMessageQueue_dataOut_readSource = _readMessageQueue_fifo_data_out[5:2];
  assign readMessageQueue_deq_bits_readSource = readMessageQueue_dataOut_readSource;
  wire [1:0]        readMessageQueue_deq_bits_dataOffset = readMessageQueue_dataOut_dataOffset;
  wire              readMessageQueue_enq_ready = ~_readMessageQueue_fifo_full;
  wire              readMessageQueue_enq_valid;
  assign deqAllocate = ~readValid | reorderStageValid & reorderStageState_0 != reorderStageNeed_0;
  assign reorderQueueVec_0_deq_ready = deqAllocate;
  assign sourceLane = 4'h1 << _readCrossBar_output_0_bits_writeIndex;
  assign readMessageQueue_enq_bits_readSource = sourceLane;
  wire              readChannel_0_valid_0 = maskDestinationType ? _maskedWrite_readChannel_0_valid : _readCrossBar_output_0_valid & readMessageQueue_enq_ready;
  wire [4:0]        readChannel_0_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_0_bits_vs : _readCrossBar_output_0_bits_vs;
  wire              readChannel_0_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_0_bits_offset : _readCrossBar_output_0_bits_offset;
  assign readMessageQueue_enq_valid = readChannel_0_ready_0 & readChannel_0_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_0_enq_bits_data = readResult_0_bits >> {27'h0, readMessageQueue_deq_bits_dataOffset, 3'h0};
  wire [3:0]        write1HPipe_0 = _write1HPipe_0_T & ~maskDestinationType ? reorderQueueVec_0_deq_bits_write1H : 4'h0;
  wire [3:0]        sourceLane_1;
  wire              readMessageQueue_1_deq_valid;
  assign readMessageQueue_1_deq_valid = ~_readMessageQueue_fifo_1_empty;
  wire [3:0]        readMessageQueue_dataOut_1_readSource;
  assign reorderQueueVec_1_enq_bits_write1H = readMessageQueue_1_deq_bits_readSource;
  wire [1:0]        readMessageQueue_dataOut_1_dataOffset;
  wire [3:0]        readMessageQueue_1_enq_bits_readSource;
  wire [1:0]        readMessageQueue_1_enq_bits_dataOffset;
  wire [5:0]        readMessageQueue_dataIn_1 = {readMessageQueue_1_enq_bits_readSource, readMessageQueue_1_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_1_dataOffset = _readMessageQueue_fifo_1_data_out[1:0];
  assign readMessageQueue_dataOut_1_readSource = _readMessageQueue_fifo_1_data_out[5:2];
  assign readMessageQueue_1_deq_bits_readSource = readMessageQueue_dataOut_1_readSource;
  wire [1:0]        readMessageQueue_1_deq_bits_dataOffset = readMessageQueue_dataOut_1_dataOffset;
  wire              readMessageQueue_1_enq_ready = ~_readMessageQueue_fifo_1_full;
  wire              readMessageQueue_1_enq_valid;
  assign deqAllocate_1 = ~readValid | reorderStageValid & reorderStageState_1 != reorderStageNeed_1;
  assign reorderQueueVec_1_deq_ready = deqAllocate_1;
  assign sourceLane_1 = 4'h1 << _readCrossBar_output_1_bits_writeIndex;
  assign readMessageQueue_1_enq_bits_readSource = sourceLane_1;
  wire              readChannel_1_valid_0 = maskDestinationType ? _maskedWrite_readChannel_1_valid : _readCrossBar_output_1_valid & readMessageQueue_1_enq_ready;
  wire [4:0]        readChannel_1_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_1_bits_vs : _readCrossBar_output_1_bits_vs;
  wire              readChannel_1_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_1_bits_offset : _readCrossBar_output_1_bits_offset;
  assign readMessageQueue_1_enq_valid = readChannel_1_ready_0 & readChannel_1_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_1_enq_bits_data = readResult_1_bits >> {27'h0, readMessageQueue_1_deq_bits_dataOffset, 3'h0};
  wire [3:0]        write1HPipe_1 = _write1HPipe_1_T & ~maskDestinationType ? reorderQueueVec_1_deq_bits_write1H : 4'h0;
  wire [3:0]        sourceLane_2;
  wire              readMessageQueue_2_deq_valid;
  assign readMessageQueue_2_deq_valid = ~_readMessageQueue_fifo_2_empty;
  wire [3:0]        readMessageQueue_dataOut_2_readSource;
  assign reorderQueueVec_2_enq_bits_write1H = readMessageQueue_2_deq_bits_readSource;
  wire [1:0]        readMessageQueue_dataOut_2_dataOffset;
  wire [3:0]        readMessageQueue_2_enq_bits_readSource;
  wire [1:0]        readMessageQueue_2_enq_bits_dataOffset;
  wire [5:0]        readMessageQueue_dataIn_2 = {readMessageQueue_2_enq_bits_readSource, readMessageQueue_2_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_2_dataOffset = _readMessageQueue_fifo_2_data_out[1:0];
  assign readMessageQueue_dataOut_2_readSource = _readMessageQueue_fifo_2_data_out[5:2];
  assign readMessageQueue_2_deq_bits_readSource = readMessageQueue_dataOut_2_readSource;
  wire [1:0]        readMessageQueue_2_deq_bits_dataOffset = readMessageQueue_dataOut_2_dataOffset;
  wire              readMessageQueue_2_enq_ready = ~_readMessageQueue_fifo_2_full;
  wire              readMessageQueue_2_enq_valid;
  assign deqAllocate_2 = ~readValid | reorderStageValid & reorderStageState_2 != reorderStageNeed_2;
  assign reorderQueueVec_2_deq_ready = deqAllocate_2;
  assign sourceLane_2 = 4'h1 << _readCrossBar_output_2_bits_writeIndex;
  assign readMessageQueue_2_enq_bits_readSource = sourceLane_2;
  wire              readChannel_2_valid_0 = maskDestinationType ? _maskedWrite_readChannel_2_valid : _readCrossBar_output_2_valid & readMessageQueue_2_enq_ready;
  wire [4:0]        readChannel_2_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_2_bits_vs : _readCrossBar_output_2_bits_vs;
  wire              readChannel_2_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_2_bits_offset : _readCrossBar_output_2_bits_offset;
  assign readMessageQueue_2_enq_valid = readChannel_2_ready_0 & readChannel_2_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_2_enq_bits_data = readResult_2_bits >> {27'h0, readMessageQueue_2_deq_bits_dataOffset, 3'h0};
  wire [3:0]        write1HPipe_2 = _write1HPipe_2_T & ~maskDestinationType ? reorderQueueVec_2_deq_bits_write1H : 4'h0;
  wire [3:0]        sourceLane_3;
  wire              readMessageQueue_3_deq_valid;
  assign readMessageQueue_3_deq_valid = ~_readMessageQueue_fifo_3_empty;
  wire [3:0]        readMessageQueue_dataOut_3_readSource;
  assign reorderQueueVec_3_enq_bits_write1H = readMessageQueue_3_deq_bits_readSource;
  wire [1:0]        readMessageQueue_dataOut_3_dataOffset;
  wire [3:0]        readMessageQueue_3_enq_bits_readSource;
  wire [1:0]        readMessageQueue_3_enq_bits_dataOffset;
  wire [5:0]        readMessageQueue_dataIn_3 = {readMessageQueue_3_enq_bits_readSource, readMessageQueue_3_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_3_dataOffset = _readMessageQueue_fifo_3_data_out[1:0];
  assign readMessageQueue_dataOut_3_readSource = _readMessageQueue_fifo_3_data_out[5:2];
  assign readMessageQueue_3_deq_bits_readSource = readMessageQueue_dataOut_3_readSource;
  wire [1:0]        readMessageQueue_3_deq_bits_dataOffset = readMessageQueue_dataOut_3_dataOffset;
  wire              readMessageQueue_3_enq_ready = ~_readMessageQueue_fifo_3_full;
  wire              readMessageQueue_3_enq_valid;
  assign deqAllocate_3 = ~readValid | reorderStageValid & reorderStageState_3 != reorderStageNeed_3;
  assign reorderQueueVec_3_deq_ready = deqAllocate_3;
  assign sourceLane_3 = 4'h1 << _readCrossBar_output_3_bits_writeIndex;
  assign readMessageQueue_3_enq_bits_readSource = sourceLane_3;
  wire              readChannel_3_valid_0 = maskDestinationType ? _maskedWrite_readChannel_3_valid : _readCrossBar_output_3_valid & readMessageQueue_3_enq_ready;
  wire [4:0]        readChannel_3_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_3_bits_vs : _readCrossBar_output_3_bits_vs;
  wire              readChannel_3_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_3_bits_offset : _readCrossBar_output_3_bits_offset;
  assign readMessageQueue_3_enq_valid = readChannel_3_ready_0 & readChannel_3_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_3_enq_bits_data = readResult_3_bits >> {27'h0, readMessageQueue_3_deq_bits_dataOffset, 3'h0};
  wire [3:0]        write1HPipe_3 = _write1HPipe_3_T & ~maskDestinationType ? reorderQueueVec_3_deq_bits_write1H : 4'h0;
  wire [31:0]       readData_data;
  wire              readData_readDataQueue_enq_ready = ~_readData_readDataQueue_fifo_full;
  wire              readData_readDataQueue_deq_ready;
  wire              readData_readDataQueue_enq_valid;
  wire              readData_readDataQueue_deq_valid = ~_readData_readDataQueue_fifo_empty | readData_readDataQueue_enq_valid;
  wire [31:0]       readData_readDataQueue_enq_bits;
  wire [31:0]       readData_readDataQueue_deq_bits = _readData_readDataQueue_fifo_empty ? readData_readDataQueue_enq_bits : _readData_readDataQueue_fifo_data_out;
  wire [1:0]        readData_readResultSelect_lo = {write1HPipe_1[0], write1HPipe_0[0]};
  wire [1:0]        readData_readResultSelect_hi = {write1HPipe_3[0], write1HPipe_2[0]};
  wire [3:0]        readData_readResultSelect = {readData_readResultSelect_hi, readData_readResultSelect_lo};
  assign readData_data =
    (readData_readResultSelect[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect[3] ? dataAfterReorderCheck_3 : 32'h0);
  assign readData_readDataQueue_enq_bits = readData_data;
  wire              readTokenRelease_0 = readData_readDataQueue_deq_ready & readData_readDataQueue_deq_valid;
  assign readData_readDataQueue_enq_valid = |readData_readResultSelect;
  wire [31:0]       readData_data_1;
  wire              isWaiteForThisData_1;
  wire              readData_readDataQueue_1_enq_ready = ~_readData_readDataQueue_fifo_1_full;
  wire              readData_readDataQueue_1_deq_ready;
  wire              readData_readDataQueue_1_enq_valid;
  wire              readData_readDataQueue_1_deq_valid = ~_readData_readDataQueue_fifo_1_empty | readData_readDataQueue_1_enq_valid;
  wire [31:0]       readData_readDataQueue_1_enq_bits;
  wire [31:0]       readData_readDataQueue_1_deq_bits = _readData_readDataQueue_fifo_1_empty ? readData_readDataQueue_1_enq_bits : _readData_readDataQueue_fifo_1_data_out;
  wire [1:0]        readData_readResultSelect_lo_1 = {write1HPipe_1[1], write1HPipe_0[1]};
  wire [1:0]        readData_readResultSelect_hi_1 = {write1HPipe_3[1], write1HPipe_2[1]};
  wire [3:0]        readData_readResultSelect_1 = {readData_readResultSelect_hi_1, readData_readResultSelect_lo_1};
  assign readData_data_1 =
    (readData_readResultSelect_1[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_1[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_1[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_1[3] ? dataAfterReorderCheck_3 : 32'h0);
  assign readData_readDataQueue_1_enq_bits = readData_data_1;
  wire              readTokenRelease_1 = readData_readDataQueue_1_deq_ready & readData_readDataQueue_1_deq_valid;
  assign readData_readDataQueue_1_enq_valid = |readData_readResultSelect_1;
  wire [31:0]       readData_data_2;
  wire              isWaiteForThisData_2;
  wire              readData_readDataQueue_2_enq_ready = ~_readData_readDataQueue_fifo_2_full;
  wire              readData_readDataQueue_2_deq_ready;
  wire              readData_readDataQueue_2_enq_valid;
  wire              readData_readDataQueue_2_deq_valid = ~_readData_readDataQueue_fifo_2_empty | readData_readDataQueue_2_enq_valid;
  wire [31:0]       readData_readDataQueue_2_enq_bits;
  wire [31:0]       readData_readDataQueue_2_deq_bits = _readData_readDataQueue_fifo_2_empty ? readData_readDataQueue_2_enq_bits : _readData_readDataQueue_fifo_2_data_out;
  wire [1:0]        readData_readResultSelect_lo_2 = {write1HPipe_1[2], write1HPipe_0[2]};
  wire [1:0]        readData_readResultSelect_hi_2 = {write1HPipe_3[2], write1HPipe_2[2]};
  wire [3:0]        readData_readResultSelect_2 = {readData_readResultSelect_hi_2, readData_readResultSelect_lo_2};
  assign readData_data_2 =
    (readData_readResultSelect_2[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_2[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_2[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_2[3] ? dataAfterReorderCheck_3 : 32'h0);
  assign readData_readDataQueue_2_enq_bits = readData_data_2;
  wire              readTokenRelease_2 = readData_readDataQueue_2_deq_ready & readData_readDataQueue_2_deq_valid;
  assign readData_readDataQueue_2_enq_valid = |readData_readResultSelect_2;
  wire [31:0]       readData_data_3;
  wire              isWaiteForThisData_3;
  wire              readData_readDataQueue_3_enq_ready = ~_readData_readDataQueue_fifo_3_full;
  wire              readData_readDataQueue_3_deq_ready;
  wire              readData_readDataQueue_3_enq_valid;
  wire              readData_readDataQueue_3_deq_valid = ~_readData_readDataQueue_fifo_3_empty | readData_readDataQueue_3_enq_valid;
  wire [31:0]       readData_readDataQueue_3_enq_bits;
  wire [31:0]       readData_readDataQueue_3_deq_bits = _readData_readDataQueue_fifo_3_empty ? readData_readDataQueue_3_enq_bits : _readData_readDataQueue_fifo_3_data_out;
  wire [1:0]        readData_readResultSelect_lo_3 = {write1HPipe_1[3], write1HPipe_0[3]};
  wire [1:0]        readData_readResultSelect_hi_3 = {write1HPipe_3[3], write1HPipe_2[3]};
  wire [3:0]        readData_readResultSelect_3 = {readData_readResultSelect_hi_3, readData_readResultSelect_lo_3};
  assign readData_data_3 =
    (readData_readResultSelect_3[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_3[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_3[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_3[3] ? dataAfterReorderCheck_3 : 32'h0);
  assign readData_readDataQueue_3_enq_bits = readData_data_3;
  wire              readTokenRelease_3 = readData_readDataQueue_3_deq_ready & readData_readDataQueue_3_deq_valid;
  assign readData_readDataQueue_3_enq_valid = |readData_readResultSelect_3;
  reg  [6:0]        waiteReadDataPipeReg_executeGroup;
  reg  [3:0]        waiteReadDataPipeReg_sourceValid;
  reg  [3:0]        waiteReadDataPipeReg_replaceVs1;
  reg  [3:0]        waiteReadDataPipeReg_needRead;
  reg               waiteReadDataPipeReg_last;
  reg  [31:0]       waiteReadData_0;
  reg  [31:0]       waiteReadData_1;
  reg  [31:0]       waiteReadData_2;
  reg  [31:0]       waiteReadData_3;
  reg  [3:0]        waiteReadSate;
  reg               waiteReadStageValid;
  wire [1:0]        executeIndexVec_0 = waiteReadDataPipeReg_executeGroup[1:0];
  wire [1:0]        executeIndexVec_1 = {waiteReadDataPipeReg_executeGroup[0], 1'h0};
  wire              writeDataVec_data_dataIsRead = waiteReadDataPipeReg_needRead[0];
  wire              writeDataVec_data_dataIsRead_4 = waiteReadDataPipeReg_needRead[0];
  wire              writeDataVec_data_dataIsRead_8 = waiteReadDataPipeReg_needRead[0];
  wire [31:0]       _GEN_43 = waiteReadDataPipeReg_replaceVs1[0] ? instReg_readFromScala : 32'h0;
  wire [31:0]       writeDataVec_data_unreadData;
  assign writeDataVec_data_unreadData = _GEN_43;
  wire [31:0]       writeDataVec_data_unreadData_4;
  assign writeDataVec_data_unreadData_4 = _GEN_43;
  wire [31:0]       writeDataVec_data_unreadData_8;
  assign writeDataVec_data_unreadData_8 = _GEN_43;
  wire [7:0]        writeDataVec_data_dataElement = writeDataVec_data_dataIsRead ? waiteReadData_0[7:0] : writeDataVec_data_unreadData[7:0];
  wire              writeDataVec_data_dataIsRead_1 = waiteReadDataPipeReg_needRead[1];
  wire              writeDataVec_data_dataIsRead_5 = waiteReadDataPipeReg_needRead[1];
  wire              writeDataVec_data_dataIsRead_9 = waiteReadDataPipeReg_needRead[1];
  wire [31:0]       _GEN_44 = waiteReadDataPipeReg_replaceVs1[1] ? instReg_readFromScala : 32'h0;
  wire [31:0]       writeDataVec_data_unreadData_1;
  assign writeDataVec_data_unreadData_1 = _GEN_44;
  wire [31:0]       writeDataVec_data_unreadData_5;
  assign writeDataVec_data_unreadData_5 = _GEN_44;
  wire [31:0]       writeDataVec_data_unreadData_9;
  assign writeDataVec_data_unreadData_9 = _GEN_44;
  wire [7:0]        writeDataVec_data_dataElement_1 = writeDataVec_data_dataIsRead_1 ? waiteReadData_1[7:0] : writeDataVec_data_unreadData_1[7:0];
  wire              writeDataVec_data_dataIsRead_2 = waiteReadDataPipeReg_needRead[2];
  wire              writeDataVec_data_dataIsRead_6 = waiteReadDataPipeReg_needRead[2];
  wire              writeDataVec_data_dataIsRead_10 = waiteReadDataPipeReg_needRead[2];
  wire [31:0]       _GEN_45 = waiteReadDataPipeReg_replaceVs1[2] ? instReg_readFromScala : 32'h0;
  wire [31:0]       writeDataVec_data_unreadData_2;
  assign writeDataVec_data_unreadData_2 = _GEN_45;
  wire [31:0]       writeDataVec_data_unreadData_6;
  assign writeDataVec_data_unreadData_6 = _GEN_45;
  wire [31:0]       writeDataVec_data_unreadData_10;
  assign writeDataVec_data_unreadData_10 = _GEN_45;
  wire [7:0]        writeDataVec_data_dataElement_2 = writeDataVec_data_dataIsRead_2 ? waiteReadData_2[7:0] : writeDataVec_data_unreadData_2[7:0];
  wire              writeDataVec_data_dataIsRead_3 = waiteReadDataPipeReg_needRead[3];
  wire              writeDataVec_data_dataIsRead_7 = waiteReadDataPipeReg_needRead[3];
  wire              writeDataVec_data_dataIsRead_11 = waiteReadDataPipeReg_needRead[3];
  wire [31:0]       _GEN_46 = waiteReadDataPipeReg_replaceVs1[3] ? instReg_readFromScala : 32'h0;
  wire [31:0]       writeDataVec_data_unreadData_3;
  assign writeDataVec_data_unreadData_3 = _GEN_46;
  wire [31:0]       writeDataVec_data_unreadData_7;
  assign writeDataVec_data_unreadData_7 = _GEN_46;
  wire [31:0]       writeDataVec_data_unreadData_11;
  assign writeDataVec_data_unreadData_11 = _GEN_46;
  wire [7:0]        writeDataVec_data_dataElement_3 = writeDataVec_data_dataIsRead_3 ? waiteReadData_3[7:0] : writeDataVec_data_unreadData_3[7:0];
  wire [15:0]       writeDataVec_data_lo = {writeDataVec_data_dataElement_1, writeDataVec_data_dataElement};
  wire [15:0]       writeDataVec_data_hi = {writeDataVec_data_dataElement_3, writeDataVec_data_dataElement_2};
  wire [31:0]       writeDataVec_data = {writeDataVec_data_hi, writeDataVec_data_lo};
  wire [158:0]      writeDataVec_shifterData = {127'h0, writeDataVec_data} << {152'h0, executeIndexVec_0, 5'h0};
  wire [127:0]      writeDataVec_0 = writeDataVec_shifterData[127:0];
  wire [15:0]       writeDataVec_data_dataElement_4 = writeDataVec_data_dataIsRead_4 ? waiteReadData_0[15:0] : writeDataVec_data_unreadData_4[15:0];
  wire [15:0]       writeDataVec_data_dataElement_5 = writeDataVec_data_dataIsRead_5 ? waiteReadData_1[15:0] : writeDataVec_data_unreadData_5[15:0];
  wire [15:0]       writeDataVec_data_dataElement_6 = writeDataVec_data_dataIsRead_6 ? waiteReadData_2[15:0] : writeDataVec_data_unreadData_6[15:0];
  wire [15:0]       writeDataVec_data_dataElement_7 = writeDataVec_data_dataIsRead_7 ? waiteReadData_3[15:0] : writeDataVec_data_unreadData_7[15:0];
  wire [31:0]       writeDataVec_data_lo_1 = {writeDataVec_data_dataElement_5, writeDataVec_data_dataElement_4};
  wire [31:0]       writeDataVec_data_hi_1 = {writeDataVec_data_dataElement_7, writeDataVec_data_dataElement_6};
  wire [63:0]       writeDataVec_data_1 = {writeDataVec_data_hi_1, writeDataVec_data_lo_1};
  wire [190:0]      writeDataVec_shifterData_1 = {127'h0, writeDataVec_data_1} << {184'h0, executeIndexVec_1, 5'h0};
  wire [127:0]      writeDataVec_1 = writeDataVec_shifterData_1[127:0];
  wire [31:0]       writeDataVec_data_dataElement_8 = writeDataVec_data_dataIsRead_8 ? waiteReadData_0 : writeDataVec_data_unreadData_8;
  wire [31:0]       writeDataVec_data_dataElement_9 = writeDataVec_data_dataIsRead_9 ? waiteReadData_1 : writeDataVec_data_unreadData_9;
  wire [31:0]       writeDataVec_data_dataElement_10 = writeDataVec_data_dataIsRead_10 ? waiteReadData_2 : writeDataVec_data_unreadData_10;
  wire [31:0]       writeDataVec_data_dataElement_11 = writeDataVec_data_dataIsRead_11 ? waiteReadData_3 : writeDataVec_data_unreadData_11;
  wire [63:0]       writeDataVec_data_lo_2 = {writeDataVec_data_dataElement_9, writeDataVec_data_dataElement_8};
  wire [63:0]       writeDataVec_data_hi_2 = {writeDataVec_data_dataElement_11, writeDataVec_data_dataElement_10};
  wire [127:0]      writeDataVec_data_2 = {writeDataVec_data_hi_2, writeDataVec_data_lo_2};
  wire [190:0]      writeDataVec_shifterData_2 = {63'h0, writeDataVec_data_2};
  wire [127:0]      writeDataVec_2 = writeDataVec_shifterData_2[127:0];
  wire [127:0]      writeData = (sew1H[0] ? writeDataVec_0 : 128'h0) | (sew1H[1] ? writeDataVec_1 : 128'h0) | (sew1H[2] ? writeDataVec_2 : 128'h0);
  wire [1:0]        writeMaskVec_mask_lo = waiteReadDataPipeReg_sourceValid[1:0];
  wire [1:0]        writeMaskVec_mask_hi = waiteReadDataPipeReg_sourceValid[3:2];
  wire [3:0]        writeMaskVec_mask = {writeMaskVec_mask_hi, writeMaskVec_mask_lo};
  wire [18:0]       writeMaskVec_shifterMask = {15'h0, writeMaskVec_mask} << {15'h0, executeIndexVec_0, 2'h0};
  wire [15:0]       writeMaskVec_0 = writeMaskVec_shifterMask[15:0];
  wire [3:0]        writeMaskVec_mask_lo_1 = {{2{waiteReadDataPipeReg_sourceValid[1]}}, {2{waiteReadDataPipeReg_sourceValid[0]}}};
  wire [3:0]        writeMaskVec_mask_hi_1 = {{2{waiteReadDataPipeReg_sourceValid[3]}}, {2{waiteReadDataPipeReg_sourceValid[2]}}};
  wire [7:0]        writeMaskVec_mask_1 = {writeMaskVec_mask_hi_1, writeMaskVec_mask_lo_1};
  wire [22:0]       writeMaskVec_shifterMask_1 = {15'h0, writeMaskVec_mask_1} << {19'h0, executeIndexVec_1, 2'h0};
  wire [15:0]       writeMaskVec_1 = writeMaskVec_shifterMask_1[15:0];
  wire [7:0]        writeMaskVec_mask_lo_2 = {{4{waiteReadDataPipeReg_sourceValid[1]}}, {4{waiteReadDataPipeReg_sourceValid[0]}}};
  wire [7:0]        writeMaskVec_mask_hi_2 = {{4{waiteReadDataPipeReg_sourceValid[3]}}, {4{waiteReadDataPipeReg_sourceValid[2]}}};
  wire [15:0]       writeMaskVec_mask_2 = {writeMaskVec_mask_hi_2, writeMaskVec_mask_lo_2};
  wire [22:0]       writeMaskVec_shifterMask_2 = {7'h0, writeMaskVec_mask_2};
  wire [15:0]       writeMaskVec_2 = writeMaskVec_shifterMask_2[15:0];
  wire [15:0]       writeMask = (sew1H[0] ? writeMaskVec_0 : 16'h0) | (sew1H[1] ? writeMaskVec_1 : 16'h0) | (sew1H[2] ? writeMaskVec_2 : 16'h0);
  wire [9:0]        _writeRequest_res_writeData_groupCounter_T_6 = {3'h0, waiteReadDataPipeReg_executeGroup} << instReg_sew;
  wire [4:0]        writeRequest_0_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_6[6:2];
  wire [4:0]        writeRequest_1_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_6[6:2];
  wire [4:0]        writeRequest_2_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_6[6:2];
  wire [4:0]        writeRequest_3_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_6[6:2];
  wire [31:0]       writeRequest_0_writeData_data = writeData[31:0];
  wire [31:0]       writeRequest_1_writeData_data = writeData[63:32];
  wire [31:0]       writeRequest_2_writeData_data = writeData[95:64];
  wire [31:0]       writeRequest_3_writeData_data = writeData[127:96];
  wire [3:0]        writeRequest_0_writeData_mask = writeMask[3:0];
  wire [3:0]        writeRequest_1_writeData_mask = writeMask[7:4];
  wire [3:0]        writeRequest_2_writeData_mask = writeMask[11:8];
  wire [3:0]        writeRequest_3_writeData_mask = writeMask[15:12];
  wire [1:0]        WillWriteLane_lo = {|writeRequest_1_writeData_mask, |writeRequest_0_writeData_mask};
  wire [1:0]        WillWriteLane_hi = {|writeRequest_3_writeData_mask, |writeRequest_2_writeData_mask};
  wire [3:0]        WillWriteLane = {WillWriteLane_hi, WillWriteLane_lo};
  wire              waiteStageDeqValid = waiteReadStageValid & (waiteReadSate == waiteReadDataPipeReg_needRead | waiteReadDataPipeReg_needRead == 4'h0);
  wire              waiteStageDeqReady;
  wire              waiteStageDeqFire = waiteStageDeqValid & waiteStageDeqReady;
  assign waiteStageEnqReady = ~waiteReadStageValid | waiteStageDeqFire;
  assign readWaitQueue_deq_ready = waiteStageEnqReady;
  wire              waiteStageEnqFire = readWaitQueue_deq_valid & waiteStageEnqReady;
  wire              isWaiteForThisData = waiteReadDataPipeReg_needRead[0] & ~(waiteReadSate[0]) & waiteReadStageValid;
  assign readData_readDataQueue_deq_ready = isWaiteForThisData | unitType[2] | compress | gatherWaiteRead | mvRd;
  assign isWaiteForThisData_1 = waiteReadDataPipeReg_needRead[1] & ~(waiteReadSate[1]) & waiteReadStageValid;
  assign readData_readDataQueue_1_deq_ready = isWaiteForThisData_1;
  assign isWaiteForThisData_2 = waiteReadDataPipeReg_needRead[2] & ~(waiteReadSate[2]) & waiteReadStageValid;
  assign readData_readDataQueue_2_deq_ready = isWaiteForThisData_2;
  assign isWaiteForThisData_3 = waiteReadDataPipeReg_needRead[3] & ~(waiteReadSate[3]) & waiteReadStageValid;
  assign readData_readDataQueue_3_deq_ready = isWaiteForThisData_3;
  wire [1:0]        readResultValid_lo = {readTokenRelease_1, readTokenRelease_0};
  wire [1:0]        readResultValid_hi = {readTokenRelease_3, readTokenRelease_2};
  wire [3:0]        readResultValid = {readResultValid_hi, readResultValid_lo};
  wire              executeEnqValid = otherTypeRequestDeq & ~readType;
  wire [63:0]       source2_lo = {exeReqReg_1_bits_source2, exeReqReg_0_bits_source2};
  wire [63:0]       source2_hi = {exeReqReg_3_bits_source2, exeReqReg_2_bits_source2};
  wire [127:0]      source2 = {source2_hi, source2_lo};
  wire [127:0]      source1 = {source1_hi, source1_lo};
  wire              vs1Split_0_2 = vs1Split_vs1SetIndex;
  wire [1:0]        vs1Split_vs1SetIndex_1 = requestCounter[1:0];
  wire              vs1Split_1_2 = &vs1Split_vs1SetIndex_1;
  wire [2:0]        vs1Split_vs1SetIndex_2 = requestCounter[2:0];
  wire              vs1Split_2_2 = &vs1Split_vs1SetIndex_2;
  wire [15:0]       _compressSource1_T_3 = sew1H[0] ? (vs1Split_vs1SetIndex ? readVS1Reg_data[31:16] : readVS1Reg_data[15:0]) : 16'h0;
  wire [3:0][7:0]   _GEN_47 = {{readVS1Reg_data[31:24]}, {readVS1Reg_data[23:16]}, {readVS1Reg_data[15:8]}, {readVS1Reg_data[7:0]}};
  wire [7:0][3:0]   _GEN_51 = {{readVS1Reg_data[31:28]}, {readVS1Reg_data[27:24]}, {readVS1Reg_data[23:20]}, {readVS1Reg_data[19:16]}, {readVS1Reg_data[15:12]}, {readVS1Reg_data[11:8]}, {readVS1Reg_data[7:4]}, {readVS1Reg_data[3:0]}};
  wire [7:0]        _GEN_52 = _compressSource1_T_3[7:0] | (sew1H[1] ? _GEN_47[vs1Split_vs1SetIndex_1] : 8'h0);
  wire [15:0]       compressSource1 = {_compressSource1_T_3[15:8], _GEN_52[7:4], _GEN_52[3:0] | (sew1H[2] ? _GEN_51[vs1Split_vs1SetIndex_2] : 4'h0)};
  wire [31:0]       source1Select = mv ? readVS1Reg_data : {16'h0, compressSource1};
  wire              source1Change = sew1H[0] & vs1Split_0_2 | sew1H[1] & vs1Split_1_2 | sew1H[2] & vs1Split_2_2;
  assign viotaCounterAdd = executeEnqValid & unitType[1];
  wire [1:0]        view__in_bits_ffoInput_lo = {exeReqReg_1_bits_ffo, exeReqReg_0_bits_ffo};
  wire [1:0]        view__in_bits_ffoInput_hi = {exeReqReg_3_bits_ffo, exeReqReg_2_bits_ffo};
  wire              reduceUnit_in_valid = executeEnqValid & unitType[2];
  wire              _view__firstGroup_T_1 = _reduceUnit_in_ready & reduceUnit_in_valid;
  wire [6:0]        extendGroupCount = extendType ? (subType[2] ? _extendGroupCount_T_1 : {1'h0, requestCounter, executeIndex[1]}) : {2'h0, requestCounter};
  wire [127:0]      _executeResult_T_4 = unitType[1] ? compressUnitResultQueue_deq_bits_data : 128'h0;
  wire [127:0]      executeResult = {_executeResult_T_4[127:32], _executeResult_T_4[31:0] | (unitType[2] ? _reduceUnit_out_bits_data : 32'h0)} | (unitType[3] ? _extendUnit_out : 128'h0);
  assign executeReady = readType | unitType[1] | unitType[2] & _reduceUnit_in_ready & readVS1Reg_dataValid | unitType[3] & executeEnqValid;
  assign compressUnitResultQueue_deq_ready = &{compressUnitResultQueue_deq_ready_hi, compressUnitResultQueue_deq_ready_lo};
  wire              compressDeq = compressUnitResultQueue_deq_ready & compressUnitResultQueue_deq_valid;
  wire              executeValid = unitType[1] & compressDeq | unitType[3] & executeEnqValid;
  assign executeGroupCounter = (unitType[1] | unitType[2] ? requestCounter : 5'h0) | (unitType[3] ? extendGroupCount[4:0] : 5'h0);
  wire [6:0]        executeDeqGroupCounter = {2'h0, (unitType[1] ? compressUnitResultQueue_deq_bits_groupCounter : 5'h0) | (unitType[2] ? requestCounter : 5'h0)} | (unitType[3] ? extendGroupCount : 7'h0);
  wire [15:0]       executeWriteByteMask = compress | ffo | mvVd ? compressUnitResultQueue_deq_bits_mask : executeByteMask;
  wire              maskFilter = |{~maskDestinationType, currentMaskGroupForDestination[31:0]};
  wire              maskFilter_1 = |{~maskDestinationType, currentMaskGroupForDestination[63:32]};
  wire              maskFilter_2 = |{~maskDestinationType, currentMaskGroupForDestination[95:64]};
  wire              maskFilter_3 = |{~maskDestinationType, currentMaskGroupForDestination[127:96]};
  assign writeQueue_0_deq_valid = ~_writeQueue_fifo_empty;
  wire              exeResp_0_valid_0 = writeQueue_0_deq_valid;
  wire              writeQueue_dataOut_ffoByOther;
  wire [31:0]       writeQueue_dataOut_writeData_data;
  wire [31:0]       exeResp_0_bits_data_0 = writeQueue_0_deq_bits_writeData_data;
  wire [3:0]        writeQueue_dataOut_writeData_mask;
  wire [3:0]        exeResp_0_bits_mask_0 = writeQueue_0_deq_bits_writeData_mask;
  wire [4:0]        writeQueue_dataOut_writeData_groupCounter;
  wire [4:0]        writeQueue_dataOut_writeData_vd;
  wire [2:0]        writeQueue_dataOut_index;
  wire [4:0]        writeQueue_0_enq_bits_writeData_groupCounter;
  wire [4:0]        writeQueue_0_enq_bits_writeData_vd;
  wire [9:0]        writeQueue_dataIn_lo = {writeQueue_0_enq_bits_writeData_groupCounter, writeQueue_0_enq_bits_writeData_vd};
  wire [31:0]       writeQueue_0_enq_bits_writeData_data;
  wire [3:0]        writeQueue_0_enq_bits_writeData_mask;
  wire [35:0]       writeQueue_dataIn_hi = {writeQueue_0_enq_bits_writeData_data, writeQueue_0_enq_bits_writeData_mask};
  wire              writeQueue_0_enq_bits_ffoByOther;
  wire [46:0]       writeQueue_dataIn_hi_1 = {writeQueue_0_enq_bits_ffoByOther, writeQueue_dataIn_hi, writeQueue_dataIn_lo};
  wire [49:0]       writeQueue_dataIn = {writeQueue_dataIn_hi_1, writeQueue_0_enq_bits_index};
  assign writeQueue_dataOut_index = _writeQueue_fifo_data_out[2:0];
  assign writeQueue_dataOut_writeData_vd = _writeQueue_fifo_data_out[7:3];
  assign writeQueue_dataOut_writeData_groupCounter = _writeQueue_fifo_data_out[12:8];
  assign writeQueue_dataOut_writeData_mask = _writeQueue_fifo_data_out[16:13];
  assign writeQueue_dataOut_writeData_data = _writeQueue_fifo_data_out[48:17];
  assign writeQueue_dataOut_ffoByOther = _writeQueue_fifo_data_out[49];
  wire              writeQueue_0_deq_bits_ffoByOther = writeQueue_dataOut_ffoByOther;
  assign writeQueue_0_deq_bits_writeData_data = writeQueue_dataOut_writeData_data;
  assign writeQueue_0_deq_bits_writeData_mask = writeQueue_dataOut_writeData_mask;
  wire [4:0]        writeQueue_0_deq_bits_writeData_groupCounter = writeQueue_dataOut_writeData_groupCounter;
  wire [4:0]        writeQueue_0_deq_bits_writeData_vd = writeQueue_dataOut_writeData_vd;
  wire [2:0]        writeQueue_0_deq_bits_index = writeQueue_dataOut_index;
  wire              writeQueue_0_enq_ready = ~_writeQueue_fifo_full;
  wire              writeQueue_0_enq_valid;
  assign writeQueue_1_deq_valid = ~_writeQueue_fifo_1_empty;
  wire              exeResp_1_valid_0 = writeQueue_1_deq_valid;
  wire              writeQueue_dataOut_1_ffoByOther;
  wire [31:0]       writeQueue_dataOut_1_writeData_data;
  wire [31:0]       exeResp_1_bits_data_0 = writeQueue_1_deq_bits_writeData_data;
  wire [3:0]        writeQueue_dataOut_1_writeData_mask;
  wire [3:0]        exeResp_1_bits_mask_0 = writeQueue_1_deq_bits_writeData_mask;
  wire [4:0]        writeQueue_dataOut_1_writeData_groupCounter;
  wire [4:0]        writeQueue_dataOut_1_writeData_vd;
  wire [2:0]        writeQueue_dataOut_1_index;
  wire [4:0]        writeQueue_1_enq_bits_writeData_groupCounter;
  wire [4:0]        writeQueue_1_enq_bits_writeData_vd;
  wire [9:0]        writeQueue_dataIn_lo_1 = {writeQueue_1_enq_bits_writeData_groupCounter, writeQueue_1_enq_bits_writeData_vd};
  wire [31:0]       writeQueue_1_enq_bits_writeData_data;
  wire [3:0]        writeQueue_1_enq_bits_writeData_mask;
  wire [35:0]       writeQueue_dataIn_hi_2 = {writeQueue_1_enq_bits_writeData_data, writeQueue_1_enq_bits_writeData_mask};
  wire              writeQueue_1_enq_bits_ffoByOther;
  wire [46:0]       writeQueue_dataIn_hi_3 = {writeQueue_1_enq_bits_ffoByOther, writeQueue_dataIn_hi_2, writeQueue_dataIn_lo_1};
  wire [49:0]       writeQueue_dataIn_1 = {writeQueue_dataIn_hi_3, writeQueue_1_enq_bits_index};
  assign writeQueue_dataOut_1_index = _writeQueue_fifo_1_data_out[2:0];
  assign writeQueue_dataOut_1_writeData_vd = _writeQueue_fifo_1_data_out[7:3];
  assign writeQueue_dataOut_1_writeData_groupCounter = _writeQueue_fifo_1_data_out[12:8];
  assign writeQueue_dataOut_1_writeData_mask = _writeQueue_fifo_1_data_out[16:13];
  assign writeQueue_dataOut_1_writeData_data = _writeQueue_fifo_1_data_out[48:17];
  assign writeQueue_dataOut_1_ffoByOther = _writeQueue_fifo_1_data_out[49];
  wire              writeQueue_1_deq_bits_ffoByOther = writeQueue_dataOut_1_ffoByOther;
  assign writeQueue_1_deq_bits_writeData_data = writeQueue_dataOut_1_writeData_data;
  assign writeQueue_1_deq_bits_writeData_mask = writeQueue_dataOut_1_writeData_mask;
  wire [4:0]        writeQueue_1_deq_bits_writeData_groupCounter = writeQueue_dataOut_1_writeData_groupCounter;
  wire [4:0]        writeQueue_1_deq_bits_writeData_vd = writeQueue_dataOut_1_writeData_vd;
  wire [2:0]        writeQueue_1_deq_bits_index = writeQueue_dataOut_1_index;
  wire              writeQueue_1_enq_ready = ~_writeQueue_fifo_1_full;
  wire              writeQueue_1_enq_valid;
  assign writeQueue_2_deq_valid = ~_writeQueue_fifo_2_empty;
  wire              exeResp_2_valid_0 = writeQueue_2_deq_valid;
  wire              writeQueue_dataOut_2_ffoByOther;
  wire [31:0]       writeQueue_dataOut_2_writeData_data;
  wire [31:0]       exeResp_2_bits_data_0 = writeQueue_2_deq_bits_writeData_data;
  wire [3:0]        writeQueue_dataOut_2_writeData_mask;
  wire [3:0]        exeResp_2_bits_mask_0 = writeQueue_2_deq_bits_writeData_mask;
  wire [4:0]        writeQueue_dataOut_2_writeData_groupCounter;
  wire [4:0]        writeQueue_dataOut_2_writeData_vd;
  wire [2:0]        writeQueue_dataOut_2_index;
  wire [4:0]        writeQueue_2_enq_bits_writeData_groupCounter;
  wire [4:0]        writeQueue_2_enq_bits_writeData_vd;
  wire [9:0]        writeQueue_dataIn_lo_2 = {writeQueue_2_enq_bits_writeData_groupCounter, writeQueue_2_enq_bits_writeData_vd};
  wire [31:0]       writeQueue_2_enq_bits_writeData_data;
  wire [3:0]        writeQueue_2_enq_bits_writeData_mask;
  wire [35:0]       writeQueue_dataIn_hi_4 = {writeQueue_2_enq_bits_writeData_data, writeQueue_2_enq_bits_writeData_mask};
  wire              writeQueue_2_enq_bits_ffoByOther;
  wire [46:0]       writeQueue_dataIn_hi_5 = {writeQueue_2_enq_bits_ffoByOther, writeQueue_dataIn_hi_4, writeQueue_dataIn_lo_2};
  wire [49:0]       writeQueue_dataIn_2 = {writeQueue_dataIn_hi_5, writeQueue_2_enq_bits_index};
  assign writeQueue_dataOut_2_index = _writeQueue_fifo_2_data_out[2:0];
  assign writeQueue_dataOut_2_writeData_vd = _writeQueue_fifo_2_data_out[7:3];
  assign writeQueue_dataOut_2_writeData_groupCounter = _writeQueue_fifo_2_data_out[12:8];
  assign writeQueue_dataOut_2_writeData_mask = _writeQueue_fifo_2_data_out[16:13];
  assign writeQueue_dataOut_2_writeData_data = _writeQueue_fifo_2_data_out[48:17];
  assign writeQueue_dataOut_2_ffoByOther = _writeQueue_fifo_2_data_out[49];
  wire              writeQueue_2_deq_bits_ffoByOther = writeQueue_dataOut_2_ffoByOther;
  assign writeQueue_2_deq_bits_writeData_data = writeQueue_dataOut_2_writeData_data;
  assign writeQueue_2_deq_bits_writeData_mask = writeQueue_dataOut_2_writeData_mask;
  wire [4:0]        writeQueue_2_deq_bits_writeData_groupCounter = writeQueue_dataOut_2_writeData_groupCounter;
  wire [4:0]        writeQueue_2_deq_bits_writeData_vd = writeQueue_dataOut_2_writeData_vd;
  wire [2:0]        writeQueue_2_deq_bits_index = writeQueue_dataOut_2_index;
  wire              writeQueue_2_enq_ready = ~_writeQueue_fifo_2_full;
  wire              writeQueue_2_enq_valid;
  assign writeQueue_3_deq_valid = ~_writeQueue_fifo_3_empty;
  wire              exeResp_3_valid_0 = writeQueue_3_deq_valid;
  wire              writeQueue_dataOut_3_ffoByOther;
  wire [31:0]       writeQueue_dataOut_3_writeData_data;
  wire [31:0]       exeResp_3_bits_data_0 = writeQueue_3_deq_bits_writeData_data;
  wire [3:0]        writeQueue_dataOut_3_writeData_mask;
  wire [3:0]        exeResp_3_bits_mask_0 = writeQueue_3_deq_bits_writeData_mask;
  wire [4:0]        writeQueue_dataOut_3_writeData_groupCounter;
  wire [4:0]        writeQueue_dataOut_3_writeData_vd;
  wire [2:0]        writeQueue_dataOut_3_index;
  wire [4:0]        writeQueue_3_enq_bits_writeData_groupCounter;
  wire [4:0]        writeQueue_3_enq_bits_writeData_vd;
  wire [9:0]        writeQueue_dataIn_lo_3 = {writeQueue_3_enq_bits_writeData_groupCounter, writeQueue_3_enq_bits_writeData_vd};
  wire [31:0]       writeQueue_3_enq_bits_writeData_data;
  wire [3:0]        writeQueue_3_enq_bits_writeData_mask;
  wire [35:0]       writeQueue_dataIn_hi_6 = {writeQueue_3_enq_bits_writeData_data, writeQueue_3_enq_bits_writeData_mask};
  wire              writeQueue_3_enq_bits_ffoByOther;
  wire [46:0]       writeQueue_dataIn_hi_7 = {writeQueue_3_enq_bits_ffoByOther, writeQueue_dataIn_hi_6, writeQueue_dataIn_lo_3};
  wire [49:0]       writeQueue_dataIn_3 = {writeQueue_dataIn_hi_7, writeQueue_3_enq_bits_index};
  assign writeQueue_dataOut_3_index = _writeQueue_fifo_3_data_out[2:0];
  assign writeQueue_dataOut_3_writeData_vd = _writeQueue_fifo_3_data_out[7:3];
  assign writeQueue_dataOut_3_writeData_groupCounter = _writeQueue_fifo_3_data_out[12:8];
  assign writeQueue_dataOut_3_writeData_mask = _writeQueue_fifo_3_data_out[16:13];
  assign writeQueue_dataOut_3_writeData_data = _writeQueue_fifo_3_data_out[48:17];
  assign writeQueue_dataOut_3_ffoByOther = _writeQueue_fifo_3_data_out[49];
  wire              writeQueue_3_deq_bits_ffoByOther = writeQueue_dataOut_3_ffoByOther;
  assign writeQueue_3_deq_bits_writeData_data = writeQueue_dataOut_3_writeData_data;
  assign writeQueue_3_deq_bits_writeData_mask = writeQueue_dataOut_3_writeData_mask;
  wire [4:0]        writeQueue_3_deq_bits_writeData_groupCounter = writeQueue_dataOut_3_writeData_groupCounter;
  wire [4:0]        writeQueue_3_deq_bits_writeData_vd = writeQueue_dataOut_3_writeData_vd;
  wire [2:0]        writeQueue_3_deq_bits_index = writeQueue_dataOut_3_index;
  wire              writeQueue_3_enq_ready = ~_writeQueue_fifo_3_full;
  wire              writeQueue_3_enq_valid;
  wire              dataNotInShifter_readTypeWriteVrf = waiteStageDeqFire & WillWriteLane[0];
  assign writeQueue_0_enq_valid = _maskedWrite_out_0_valid | dataNotInShifter_readTypeWriteVrf;
  assign writeQueue_0_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf ? writeRequest_0_writeData_vd : 5'h0;
  assign writeQueue_0_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf ? writeRequest_0_writeData_groupCounter : _maskedWrite_out_0_bits_writeData_groupCounter;
  assign writeQueue_0_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf ? writeRequest_0_writeData_mask : _maskedWrite_out_0_bits_writeData_mask;
  assign writeQueue_0_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf ? writeRequest_0_writeData_data : _maskedWrite_out_0_bits_writeData_data;
  assign writeQueue_0_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf & _maskedWrite_out_0_bits_ffoByOther;
  wire [4:0]        exeResp_0_bits_vd_0 = instReg_vd + {1'h0, writeQueue_0_deq_bits_writeData_groupCounter[4:1]};
  wire              exeResp_0_bits_offset_0 = writeQueue_0_deq_bits_writeData_groupCounter[0];
  reg  [2:0]        dataNotInShifter_writeTokenCounter;
  wire              _dataNotInShifter_T = exeResp_0_ready_0 & exeResp_0_valid_0;
  wire [2:0]        dataNotInShifter_writeTokenChange = _dataNotInShifter_T ? 3'h1 : 3'h7;
  wire              dataNotInShifter_readTypeWriteVrf_1 = waiteStageDeqFire & WillWriteLane[1];
  assign writeQueue_1_enq_valid = _maskedWrite_out_1_valid | dataNotInShifter_readTypeWriteVrf_1;
  assign writeQueue_1_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_1 ? writeRequest_1_writeData_vd : 5'h0;
  assign writeQueue_1_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_1 ? writeRequest_1_writeData_groupCounter : _maskedWrite_out_1_bits_writeData_groupCounter;
  assign writeQueue_1_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_1 ? writeRequest_1_writeData_mask : _maskedWrite_out_1_bits_writeData_mask;
  assign writeQueue_1_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_1 ? writeRequest_1_writeData_data : _maskedWrite_out_1_bits_writeData_data;
  assign writeQueue_1_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_1 & _maskedWrite_out_1_bits_ffoByOther;
  wire [4:0]        exeResp_1_bits_vd_0 = instReg_vd + {1'h0, writeQueue_1_deq_bits_writeData_groupCounter[4:1]};
  wire              exeResp_1_bits_offset_0 = writeQueue_1_deq_bits_writeData_groupCounter[0];
  reg  [2:0]        dataNotInShifter_writeTokenCounter_1;
  wire              _dataNotInShifter_T_3 = exeResp_1_ready_0 & exeResp_1_valid_0;
  wire [2:0]        dataNotInShifter_writeTokenChange_1 = _dataNotInShifter_T_3 ? 3'h1 : 3'h7;
  wire              dataNotInShifter_readTypeWriteVrf_2 = waiteStageDeqFire & WillWriteLane[2];
  assign writeQueue_2_enq_valid = _maskedWrite_out_2_valid | dataNotInShifter_readTypeWriteVrf_2;
  assign writeQueue_2_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_2 ? writeRequest_2_writeData_vd : 5'h0;
  assign writeQueue_2_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_2 ? writeRequest_2_writeData_groupCounter : _maskedWrite_out_2_bits_writeData_groupCounter;
  assign writeQueue_2_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_2 ? writeRequest_2_writeData_mask : _maskedWrite_out_2_bits_writeData_mask;
  assign writeQueue_2_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_2 ? writeRequest_2_writeData_data : _maskedWrite_out_2_bits_writeData_data;
  assign writeQueue_2_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_2 & _maskedWrite_out_2_bits_ffoByOther;
  wire [4:0]        exeResp_2_bits_vd_0 = instReg_vd + {1'h0, writeQueue_2_deq_bits_writeData_groupCounter[4:1]};
  wire              exeResp_2_bits_offset_0 = writeQueue_2_deq_bits_writeData_groupCounter[0];
  reg  [2:0]        dataNotInShifter_writeTokenCounter_2;
  wire              _dataNotInShifter_T_6 = exeResp_2_ready_0 & exeResp_2_valid_0;
  wire [2:0]        dataNotInShifter_writeTokenChange_2 = _dataNotInShifter_T_6 ? 3'h1 : 3'h7;
  wire              dataNotInShifter_readTypeWriteVrf_3 = waiteStageDeqFire & WillWriteLane[3];
  assign writeQueue_3_enq_valid = _maskedWrite_out_3_valid | dataNotInShifter_readTypeWriteVrf_3;
  assign writeQueue_3_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_3 ? writeRequest_3_writeData_vd : 5'h0;
  assign writeQueue_3_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_3 ? writeRequest_3_writeData_groupCounter : _maskedWrite_out_3_bits_writeData_groupCounter;
  assign writeQueue_3_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_3 ? writeRequest_3_writeData_mask : _maskedWrite_out_3_bits_writeData_mask;
  assign writeQueue_3_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_3 ? writeRequest_3_writeData_data : _maskedWrite_out_3_bits_writeData_data;
  assign writeQueue_3_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_3 & _maskedWrite_out_3_bits_ffoByOther;
  wire [4:0]        exeResp_3_bits_vd_0 = instReg_vd + {1'h0, writeQueue_3_deq_bits_writeData_groupCounter[4:1]};
  wire              exeResp_3_bits_offset_0 = writeQueue_3_deq_bits_writeData_groupCounter[0];
  reg  [2:0]        dataNotInShifter_writeTokenCounter_3;
  wire              _dataNotInShifter_T_9 = exeResp_3_ready_0 & exeResp_3_valid_0;
  wire [2:0]        dataNotInShifter_writeTokenChange_3 = _dataNotInShifter_T_9 ? 3'h1 : 3'h7;
  wire              dataNotInShifter = dataNotInShifter_writeTokenCounter == 3'h0 & dataNotInShifter_writeTokenCounter_1 == 3'h0 & dataNotInShifter_writeTokenCounter_2 == 3'h0 & dataNotInShifter_writeTokenCounter_3 == 3'h0;
  assign waiteStageDeqReady = (~(WillWriteLane[0]) | writeQueue_0_enq_ready) & (~(WillWriteLane[1]) | writeQueue_1_enq_ready) & (~(WillWriteLane[2]) | writeQueue_2_enq_ready) & (~(WillWriteLane[3]) | writeQueue_3_enq_ready);
  reg               waiteLastRequest;
  reg               waitQueueClear;
  wire              lastReportValid = waitQueueClear & ~(writeQueue_0_deq_valid | writeQueue_1_deq_valid | writeQueue_2_deq_valid | writeQueue_3_deq_valid) & dataNotInShifter;
  wire              executeStageInvalid = unitType[1] & ~compressUnitResultQueue_deq_valid & ~_compressUnit_stageValid | unitType[2] & _reduceUnit_in_ready | unitType[3];
  wire              executeStageClean = readType ? waiteStageDeqFire & waiteReadDataPipeReg_last : waiteLastRequest & _maskedWrite_stageClear & executeStageInvalid;
  wire              invalidEnq = instReq_valid & instReq_bits_vl == 9'h0 & ~enqMvRD;
  wire [7:0]        _lastReport_output = lastReportValid ? 8'h1 << instReg_instructionIndex : 8'h0;
  wire [31:0]       gatherData_bits_0 = readVS1Reg_dataValid ? readVS1Reg_data : 32'h0;
  always @(posedge clock) begin
    if (reset) begin
      v0_0 <= 32'h0;
      v0_1 <= 32'h0;
      v0_2 <= 32'h0;
      v0_3 <= 32'h0;
      v0_4 <= 32'h0;
      v0_5 <= 32'h0;
      v0_6 <= 32'h0;
      v0_7 <= 32'h0;
      gatherReadState <= 2'h0;
      gatherDatOffset <= 2'h0;
      gatherLane <= 2'h0;
      gatherOffset <= 1'h0;
      gatherGrowth <= 3'h0;
      instReg_instructionIndex <= 3'h0;
      instReg_decodeResult_specialSlot <= 1'h0;
      instReg_decodeResult_topUop <= 5'h0;
      instReg_decodeResult_popCount <= 1'h0;
      instReg_decodeResult_ffo <= 1'h0;
      instReg_decodeResult_average <= 1'h0;
      instReg_decodeResult_reverse <= 1'h0;
      instReg_decodeResult_dontNeedExecuteInLane <= 1'h0;
      instReg_decodeResult_scheduler <= 1'h0;
      instReg_decodeResult_sReadVD <= 1'h0;
      instReg_decodeResult_vtype <= 1'h0;
      instReg_decodeResult_sWrite <= 1'h0;
      instReg_decodeResult_crossRead <= 1'h0;
      instReg_decodeResult_crossWrite <= 1'h0;
      instReg_decodeResult_maskUnit <= 1'h0;
      instReg_decodeResult_special <= 1'h0;
      instReg_decodeResult_saturate <= 1'h0;
      instReg_decodeResult_vwmacc <= 1'h0;
      instReg_decodeResult_readOnly <= 1'h0;
      instReg_decodeResult_maskSource <= 1'h0;
      instReg_decodeResult_maskDestination <= 1'h0;
      instReg_decodeResult_maskLogic <= 1'h0;
      instReg_decodeResult_uop <= 4'h0;
      instReg_decodeResult_iota <= 1'h0;
      instReg_decodeResult_mv <= 1'h0;
      instReg_decodeResult_extend <= 1'h0;
      instReg_decodeResult_unOrderWrite <= 1'h0;
      instReg_decodeResult_compress <= 1'h0;
      instReg_decodeResult_gather16 <= 1'h0;
      instReg_decodeResult_gather <= 1'h0;
      instReg_decodeResult_slid <= 1'h0;
      instReg_decodeResult_targetRd <= 1'h0;
      instReg_decodeResult_widenReduce <= 1'h0;
      instReg_decodeResult_red <= 1'h0;
      instReg_decodeResult_nr <= 1'h0;
      instReg_decodeResult_itype <= 1'h0;
      instReg_decodeResult_unsigned1 <= 1'h0;
      instReg_decodeResult_unsigned0 <= 1'h0;
      instReg_decodeResult_other <= 1'h0;
      instReg_decodeResult_multiCycle <= 1'h0;
      instReg_decodeResult_divider <= 1'h0;
      instReg_decodeResult_multiplier <= 1'h0;
      instReg_decodeResult_shift <= 1'h0;
      instReg_decodeResult_adder <= 1'h0;
      instReg_decodeResult_logic <= 1'h0;
      instReg_readFromScala <= 32'h0;
      instReg_sew <= 2'h0;
      instReg_vlmul <= 3'h0;
      instReg_maskType <= 1'h0;
      instReg_vxrm <= 3'h0;
      instReg_vs2 <= 5'h0;
      instReg_vs1 <= 5'h0;
      instReg_vd <= 5'h0;
      instReg_vl <= 9'h0;
      instVlValid <= 1'h0;
      readVS1Reg_dataValid <= 1'h0;
      readVS1Reg_requestSend <= 1'h0;
      readVS1Reg_sendToExecution <= 1'h0;
      readVS1Reg_data <= 32'h0;
      readVS1Reg_readIndex <= 4'h0;
      exeReqReg_0_valid <= 1'h0;
      exeReqReg_0_bits_source1 <= 32'h0;
      exeReqReg_0_bits_source2 <= 32'h0;
      exeReqReg_0_bits_index <= 3'h0;
      exeReqReg_0_bits_ffo <= 1'h0;
      exeReqReg_1_valid <= 1'h0;
      exeReqReg_1_bits_source1 <= 32'h0;
      exeReqReg_1_bits_source2 <= 32'h0;
      exeReqReg_1_bits_index <= 3'h0;
      exeReqReg_1_bits_ffo <= 1'h0;
      exeReqReg_2_valid <= 1'h0;
      exeReqReg_2_bits_source1 <= 32'h0;
      exeReqReg_2_bits_source2 <= 32'h0;
      exeReqReg_2_bits_index <= 3'h0;
      exeReqReg_2_bits_ffo <= 1'h0;
      exeReqReg_3_valid <= 1'h0;
      exeReqReg_3_bits_source1 <= 32'h0;
      exeReqReg_3_bits_source2 <= 32'h0;
      exeReqReg_3_bits_index <= 3'h0;
      exeReqReg_3_bits_ffo <= 1'h0;
      requestCounter <= 5'h0;
      executeIndex <= 2'h0;
      readIssueStageState_groupReadState <= 4'h0;
      readIssueStageState_needRead <= 4'h0;
      readIssueStageState_elementValid <= 4'h0;
      readIssueStageState_replaceVs1 <= 4'h0;
      readIssueStageState_readOffset <= 4'h0;
      readIssueStageState_accessLane_0 <= 2'h0;
      readIssueStageState_accessLane_1 <= 2'h0;
      readIssueStageState_accessLane_2 <= 2'h0;
      readIssueStageState_accessLane_3 <= 2'h0;
      readIssueStageState_vsGrowth_0 <= 3'h0;
      readIssueStageState_vsGrowth_1 <= 3'h0;
      readIssueStageState_vsGrowth_2 <= 3'h0;
      readIssueStageState_vsGrowth_3 <= 3'h0;
      readIssueStageState_executeGroup <= 7'h0;
      readIssueStageState_readDataOffset <= 8'h0;
      readIssueStageState_last <= 1'h0;
      readIssueStageValid <= 1'h0;
      tokenCheck_counter <= 4'h0;
      tokenCheck_counter_1 <= 4'h0;
      tokenCheck_counter_2 <= 4'h0;
      tokenCheck_counter_3 <= 4'h0;
      reorderQueueAllocate_counter <= 4'h0;
      reorderQueueAllocate_counterWillUpdate <= 4'h0;
      reorderQueueAllocate_counter_1 <= 4'h0;
      reorderQueueAllocate_counterWillUpdate_1 <= 4'h0;
      reorderQueueAllocate_counter_2 <= 4'h0;
      reorderQueueAllocate_counterWillUpdate_2 <= 4'h0;
      reorderQueueAllocate_counter_3 <= 4'h0;
      reorderQueueAllocate_counterWillUpdate_3 <= 4'h0;
      reorderStageValid <= 1'h0;
      reorderStageState_0 <= 3'h0;
      reorderStageState_1 <= 3'h0;
      reorderStageState_2 <= 3'h0;
      reorderStageState_3 <= 3'h0;
      reorderStageNeed_0 <= 3'h0;
      reorderStageNeed_1 <= 3'h0;
      reorderStageNeed_2 <= 3'h0;
      reorderStageNeed_3 <= 3'h0;
      waiteReadDataPipeReg_executeGroup <= 7'h0;
      waiteReadDataPipeReg_sourceValid <= 4'h0;
      waiteReadDataPipeReg_replaceVs1 <= 4'h0;
      waiteReadDataPipeReg_needRead <= 4'h0;
      waiteReadDataPipeReg_last <= 1'h0;
      waiteReadData_0 <= 32'h0;
      waiteReadData_1 <= 32'h0;
      waiteReadData_2 <= 32'h0;
      waiteReadData_3 <= 32'h0;
      waiteReadSate <= 4'h0;
      waiteReadStageValid <= 1'h0;
      dataNotInShifter_writeTokenCounter <= 3'h0;
      dataNotInShifter_writeTokenCounter_1 <= 3'h0;
      dataNotInShifter_writeTokenCounter_2 <= 3'h0;
      dataNotInShifter_writeTokenCounter_3 <= 3'h0;
      waiteLastRequest <= 1'h0;
      waitQueueClear <= 1'h0;
    end
    else begin
      automatic logic _GEN_48 = instReq_valid & (viotaReq | enqMvRD) | gatherRequestFire;
      automatic logic _GEN_49;
      automatic logic _GEN_50 = source1Change & viotaCounterAdd;
      _GEN_49 = instReq_valid | gatherRequestFire;
      if (v0UpdateVec_0_valid & ~v0UpdateVec_0_bits_offset)
        v0_0 <= v0_0 & ~maskExt | maskExt & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & ~v0UpdateVec_1_bits_offset)
        v0_1 <= v0_1 & ~maskExt_1 | maskExt_1 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & ~v0UpdateVec_2_bits_offset)
        v0_2 <= v0_2 & ~maskExt_2 | maskExt_2 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & ~v0UpdateVec_3_bits_offset)
        v0_3 <= v0_3 & ~maskExt_3 | maskExt_3 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset)
        v0_4 <= v0_4 & ~maskExt_4 | maskExt_4 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset)
        v0_5 <= v0_5 & ~maskExt_5 | maskExt_5 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset)
        v0_6 <= v0_6 & ~maskExt_6 | maskExt_6 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset)
        v0_7 <= v0_7 & ~maskExt_7 | maskExt_7 & v0UpdateVec_3_bits_data;
      if (gatherData_ready_0 & gatherData_valid_0)
        gatherReadState <= 2'h0;
      else if (_tokenCheck_T & gatherSRead)
        gatherReadState <= 2'h2;
      else if (gatherRequestFire)
        gatherReadState <= {notNeedRead, 1'h1};
      else if (readTokenRelease_0 & gatherWaiteRead)
        gatherReadState <= 2'h3;
      if (gatherRequestFire) begin
        gatherDatOffset <= dataOffset;
        gatherLane <= accessLane;
        gatherOffset <= offset;
        gatherGrowth <= reallyGrowth;
      end
      if (_GEN_48 | instReq_valid)
        instReg_instructionIndex <= instReq_bits_instructionIndex;
      if (instReq_valid) begin
        instReg_decodeResult_specialSlot <= instReq_bits_decodeResult_specialSlot;
        instReg_decodeResult_topUop <= instReq_bits_decodeResult_topUop;
        instReg_decodeResult_popCount <= instReq_bits_decodeResult_popCount;
        instReg_decodeResult_ffo <= instReq_bits_decodeResult_ffo;
        instReg_decodeResult_average <= instReq_bits_decodeResult_average;
        instReg_decodeResult_reverse <= instReq_bits_decodeResult_reverse;
        instReg_decodeResult_dontNeedExecuteInLane <= instReq_bits_decodeResult_dontNeedExecuteInLane;
        instReg_decodeResult_scheduler <= instReq_bits_decodeResult_scheduler;
        instReg_decodeResult_sReadVD <= instReq_bits_decodeResult_sReadVD;
        instReg_decodeResult_vtype <= instReq_bits_decodeResult_vtype;
        instReg_decodeResult_sWrite <= instReq_bits_decodeResult_sWrite;
        instReg_decodeResult_crossRead <= instReq_bits_decodeResult_crossRead;
        instReg_decodeResult_crossWrite <= instReq_bits_decodeResult_crossWrite;
        instReg_decodeResult_maskUnit <= instReq_bits_decodeResult_maskUnit;
        instReg_decodeResult_special <= instReq_bits_decodeResult_special;
        instReg_decodeResult_saturate <= instReq_bits_decodeResult_saturate;
        instReg_decodeResult_vwmacc <= instReq_bits_decodeResult_vwmacc;
        instReg_decodeResult_readOnly <= instReq_bits_decodeResult_readOnly;
        instReg_decodeResult_maskSource <= instReq_bits_decodeResult_maskSource;
        instReg_decodeResult_maskDestination <= instReq_bits_decodeResult_maskDestination;
        instReg_decodeResult_maskLogic <= instReq_bits_decodeResult_maskLogic;
        instReg_decodeResult_uop <= instReq_bits_decodeResult_uop;
        instReg_decodeResult_iota <= instReq_bits_decodeResult_iota;
        instReg_decodeResult_mv <= instReq_bits_decodeResult_mv;
        instReg_decodeResult_extend <= instReq_bits_decodeResult_extend;
        instReg_decodeResult_unOrderWrite <= instReq_bits_decodeResult_unOrderWrite;
        instReg_decodeResult_compress <= instReq_bits_decodeResult_compress;
        instReg_decodeResult_gather16 <= instReq_bits_decodeResult_gather16;
        instReg_decodeResult_gather <= instReq_bits_decodeResult_gather;
        instReg_decodeResult_slid <= instReq_bits_decodeResult_slid;
        instReg_decodeResult_targetRd <= instReq_bits_decodeResult_targetRd;
        instReg_decodeResult_widenReduce <= instReq_bits_decodeResult_widenReduce;
        instReg_decodeResult_red <= instReq_bits_decodeResult_red;
        instReg_decodeResult_nr <= instReq_bits_decodeResult_nr;
        instReg_decodeResult_itype <= instReq_bits_decodeResult_itype;
        instReg_decodeResult_unsigned1 <= instReq_bits_decodeResult_unsigned1;
        instReg_decodeResult_unsigned0 <= instReq_bits_decodeResult_unsigned0;
        instReg_decodeResult_other <= instReq_bits_decodeResult_other;
        instReg_decodeResult_multiCycle <= instReq_bits_decodeResult_multiCycle;
        instReg_decodeResult_divider <= instReq_bits_decodeResult_divider;
        instReg_decodeResult_multiplier <= instReq_bits_decodeResult_multiplier;
        instReg_decodeResult_shift <= instReq_bits_decodeResult_shift;
        instReg_decodeResult_adder <= instReq_bits_decodeResult_adder;
        instReg_decodeResult_logic <= instReq_bits_decodeResult_logic;
        instReg_readFromScala <= instReq_bits_readFromScala;
        instReg_sew <= instReq_bits_sew;
        instReg_vlmul <= instReq_bits_vlmul;
        instReg_maskType <= instReq_bits_maskType;
        instReg_vxrm <= instReq_bits_vxrm;
        instReg_vs2 <= instReq_bits_vs2;
        instReg_vd <= instReq_bits_vd;
        instReg_vl <= instReq_bits_vl;
      end
      if (_GEN_48)
        instReg_vs1 <= instReq_bits_vs2;
      else if (instReq_valid)
        instReg_vs1 <= instReq_bits_vs1;
      if (|{instReq_valid, _lastReport_output})
        instVlValid <= ((|instReq_bits_vl) | enqMvRD) & instReq_valid;
      readVS1Reg_dataValid <= ~_GEN_50 & (readTokenRelease_0 | ~_GEN_49 & readVS1Reg_dataValid);
      readVS1Reg_requestSend <= ~_GEN_50 & (_tokenCheck_T | ~_GEN_49 & readVS1Reg_requestSend);
      readVS1Reg_sendToExecution <= _view__firstGroup_T_1 | viotaCounterAdd | ~_GEN_49 & readVS1Reg_sendToExecution;
      if (readTokenRelease_0) begin
        readVS1Reg_data <= readData_readDataQueue_deq_bits;
        waiteReadData_0 <= readData_readDataQueue_deq_bits;
      end
      if (_GEN_50)
        readVS1Reg_readIndex <= readVS1Reg_readIndex + 4'h1;
      else if (_GEN_49)
        readVS1Reg_readIndex <= 4'h0;
      if (tokenIO_0_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_0_valid <= tokenIO_0_maskRequestRelease_0 & ~viota;
      if (tokenIO_0_maskRequestRelease_0) begin
        exeReqReg_0_bits_source1 <= exeRequestQueue_0_deq_bits_source1;
        exeReqReg_0_bits_source2 <= exeRequestQueue_0_deq_bits_source2;
        exeReqReg_0_bits_index <= exeRequestQueue_0_deq_bits_index;
        exeReqReg_0_bits_ffo <= exeRequestQueue_0_deq_bits_ffo;
      end
      if (tokenIO_1_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_1_valid <= tokenIO_1_maskRequestRelease_0 & ~viota;
      if (tokenIO_1_maskRequestRelease_0) begin
        exeReqReg_1_bits_source1 <= exeRequestQueue_1_deq_bits_source1;
        exeReqReg_1_bits_source2 <= exeRequestQueue_1_deq_bits_source2;
        exeReqReg_1_bits_index <= exeRequestQueue_1_deq_bits_index;
        exeReqReg_1_bits_ffo <= exeRequestQueue_1_deq_bits_ffo;
      end
      if (tokenIO_2_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_2_valid <= tokenIO_2_maskRequestRelease_0 & ~viota;
      if (tokenIO_2_maskRequestRelease_0) begin
        exeReqReg_2_bits_source1 <= exeRequestQueue_2_deq_bits_source1;
        exeReqReg_2_bits_source2 <= exeRequestQueue_2_deq_bits_source2;
        exeReqReg_2_bits_index <= exeRequestQueue_2_deq_bits_index;
        exeReqReg_2_bits_ffo <= exeRequestQueue_2_deq_bits_ffo;
      end
      if (tokenIO_3_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_3_valid <= tokenIO_3_maskRequestRelease_0 & ~viota;
      if (tokenIO_3_maskRequestRelease_0) begin
        exeReqReg_3_bits_source1 <= exeRequestQueue_3_deq_bits_source1;
        exeReqReg_3_bits_source2 <= exeRequestQueue_3_deq_bits_source2;
        exeReqReg_3_bits_index <= exeRequestQueue_3_deq_bits_index;
        exeReqReg_3_bits_ffo <= exeRequestQueue_3_deq_bits_ffo;
      end
      if (instReq_valid | groupCounterAdd)
        requestCounter <= instReq_valid ? 5'h0 : requestCounter + 5'h1;
      if (requestStageDeq & anyDataValid)
        executeIndex <= executeIndex + executeIndexGrowth[1:0];
      if (readIssueStageEnq) begin
        readIssueStageState_groupReadState <= 4'h0;
        readIssueStageState_needRead <= _GEN_41 ? _slideAddressGen_indexDeq_bits_needRead : ~notReadSelect;
        readIssueStageState_elementValid <= _GEN_41 ? _slideAddressGen_indexDeq_bits_elementValid : elementValidSelect;
        readIssueStageState_replaceVs1 <= _GEN_41 ? _slideAddressGen_indexDeq_bits_replaceVs1 : 4'h0;
        readIssueStageState_readOffset <= _GEN_41 ? _slideAddressGen_indexDeq_bits_readOffset : offsetSelect;
        readIssueStageState_accessLane_0 <= _GEN_41 ? _slideAddressGen_indexDeq_bits_accessLane_0 : accessLaneSelect[1:0];
        readIssueStageState_accessLane_1 <= _GEN_41 ? _slideAddressGen_indexDeq_bits_accessLane_1 : accessLaneSelect[3:2];
        readIssueStageState_accessLane_2 <= _GEN_41 ? _slideAddressGen_indexDeq_bits_accessLane_2 : accessLaneSelect[5:4];
        readIssueStageState_accessLane_3 <= _GEN_41 ? _slideAddressGen_indexDeq_bits_accessLane_3 : accessLaneSelect[7:6];
        readIssueStageState_vsGrowth_0 <= _GEN_41 ? _slideAddressGen_indexDeq_bits_vsGrowth_0 : growthSelect[2:0];
        readIssueStageState_vsGrowth_1 <= _GEN_41 ? _slideAddressGen_indexDeq_bits_vsGrowth_1 : growthSelect[5:3];
        readIssueStageState_vsGrowth_2 <= _GEN_41 ? _slideAddressGen_indexDeq_bits_vsGrowth_2 : growthSelect[8:6];
        readIssueStageState_vsGrowth_3 <= _GEN_41 ? _slideAddressGen_indexDeq_bits_vsGrowth_3 : growthSelect[11:9];
        readIssueStageState_executeGroup <= _GEN_41 ? _slideAddressGen_indexDeq_bits_executeGroup : executeGroup;
        readIssueStageState_readDataOffset <= _GEN_41 ? _slideAddressGen_indexDeq_bits_readDataOffset : dataOffsetSelect;
        readIssueStageState_last <= _GEN_41 ? _slideAddressGen_indexDeq_bits_last : isVlBoundary;
      end
      else if (anyReadFire)
        readIssueStageState_groupReadState <= readStateUpdate;
      if (readTypeRequestDeq ^ readIssueStageEnq)
        readIssueStageValid <= readIssueStageEnq;
      if (_tokenCheck_T ^ readTokenRelease_0)
        tokenCheck_counter <= tokenCheck_counter + tokenCheck_counterChange;
      if (pipeReadFire_1 ^ readTokenRelease_1)
        tokenCheck_counter_1 <= tokenCheck_counter_1 + tokenCheck_counterChange_1;
      if (pipeReadFire_2 ^ readTokenRelease_2)
        tokenCheck_counter_2 <= tokenCheck_counter_2 + tokenCheck_counterChange_2;
      if (pipeReadFire_3 ^ readTokenRelease_3)
        tokenCheck_counter_3 <= tokenCheck_counter_3 + tokenCheck_counterChange_3;
      if (reorderQueueAllocate_release | readIssueStageEnq) begin
        reorderQueueAllocate_counter <= reorderQueueAllocate_counterUpdate;
        reorderQueueAllocate_counterWillUpdate <= reorderQueueAllocate_counterUpdate + 4'h4;
      end
      if (reorderQueueAllocate_release_1 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_1 <= reorderQueueAllocate_counterUpdate_1;
        reorderQueueAllocate_counterWillUpdate_1 <= reorderQueueAllocate_counterUpdate_1 + 4'h4;
      end
      if (reorderQueueAllocate_release_2 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_2 <= reorderQueueAllocate_counterUpdate_2;
        reorderQueueAllocate_counterWillUpdate_2 <= reorderQueueAllocate_counterUpdate_2 + 4'h4;
      end
      if (reorderQueueAllocate_release_3 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_3 <= reorderQueueAllocate_counterUpdate_3;
        reorderQueueAllocate_counterWillUpdate_3 <= reorderQueueAllocate_counterUpdate_3 + 4'h4;
      end
      if (reorderStageEnqFire ^ reorderStageDeqFire)
        reorderStageValid <= reorderStageEnqFire;
      if (_write1HPipe_0_T & readType)
        reorderStageState_0 <= reorderStageState_0 + 3'h1;
      else if (reorderStageEnqFire)
        reorderStageState_0 <= 3'h0;
      if (_write1HPipe_1_T & readType)
        reorderStageState_1 <= reorderStageState_1 + 3'h1;
      else if (reorderStageEnqFire)
        reorderStageState_1 <= 3'h0;
      if (_write1HPipe_2_T & readType)
        reorderStageState_2 <= reorderStageState_2 + 3'h1;
      else if (reorderStageEnqFire)
        reorderStageState_2 <= 3'h0;
      if (_write1HPipe_3_T & readType)
        reorderStageState_3 <= reorderStageState_3 + 3'h1;
      else if (reorderStageEnqFire)
        reorderStageState_3 <= 3'h0;
      if (reorderStageEnqFire) begin
        reorderStageNeed_0 <= accessCountQueue_deq_bits_0;
        reorderStageNeed_1 <= accessCountQueue_deq_bits_1;
        reorderStageNeed_2 <= accessCountQueue_deq_bits_2;
        reorderStageNeed_3 <= accessCountQueue_deq_bits_3;
      end
      if (waiteStageEnqFire) begin
        waiteReadDataPipeReg_executeGroup <= readWaitQueue_deq_bits_executeGroup;
        waiteReadDataPipeReg_sourceValid <= readWaitQueue_deq_bits_sourceValid;
        waiteReadDataPipeReg_replaceVs1 <= readWaitQueue_deq_bits_replaceVs1;
        waiteReadDataPipeReg_needRead <= readWaitQueue_deq_bits_needRead;
        waiteReadDataPipeReg_last <= readWaitQueue_deq_bits_last;
      end
      if (readTokenRelease_1)
        waiteReadData_1 <= readData_readDataQueue_1_deq_bits;
      if (readTokenRelease_2)
        waiteReadData_2 <= readData_readDataQueue_2_deq_bits;
      if (readTokenRelease_3)
        waiteReadData_3 <= readData_readDataQueue_3_deq_bits;
      if (waiteStageEnqFire & (|readResultValid))
        waiteReadSate <= readResultValid;
      else if (|readResultValid)
        waiteReadSate <= waiteReadSate | readResultValid;
      else if (waiteStageEnqFire)
        waiteReadSate <= 4'h0;
      if (waiteStageDeqFire ^ waiteStageEnqFire)
        waiteReadStageValid <= waiteStageEnqFire;
      if (_dataNotInShifter_T ^ writeRelease_0)
        dataNotInShifter_writeTokenCounter <= dataNotInShifter_writeTokenCounter + dataNotInShifter_writeTokenChange;
      if (_dataNotInShifter_T_3 ^ writeRelease_1)
        dataNotInShifter_writeTokenCounter_1 <= dataNotInShifter_writeTokenCounter_1 + dataNotInShifter_writeTokenChange_1;
      if (_dataNotInShifter_T_6 ^ writeRelease_2)
        dataNotInShifter_writeTokenCounter_2 <= dataNotInShifter_writeTokenCounter_2 + dataNotInShifter_writeTokenChange_2;
      if (_dataNotInShifter_T_9 ^ writeRelease_3)
        dataNotInShifter_writeTokenCounter_3 <= dataNotInShifter_writeTokenCounter_3 + dataNotInShifter_writeTokenChange_3;
      waiteLastRequest <= ~readType & requestStageDeq & lastGroup | ~lastReportValid & waiteLastRequest;
      waitQueueClear <= executeStageClean | invalidEnq | ~lastReportValid & waitQueueClear;
    end
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:31];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [5:0] i = 6'h0; i < 6'h20; i += 6'h1) begin
          _RANDOM[i[4:0]] = `RANDOM;
        end
        v0_0 = _RANDOM[5'h0];
        v0_1 = _RANDOM[5'h1];
        v0_2 = _RANDOM[5'h2];
        v0_3 = _RANDOM[5'h3];
        v0_4 = _RANDOM[5'h4];
        v0_5 = _RANDOM[5'h5];
        v0_6 = _RANDOM[5'h6];
        v0_7 = _RANDOM[5'h7];
        gatherReadState = _RANDOM[5'h8][1:0];
        gatherDatOffset = _RANDOM[5'h8][3:2];
        gatherLane = _RANDOM[5'h8][5:4];
        gatherOffset = _RANDOM[5'h8][6];
        gatherGrowth = _RANDOM[5'h8][9:7];
        instReg_instructionIndex = _RANDOM[5'h8][12:10];
        instReg_decodeResult_specialSlot = _RANDOM[5'h8][13];
        instReg_decodeResult_topUop = _RANDOM[5'h8][18:14];
        instReg_decodeResult_popCount = _RANDOM[5'h8][19];
        instReg_decodeResult_ffo = _RANDOM[5'h8][20];
        instReg_decodeResult_average = _RANDOM[5'h8][21];
        instReg_decodeResult_reverse = _RANDOM[5'h8][22];
        instReg_decodeResult_dontNeedExecuteInLane = _RANDOM[5'h8][23];
        instReg_decodeResult_scheduler = _RANDOM[5'h8][24];
        instReg_decodeResult_sReadVD = _RANDOM[5'h8][25];
        instReg_decodeResult_vtype = _RANDOM[5'h8][26];
        instReg_decodeResult_sWrite = _RANDOM[5'h8][27];
        instReg_decodeResult_crossRead = _RANDOM[5'h8][28];
        instReg_decodeResult_crossWrite = _RANDOM[5'h8][29];
        instReg_decodeResult_maskUnit = _RANDOM[5'h8][30];
        instReg_decodeResult_special = _RANDOM[5'h8][31];
        instReg_decodeResult_saturate = _RANDOM[5'h9][0];
        instReg_decodeResult_vwmacc = _RANDOM[5'h9][1];
        instReg_decodeResult_readOnly = _RANDOM[5'h9][2];
        instReg_decodeResult_maskSource = _RANDOM[5'h9][3];
        instReg_decodeResult_maskDestination = _RANDOM[5'h9][4];
        instReg_decodeResult_maskLogic = _RANDOM[5'h9][5];
        instReg_decodeResult_uop = _RANDOM[5'h9][9:6];
        instReg_decodeResult_iota = _RANDOM[5'h9][10];
        instReg_decodeResult_mv = _RANDOM[5'h9][11];
        instReg_decodeResult_extend = _RANDOM[5'h9][12];
        instReg_decodeResult_unOrderWrite = _RANDOM[5'h9][13];
        instReg_decodeResult_compress = _RANDOM[5'h9][14];
        instReg_decodeResult_gather16 = _RANDOM[5'h9][15];
        instReg_decodeResult_gather = _RANDOM[5'h9][16];
        instReg_decodeResult_slid = _RANDOM[5'h9][17];
        instReg_decodeResult_targetRd = _RANDOM[5'h9][18];
        instReg_decodeResult_widenReduce = _RANDOM[5'h9][19];
        instReg_decodeResult_red = _RANDOM[5'h9][20];
        instReg_decodeResult_nr = _RANDOM[5'h9][21];
        instReg_decodeResult_itype = _RANDOM[5'h9][22];
        instReg_decodeResult_unsigned1 = _RANDOM[5'h9][23];
        instReg_decodeResult_unsigned0 = _RANDOM[5'h9][24];
        instReg_decodeResult_other = _RANDOM[5'h9][25];
        instReg_decodeResult_multiCycle = _RANDOM[5'h9][26];
        instReg_decodeResult_divider = _RANDOM[5'h9][27];
        instReg_decodeResult_multiplier = _RANDOM[5'h9][28];
        instReg_decodeResult_shift = _RANDOM[5'h9][29];
        instReg_decodeResult_adder = _RANDOM[5'h9][30];
        instReg_decodeResult_logic = _RANDOM[5'h9][31];
        instReg_readFromScala = _RANDOM[5'hA];
        instReg_sew = _RANDOM[5'hB][1:0];
        instReg_vlmul = _RANDOM[5'hB][4:2];
        instReg_maskType = _RANDOM[5'hB][5];
        instReg_vxrm = _RANDOM[5'hB][8:6];
        instReg_vs2 = _RANDOM[5'hB][13:9];
        instReg_vs1 = _RANDOM[5'hB][18:14];
        instReg_vd = _RANDOM[5'hB][23:19];
        instReg_vl = {_RANDOM[5'hB][31:24], _RANDOM[5'hC][0]};
        instVlValid = _RANDOM[5'hC][1];
        readVS1Reg_dataValid = _RANDOM[5'hC][2];
        readVS1Reg_requestSend = _RANDOM[5'hC][3];
        readVS1Reg_sendToExecution = _RANDOM[5'hC][4];
        readVS1Reg_data = {_RANDOM[5'hC][31:5], _RANDOM[5'hD][4:0]};
        readVS1Reg_readIndex = _RANDOM[5'hD][8:5];
        exeReqReg_0_valid = _RANDOM[5'hD][13];
        exeReqReg_0_bits_source1 = {_RANDOM[5'hD][31:14], _RANDOM[5'hE][13:0]};
        exeReqReg_0_bits_source2 = {_RANDOM[5'hE][31:14], _RANDOM[5'hF][13:0]};
        exeReqReg_0_bits_index = _RANDOM[5'hF][16:14];
        exeReqReg_0_bits_ffo = _RANDOM[5'hF][17];
        exeReqReg_1_valid = _RANDOM[5'hF][18];
        exeReqReg_1_bits_source1 = {_RANDOM[5'hF][31:19], _RANDOM[5'h10][18:0]};
        exeReqReg_1_bits_source2 = {_RANDOM[5'h10][31:19], _RANDOM[5'h11][18:0]};
        exeReqReg_1_bits_index = _RANDOM[5'h11][21:19];
        exeReqReg_1_bits_ffo = _RANDOM[5'h11][22];
        exeReqReg_2_valid = _RANDOM[5'h11][23];
        exeReqReg_2_bits_source1 = {_RANDOM[5'h11][31:24], _RANDOM[5'h12][23:0]};
        exeReqReg_2_bits_source2 = {_RANDOM[5'h12][31:24], _RANDOM[5'h13][23:0]};
        exeReqReg_2_bits_index = _RANDOM[5'h13][26:24];
        exeReqReg_2_bits_ffo = _RANDOM[5'h13][27];
        exeReqReg_3_valid = _RANDOM[5'h13][28];
        exeReqReg_3_bits_source1 = {_RANDOM[5'h13][31:29], _RANDOM[5'h14][28:0]};
        exeReqReg_3_bits_source2 = {_RANDOM[5'h14][31:29], _RANDOM[5'h15][28:0]};
        exeReqReg_3_bits_index = _RANDOM[5'h15][31:29];
        exeReqReg_3_bits_ffo = _RANDOM[5'h16][0];
        requestCounter = _RANDOM[5'h16][5:1];
        executeIndex = _RANDOM[5'h16][7:6];
        readIssueStageState_groupReadState = _RANDOM[5'h16][11:8];
        readIssueStageState_needRead = _RANDOM[5'h16][15:12];
        readIssueStageState_elementValid = _RANDOM[5'h16][19:16];
        readIssueStageState_replaceVs1 = _RANDOM[5'h16][23:20];
        readIssueStageState_readOffset = _RANDOM[5'h16][27:24];
        readIssueStageState_accessLane_0 = _RANDOM[5'h16][29:28];
        readIssueStageState_accessLane_1 = _RANDOM[5'h16][31:30];
        readIssueStageState_accessLane_2 = _RANDOM[5'h17][1:0];
        readIssueStageState_accessLane_3 = _RANDOM[5'h17][3:2];
        readIssueStageState_vsGrowth_0 = _RANDOM[5'h17][6:4];
        readIssueStageState_vsGrowth_1 = _RANDOM[5'h17][9:7];
        readIssueStageState_vsGrowth_2 = _RANDOM[5'h17][12:10];
        readIssueStageState_vsGrowth_3 = _RANDOM[5'h17][15:13];
        readIssueStageState_executeGroup = _RANDOM[5'h17][22:16];
        readIssueStageState_readDataOffset = _RANDOM[5'h17][30:23];
        readIssueStageState_last = _RANDOM[5'h17][31];
        readIssueStageValid = _RANDOM[5'h18][0];
        tokenCheck_counter = _RANDOM[5'h18][4:1];
        tokenCheck_counter_1 = _RANDOM[5'h18][8:5];
        tokenCheck_counter_2 = _RANDOM[5'h18][12:9];
        tokenCheck_counter_3 = _RANDOM[5'h18][16:13];
        reorderQueueAllocate_counter = _RANDOM[5'h18][20:17];
        reorderQueueAllocate_counterWillUpdate = _RANDOM[5'h18][24:21];
        reorderQueueAllocate_counter_1 = _RANDOM[5'h18][28:25];
        reorderQueueAllocate_counterWillUpdate_1 = {_RANDOM[5'h18][31:29], _RANDOM[5'h19][0]};
        reorderQueueAllocate_counter_2 = _RANDOM[5'h19][4:1];
        reorderQueueAllocate_counterWillUpdate_2 = _RANDOM[5'h19][8:5];
        reorderQueueAllocate_counter_3 = _RANDOM[5'h19][12:9];
        reorderQueueAllocate_counterWillUpdate_3 = _RANDOM[5'h19][16:13];
        reorderStageValid = _RANDOM[5'h19][17];
        reorderStageState_0 = _RANDOM[5'h19][20:18];
        reorderStageState_1 = _RANDOM[5'h19][23:21];
        reorderStageState_2 = _RANDOM[5'h19][26:24];
        reorderStageState_3 = _RANDOM[5'h19][29:27];
        reorderStageNeed_0 = {_RANDOM[5'h19][31:30], _RANDOM[5'h1A][0]};
        reorderStageNeed_1 = _RANDOM[5'h1A][3:1];
        reorderStageNeed_2 = _RANDOM[5'h1A][6:4];
        reorderStageNeed_3 = _RANDOM[5'h1A][9:7];
        waiteReadDataPipeReg_executeGroup = _RANDOM[5'h1A][16:10];
        waiteReadDataPipeReg_sourceValid = _RANDOM[5'h1A][20:17];
        waiteReadDataPipeReg_replaceVs1 = _RANDOM[5'h1A][24:21];
        waiteReadDataPipeReg_needRead = _RANDOM[5'h1A][28:25];
        waiteReadDataPipeReg_last = _RANDOM[5'h1A][29];
        waiteReadData_0 = {_RANDOM[5'h1A][31:30], _RANDOM[5'h1B][29:0]};
        waiteReadData_1 = {_RANDOM[5'h1B][31:30], _RANDOM[5'h1C][29:0]};
        waiteReadData_2 = {_RANDOM[5'h1C][31:30], _RANDOM[5'h1D][29:0]};
        waiteReadData_3 = {_RANDOM[5'h1D][31:30], _RANDOM[5'h1E][29:0]};
        waiteReadSate = {_RANDOM[5'h1E][31:30], _RANDOM[5'h1F][1:0]};
        waiteReadStageValid = _RANDOM[5'h1F][2];
        dataNotInShifter_writeTokenCounter = _RANDOM[5'h1F][5:3];
        dataNotInShifter_writeTokenCounter_1 = _RANDOM[5'h1F][8:6];
        dataNotInShifter_writeTokenCounter_2 = _RANDOM[5'h1F][11:9];
        dataNotInShifter_writeTokenCounter_3 = _RANDOM[5'h1F][14:12];
        waiteLastRequest = _RANDOM[5'h1F][15];
        waitQueueClear = _RANDOM[5'h1F][16];
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  wire              exeRequestQueue_0_empty;
  assign exeRequestQueue_0_empty = _exeRequestQueue_queue_fifo_empty;
  wire              exeRequestQueue_0_full;
  assign exeRequestQueue_0_full = _exeRequestQueue_queue_fifo_full;
  wire              exeRequestQueue_1_empty;
  assign exeRequestQueue_1_empty = _exeRequestQueue_queue_fifo_1_empty;
  wire              exeRequestQueue_1_full;
  assign exeRequestQueue_1_full = _exeRequestQueue_queue_fifo_1_full;
  wire              exeRequestQueue_2_empty;
  assign exeRequestQueue_2_empty = _exeRequestQueue_queue_fifo_2_empty;
  wire              exeRequestQueue_2_full;
  assign exeRequestQueue_2_full = _exeRequestQueue_queue_fifo_2_full;
  wire              exeRequestQueue_3_empty;
  assign exeRequestQueue_3_empty = _exeRequestQueue_queue_fifo_3_empty;
  wire              exeRequestQueue_3_full;
  assign exeRequestQueue_3_full = _exeRequestQueue_queue_fifo_3_full;
  wire              accessCountQueue_empty;
  assign accessCountQueue_empty = _accessCountQueue_fifo_empty;
  wire              accessCountQueue_full;
  assign accessCountQueue_full = _accessCountQueue_fifo_full;
  wire              readWaitQueue_empty;
  assign readWaitQueue_empty = _readWaitQueue_fifo_empty;
  wire              readWaitQueue_full;
  assign readWaitQueue_full = _readWaitQueue_fifo_full;
  assign compressUnitResultQueue_empty = _compressUnitResultQueue_fifo_empty;
  wire              compressUnitResultQueue_full;
  assign compressUnitResultQueue_full = _compressUnitResultQueue_fifo_full;
  wire              reorderQueueVec_0_empty;
  assign reorderQueueVec_0_empty = _reorderQueueVec_fifo_empty;
  wire              reorderQueueVec_0_full;
  assign reorderQueueVec_0_full = _reorderQueueVec_fifo_full;
  wire              reorderQueueVec_1_empty;
  assign reorderQueueVec_1_empty = _reorderQueueVec_fifo_1_empty;
  wire              reorderQueueVec_1_full;
  assign reorderQueueVec_1_full = _reorderQueueVec_fifo_1_full;
  wire              reorderQueueVec_2_empty;
  assign reorderQueueVec_2_empty = _reorderQueueVec_fifo_2_empty;
  wire              reorderQueueVec_2_full;
  assign reorderQueueVec_2_full = _reorderQueueVec_fifo_2_full;
  wire              reorderQueueVec_3_empty;
  assign reorderQueueVec_3_empty = _reorderQueueVec_fifo_3_empty;
  wire              reorderQueueVec_3_full;
  assign reorderQueueVec_3_full = _reorderQueueVec_fifo_3_full;
  wire              readMessageQueue_empty;
  assign readMessageQueue_empty = _readMessageQueue_fifo_empty;
  wire              readMessageQueue_full;
  assign readMessageQueue_full = _readMessageQueue_fifo_full;
  wire              readMessageQueue_1_empty;
  assign readMessageQueue_1_empty = _readMessageQueue_fifo_1_empty;
  wire              readMessageQueue_1_full;
  assign readMessageQueue_1_full = _readMessageQueue_fifo_1_full;
  wire              readMessageQueue_2_empty;
  assign readMessageQueue_2_empty = _readMessageQueue_fifo_2_empty;
  wire              readMessageQueue_2_full;
  assign readMessageQueue_2_full = _readMessageQueue_fifo_2_full;
  wire              readMessageQueue_3_empty;
  assign readMessageQueue_3_empty = _readMessageQueue_fifo_3_empty;
  wire              readMessageQueue_3_full;
  assign readMessageQueue_3_full = _readMessageQueue_fifo_3_full;
  wire              readData_readDataQueue_empty;
  assign readData_readDataQueue_empty = _readData_readDataQueue_fifo_empty;
  wire              readData_readDataQueue_full;
  assign readData_readDataQueue_full = _readData_readDataQueue_fifo_full;
  wire              readData_readDataQueue_1_empty;
  assign readData_readDataQueue_1_empty = _readData_readDataQueue_fifo_1_empty;
  wire              readData_readDataQueue_1_full;
  assign readData_readDataQueue_1_full = _readData_readDataQueue_fifo_1_full;
  wire              readData_readDataQueue_2_empty;
  assign readData_readDataQueue_2_empty = _readData_readDataQueue_fifo_2_empty;
  wire              readData_readDataQueue_2_full;
  assign readData_readDataQueue_2_full = _readData_readDataQueue_fifo_2_full;
  wire              readData_readDataQueue_3_empty;
  assign readData_readDataQueue_3_empty = _readData_readDataQueue_fifo_3_empty;
  wire              readData_readDataQueue_3_full;
  assign readData_readDataQueue_3_full = _readData_readDataQueue_fifo_3_full;
  assign compressUnitResultQueue_enq_valid = _compressUnit_out_compressValid;
  assign compressUnitResultQueue_enq_bits_compressValid = _compressUnit_out_compressValid;
  wire              writeQueue_0_empty;
  assign writeQueue_0_empty = _writeQueue_fifo_empty;
  wire              writeQueue_0_full;
  assign writeQueue_0_full = _writeQueue_fifo_full;
  wire              writeQueue_1_empty;
  assign writeQueue_1_empty = _writeQueue_fifo_1_empty;
  wire              writeQueue_1_full;
  assign writeQueue_1_full = _writeQueue_fifo_1_full;
  wire              writeQueue_2_empty;
  assign writeQueue_2_empty = _writeQueue_fifo_2_empty;
  wire              writeQueue_2_full;
  assign writeQueue_2_full = _writeQueue_fifo_2_full;
  wire              writeQueue_3_empty;
  assign writeQueue_3_empty = _writeQueue_fifo_3_empty;
  wire              writeQueue_3_full;
  assign writeQueue_3_full = _writeQueue_fifo_3_full;
  BitLevelMaskWrite maskedWrite (
    .clock                             (clock),
    .reset                             (reset),
    .needWAR                           (maskDestinationType),
    .vd                                (instReg_vd),
    .in_0_ready                        (_maskedWrite_in_0_ready),
    .in_0_valid                        (unitType[2] ? _reduceUnit_out_valid : executeValid & maskFilter),
    .in_0_bits_data                    (unitType[2] ? _reduceUnit_out_bits_data : executeResult[31:0]),
    .in_0_bits_bitMask                 (currentMaskGroupForDestination[31:0]),
    .in_0_bits_mask                    (unitType[2] ? _reduceUnit_out_bits_mask : executeWriteByteMask[3:0]),
    .in_0_bits_groupCounter            (unitType[2] ? 5'h0 : executeDeqGroupCounter[4:0]),
    .in_0_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[0] & ffo),
    .in_1_ready                        (_maskedWrite_in_1_ready),
    .in_1_valid                        (executeValid & maskFilter_1),
    .in_1_bits_data                    (executeResult[63:32]),
    .in_1_bits_bitMask                 (currentMaskGroupForDestination[63:32]),
    .in_1_bits_mask                    (executeWriteByteMask[7:4]),
    .in_1_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_1_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[1] & ffo),
    .in_2_ready                        (_maskedWrite_in_2_ready),
    .in_2_valid                        (executeValid & maskFilter_2),
    .in_2_bits_data                    (executeResult[95:64]),
    .in_2_bits_bitMask                 (currentMaskGroupForDestination[95:64]),
    .in_2_bits_mask                    (executeWriteByteMask[11:8]),
    .in_2_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_2_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[2] & ffo),
    .in_3_ready                        (_maskedWrite_in_3_ready),
    .in_3_valid                        (executeValid & maskFilter_3),
    .in_3_bits_data                    (executeResult[127:96]),
    .in_3_bits_bitMask                 (currentMaskGroupForDestination[127:96]),
    .in_3_bits_mask                    (executeWriteByteMask[15:12]),
    .in_3_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_3_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[3] & ffo),
    .out_0_ready                       (writeQueue_0_enq_ready),
    .out_0_valid                       (_maskedWrite_out_0_valid),
    .out_0_bits_ffoByOther             (_maskedWrite_out_0_bits_ffoByOther),
    .out_0_bits_writeData_data         (_maskedWrite_out_0_bits_writeData_data),
    .out_0_bits_writeData_mask         (_maskedWrite_out_0_bits_writeData_mask),
    .out_0_bits_writeData_groupCounter (_maskedWrite_out_0_bits_writeData_groupCounter),
    .out_1_ready                       (writeQueue_1_enq_ready),
    .out_1_valid                       (_maskedWrite_out_1_valid),
    .out_1_bits_ffoByOther             (_maskedWrite_out_1_bits_ffoByOther),
    .out_1_bits_writeData_data         (_maskedWrite_out_1_bits_writeData_data),
    .out_1_bits_writeData_mask         (_maskedWrite_out_1_bits_writeData_mask),
    .out_1_bits_writeData_groupCounter (_maskedWrite_out_1_bits_writeData_groupCounter),
    .out_2_ready                       (writeQueue_2_enq_ready),
    .out_2_valid                       (_maskedWrite_out_2_valid),
    .out_2_bits_ffoByOther             (_maskedWrite_out_2_bits_ffoByOther),
    .out_2_bits_writeData_data         (_maskedWrite_out_2_bits_writeData_data),
    .out_2_bits_writeData_mask         (_maskedWrite_out_2_bits_writeData_mask),
    .out_2_bits_writeData_groupCounter (_maskedWrite_out_2_bits_writeData_groupCounter),
    .out_3_ready                       (writeQueue_3_enq_ready),
    .out_3_valid                       (_maskedWrite_out_3_valid),
    .out_3_bits_ffoByOther             (_maskedWrite_out_3_bits_ffoByOther),
    .out_3_bits_writeData_data         (_maskedWrite_out_3_bits_writeData_data),
    .out_3_bits_writeData_mask         (_maskedWrite_out_3_bits_writeData_mask),
    .out_3_bits_writeData_groupCounter (_maskedWrite_out_3_bits_writeData_groupCounter),
    .readChannel_0_ready               (readChannel_0_ready_0),
    .readChannel_0_valid               (_maskedWrite_readChannel_0_valid),
    .readChannel_0_bits_vs             (_maskedWrite_readChannel_0_bits_vs),
    .readChannel_0_bits_offset         (_maskedWrite_readChannel_0_bits_offset),
    .readChannel_1_ready               (readChannel_1_ready_0),
    .readChannel_1_valid               (_maskedWrite_readChannel_1_valid),
    .readChannel_1_bits_vs             (_maskedWrite_readChannel_1_bits_vs),
    .readChannel_1_bits_offset         (_maskedWrite_readChannel_1_bits_offset),
    .readChannel_2_ready               (readChannel_2_ready_0),
    .readChannel_2_valid               (_maskedWrite_readChannel_2_valid),
    .readChannel_2_bits_vs             (_maskedWrite_readChannel_2_bits_vs),
    .readChannel_2_bits_offset         (_maskedWrite_readChannel_2_bits_offset),
    .readChannel_3_ready               (readChannel_3_ready_0),
    .readChannel_3_valid               (_maskedWrite_readChannel_3_valid),
    .readChannel_3_bits_vs             (_maskedWrite_readChannel_3_bits_vs),
    .readChannel_3_bits_offset         (_maskedWrite_readChannel_3_bits_offset),
    .readResult_0_valid                (readResult_0_valid),
    .readResult_0_bits                 (readResult_0_bits),
    .readResult_1_valid                (readResult_1_valid),
    .readResult_1_bits                 (readResult_1_bits),
    .readResult_2_valid                (readResult_2_valid),
    .readResult_2_bits                 (readResult_2_bits),
    .readResult_3_valid                (readResult_3_valid),
    .readResult_3_bits                 (readResult_3_bits),
    .stageClear                        (_maskedWrite_stageClear)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_0_enq_ready & exeRequestQueue_0_enq_valid & ~(_exeRequestQueue_queue_fifo_empty & exeRequestQueue_0_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_0_deq_ready & ~_exeRequestQueue_queue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn),
    .empty        (_exeRequestQueue_queue_fifo_empty),
    .almost_empty (exeRequestQueue_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_0_almostFull),
    .full         (_exeRequestQueue_queue_fifo_full),
    .error        (_exeRequestQueue_queue_fifo_error),
    .data_out     (_exeRequestQueue_queue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_1_enq_ready & exeRequestQueue_1_enq_valid & ~(_exeRequestQueue_queue_fifo_1_empty & exeRequestQueue_1_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_1_deq_ready & ~_exeRequestQueue_queue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_1),
    .empty        (_exeRequestQueue_queue_fifo_1_empty),
    .almost_empty (exeRequestQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_1_almostFull),
    .full         (_exeRequestQueue_queue_fifo_1_full),
    .error        (_exeRequestQueue_queue_fifo_1_error),
    .data_out     (_exeRequestQueue_queue_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_2_enq_ready & exeRequestQueue_2_enq_valid & ~(_exeRequestQueue_queue_fifo_2_empty & exeRequestQueue_2_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_2_deq_ready & ~_exeRequestQueue_queue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_2),
    .empty        (_exeRequestQueue_queue_fifo_2_empty),
    .almost_empty (exeRequestQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_2_almostFull),
    .full         (_exeRequestQueue_queue_fifo_2_full),
    .error        (_exeRequestQueue_queue_fifo_2_error),
    .data_out     (_exeRequestQueue_queue_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_3_enq_ready & exeRequestQueue_3_enq_valid & ~(_exeRequestQueue_queue_fifo_3_empty & exeRequestQueue_3_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_3_deq_ready & ~_exeRequestQueue_queue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_3),
    .empty        (_exeRequestQueue_queue_fifo_3_empty),
    .almost_empty (exeRequestQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_3_almostFull),
    .full         (_exeRequestQueue_queue_fifo_3_full),
    .error        (_exeRequestQueue_queue_fifo_3_error),
    .data_out     (_exeRequestQueue_queue_fifo_3_data_out)
  );
  SlideIndexGen slideAddressGen (
    .clock                              (clock),
    .reset                              (reset),
    .newInstruction                     (instReq_valid & (|instReq_bits_vl)),
    .instructionReq_decodeResult_topUop (instReg_decodeResult_topUop),
    .instructionReq_readFromScala       (instReg_readFromScala),
    .instructionReq_sew                 (instReg_sew),
    .instructionReq_vlmul               (instReg_vlmul),
    .instructionReq_maskType            (instReg_maskType),
    .instructionReq_vl                  (instReg_vl),
    .indexDeq_ready                     (slideAddressGen_indexDeq_ready),
    .indexDeq_valid                     (_slideAddressGen_indexDeq_valid),
    .indexDeq_bits_needRead             (_slideAddressGen_indexDeq_bits_needRead),
    .indexDeq_bits_elementValid         (_slideAddressGen_indexDeq_bits_elementValid),
    .indexDeq_bits_replaceVs1           (_slideAddressGen_indexDeq_bits_replaceVs1),
    .indexDeq_bits_readOffset           (_slideAddressGen_indexDeq_bits_readOffset),
    .indexDeq_bits_accessLane_0         (_slideAddressGen_indexDeq_bits_accessLane_0),
    .indexDeq_bits_accessLane_1         (_slideAddressGen_indexDeq_bits_accessLane_1),
    .indexDeq_bits_accessLane_2         (_slideAddressGen_indexDeq_bits_accessLane_2),
    .indexDeq_bits_accessLane_3         (_slideAddressGen_indexDeq_bits_accessLane_3),
    .indexDeq_bits_vsGrowth_0           (_slideAddressGen_indexDeq_bits_vsGrowth_0),
    .indexDeq_bits_vsGrowth_1           (_slideAddressGen_indexDeq_bits_vsGrowth_1),
    .indexDeq_bits_vsGrowth_2           (_slideAddressGen_indexDeq_bits_vsGrowth_2),
    .indexDeq_bits_vsGrowth_3           (_slideAddressGen_indexDeq_bits_vsGrowth_3),
    .indexDeq_bits_executeGroup         (_slideAddressGen_indexDeq_bits_executeGroup),
    .indexDeq_bits_readDataOffset       (_slideAddressGen_indexDeq_bits_readDataOffset),
    .indexDeq_bits_last                 (_slideAddressGen_indexDeq_bits_last),
    .slideGroupOut                      (_slideAddressGen_slideGroupOut),
    .slideMaskInput                     (_GEN_12[_slideAddressGen_slideGroupOut[5:0]])
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) accessCountQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(accessCountQueue_enq_ready & accessCountQueue_enq_valid)),
    .pop_req_n    (~(accessCountQueue_deq_ready & ~_accessCountQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (accessCountQueue_dataIn),
    .empty        (_accessCountQueue_fifo_empty),
    .almost_empty (accessCountQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (accessCountQueue_almostFull),
    .full         (_accessCountQueue_fifo_full),
    .error        (_accessCountQueue_fifo_error),
    .data_out     (_accessCountQueue_fifo_data_out)
  );
  MaskUnitReadCrossBar readCrossBar (
    .input_0_ready            (_readCrossBar_input_0_ready),
    .input_0_valid            (readCrossBar_input_0_valid),
    .input_0_bits_vs          (selectExecuteReq_0_bits_vs),
    .input_0_bits_offset      (selectExecuteReq_0_bits_offset),
    .input_0_bits_readLane    (selectExecuteReq_0_bits_readLane),
    .input_0_bits_dataOffset  (selectExecuteReq_0_bits_dataOffset),
    .input_1_ready            (_readCrossBar_input_1_ready),
    .input_1_valid            (readCrossBar_input_1_valid),
    .input_1_bits_vs          (selectExecuteReq_1_bits_vs),
    .input_1_bits_offset      (selectExecuteReq_1_bits_offset),
    .input_1_bits_readLane    (selectExecuteReq_1_bits_readLane),
    .input_1_bits_dataOffset  (selectExecuteReq_1_bits_dataOffset),
    .input_2_ready            (_readCrossBar_input_2_ready),
    .input_2_valid            (readCrossBar_input_2_valid),
    .input_2_bits_vs          (selectExecuteReq_2_bits_vs),
    .input_2_bits_offset      (selectExecuteReq_2_bits_offset),
    .input_2_bits_readLane    (selectExecuteReq_2_bits_readLane),
    .input_2_bits_dataOffset  (selectExecuteReq_2_bits_dataOffset),
    .input_3_ready            (_readCrossBar_input_3_ready),
    .input_3_valid            (readCrossBar_input_3_valid),
    .input_3_bits_vs          (selectExecuteReq_3_bits_vs),
    .input_3_bits_offset      (selectExecuteReq_3_bits_offset),
    .input_3_bits_readLane    (selectExecuteReq_3_bits_readLane),
    .input_3_bits_dataOffset  (selectExecuteReq_3_bits_dataOffset),
    .output_0_ready           (readChannel_0_ready_0 & readMessageQueue_enq_ready),
    .output_0_valid           (_readCrossBar_output_0_valid),
    .output_0_bits_vs         (_readCrossBar_output_0_bits_vs),
    .output_0_bits_offset     (_readCrossBar_output_0_bits_offset),
    .output_0_bits_writeIndex (_readCrossBar_output_0_bits_writeIndex),
    .output_0_bits_dataOffset (readMessageQueue_enq_bits_dataOffset),
    .output_1_ready           (readChannel_1_ready_0 & readMessageQueue_1_enq_ready),
    .output_1_valid           (_readCrossBar_output_1_valid),
    .output_1_bits_vs         (_readCrossBar_output_1_bits_vs),
    .output_1_bits_offset     (_readCrossBar_output_1_bits_offset),
    .output_1_bits_writeIndex (_readCrossBar_output_1_bits_writeIndex),
    .output_1_bits_dataOffset (readMessageQueue_1_enq_bits_dataOffset),
    .output_2_ready           (readChannel_2_ready_0 & readMessageQueue_2_enq_ready),
    .output_2_valid           (_readCrossBar_output_2_valid),
    .output_2_bits_vs         (_readCrossBar_output_2_bits_vs),
    .output_2_bits_offset     (_readCrossBar_output_2_bits_offset),
    .output_2_bits_writeIndex (_readCrossBar_output_2_bits_writeIndex),
    .output_2_bits_dataOffset (readMessageQueue_2_enq_bits_dataOffset),
    .output_3_ready           (readChannel_3_ready_0 & readMessageQueue_3_enq_ready),
    .output_3_valid           (_readCrossBar_output_3_valid),
    .output_3_bits_vs         (_readCrossBar_output_3_bits_vs),
    .output_3_bits_offset     (_readCrossBar_output_3_bits_offset),
    .output_3_bits_writeIndex (_readCrossBar_output_3_bits_writeIndex),
    .output_3_bits_dataOffset (readMessageQueue_3_enq_bits_dataOffset)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(20)
  ) readWaitQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readWaitQueue_enq_ready & readWaitQueue_enq_valid)),
    .pop_req_n    (~(readWaitQueue_deq_ready & ~_readWaitQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (readWaitQueue_dataIn),
    .empty        (_readWaitQueue_fifo_empty),
    .almost_empty (readWaitQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readWaitQueue_almostFull),
    .full         (_readWaitQueue_fifo_full),
    .error        (_readWaitQueue_fifo_error),
    .data_out     (_readWaitQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(154)
  ) compressUnitResultQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(compressUnitResultQueue_enq_ready & compressUnitResultQueue_enq_valid & ~(_compressUnitResultQueue_fifo_empty & compressUnitResultQueue_deq_ready))),
    .pop_req_n    (~(compressUnitResultQueue_deq_ready & ~_compressUnitResultQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (compressUnitResultQueue_dataIn),
    .empty        (_compressUnitResultQueue_fifo_empty),
    .almost_empty (compressUnitResultQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (compressUnitResultQueue_almostFull),
    .full         (_compressUnitResultQueue_fifo_full),
    .error        (_compressUnitResultQueue_fifo_error),
    .data_out     (_compressUnitResultQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(36)
  ) reorderQueueVec_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_0_enq_ready & reorderQueueVec_0_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_0_deq_ready & ~_reorderQueueVec_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn),
    .empty        (_reorderQueueVec_fifo_empty),
    .almost_empty (reorderQueueVec_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_0_almostFull),
    .full         (_reorderQueueVec_fifo_full),
    .error        (_reorderQueueVec_fifo_error),
    .data_out     (_reorderQueueVec_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(36)
  ) reorderQueueVec_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_1_enq_ready & reorderQueueVec_1_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_1_deq_ready & ~_reorderQueueVec_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_1),
    .empty        (_reorderQueueVec_fifo_1_empty),
    .almost_empty (reorderQueueVec_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_1_almostFull),
    .full         (_reorderQueueVec_fifo_1_full),
    .error        (_reorderQueueVec_fifo_1_error),
    .data_out     (_reorderQueueVec_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(36)
  ) reorderQueueVec_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_2_enq_ready & reorderQueueVec_2_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_2_deq_ready & ~_reorderQueueVec_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_2),
    .empty        (_reorderQueueVec_fifo_2_empty),
    .almost_empty (reorderQueueVec_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_2_almostFull),
    .full         (_reorderQueueVec_fifo_2_full),
    .error        (_reorderQueueVec_fifo_2_error),
    .data_out     (_reorderQueueVec_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(36)
  ) reorderQueueVec_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_3_enq_ready & reorderQueueVec_3_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_3_deq_ready & ~_reorderQueueVec_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_3),
    .empty        (_reorderQueueVec_fifo_3_empty),
    .almost_empty (reorderQueueVec_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_3_almostFull),
    .full         (_reorderQueueVec_fifo_3_full),
    .error        (_reorderQueueVec_fifo_3_error),
    .data_out     (_reorderQueueVec_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(6)
  ) readMessageQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_enq_ready & readMessageQueue_enq_valid)),
    .pop_req_n    (~(readMessageQueue_deq_ready & ~_readMessageQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn),
    .empty        (_readMessageQueue_fifo_empty),
    .almost_empty (readMessageQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_almostFull),
    .full         (_readMessageQueue_fifo_full),
    .error        (_readMessageQueue_fifo_error),
    .data_out     (_readMessageQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(6)
  ) readMessageQueue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_1_enq_ready & readMessageQueue_1_enq_valid)),
    .pop_req_n    (~(readMessageQueue_1_deq_ready & ~_readMessageQueue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_1),
    .empty        (_readMessageQueue_fifo_1_empty),
    .almost_empty (readMessageQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_1_almostFull),
    .full         (_readMessageQueue_fifo_1_full),
    .error        (_readMessageQueue_fifo_1_error),
    .data_out     (_readMessageQueue_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(6)
  ) readMessageQueue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_2_enq_ready & readMessageQueue_2_enq_valid)),
    .pop_req_n    (~(readMessageQueue_2_deq_ready & ~_readMessageQueue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_2),
    .empty        (_readMessageQueue_fifo_2_empty),
    .almost_empty (readMessageQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_2_almostFull),
    .full         (_readMessageQueue_fifo_2_full),
    .error        (_readMessageQueue_fifo_2_error),
    .data_out     (_readMessageQueue_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(6)
  ) readMessageQueue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_3_enq_ready & readMessageQueue_3_enq_valid)),
    .pop_req_n    (~(readMessageQueue_3_deq_ready & ~_readMessageQueue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_3),
    .empty        (_readMessageQueue_fifo_3_empty),
    .almost_empty (readMessageQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_3_almostFull),
    .full         (_readMessageQueue_fifo_3_full),
    .error        (_readMessageQueue_fifo_3_error),
    .data_out     (_readMessageQueue_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_enq_ready & readData_readDataQueue_enq_valid & ~(_readData_readDataQueue_fifo_empty & readData_readDataQueue_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_deq_ready & ~_readData_readDataQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_enq_bits),
    .empty        (_readData_readDataQueue_fifo_empty),
    .almost_empty (readData_readDataQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_almostFull),
    .full         (_readData_readDataQueue_fifo_full),
    .error        (_readData_readDataQueue_fifo_error),
    .data_out     (_readData_readDataQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_1_enq_ready & readData_readDataQueue_1_enq_valid & ~(_readData_readDataQueue_fifo_1_empty & readData_readDataQueue_1_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_1_deq_ready & ~_readData_readDataQueue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_1_enq_bits),
    .empty        (_readData_readDataQueue_fifo_1_empty),
    .almost_empty (readData_readDataQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_1_almostFull),
    .full         (_readData_readDataQueue_fifo_1_full),
    .error        (_readData_readDataQueue_fifo_1_error),
    .data_out     (_readData_readDataQueue_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_2_enq_ready & readData_readDataQueue_2_enq_valid & ~(_readData_readDataQueue_fifo_2_empty & readData_readDataQueue_2_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_2_deq_ready & ~_readData_readDataQueue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_2_enq_bits),
    .empty        (_readData_readDataQueue_fifo_2_empty),
    .almost_empty (readData_readDataQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_2_almostFull),
    .full         (_readData_readDataQueue_fifo_2_full),
    .error        (_readData_readDataQueue_fifo_2_error),
    .data_out     (_readData_readDataQueue_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_3_enq_ready & readData_readDataQueue_3_enq_valid & ~(_readData_readDataQueue_fifo_3_empty & readData_readDataQueue_3_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_3_deq_ready & ~_readData_readDataQueue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_3_enq_bits),
    .empty        (_readData_readDataQueue_fifo_3_empty),
    .almost_empty (readData_readDataQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_3_almostFull),
    .full         (_readData_readDataQueue_fifo_3_full),
    .error        (_readData_readDataQueue_fifo_3_error),
    .data_out     (_readData_readDataQueue_fifo_3_data_out)
  );
  MaskCompress compressUnit (
    .clock                  (clock),
    .reset                  (reset),
    .in_valid               (viotaCounterAdd),
    .in_bits_maskType       (instReg_maskType),
    .in_bits_eew            (instReg_sew),
    .in_bits_uop            (instReg_decodeResult_topUop[2:0]),
    .in_bits_readFromScalar (instReg_readFromScala),
    .in_bits_source1        (source1Select),
    .in_bits_mask           ({16'h0, executeElementMask}),
    .in_bits_source2        (source2),
    .in_bits_pipeData       (source1),
    .in_bits_groupCounter   (requestCounter),
    .in_bits_ffoInput       ({view__in_bits_ffoInput_hi, view__in_bits_ffoInput_lo}),
    .in_bits_validInput     ({view__in_bits_validInput_hi, view__in_bits_validInput_lo}),
    .in_bits_lastCompress   (lastGroup),
    .out_data               (compressUnitResultQueue_enq_bits_data),
    .out_mask               (compressUnitResultQueue_enq_bits_mask),
    .out_groupCounter       (compressUnitResultQueue_enq_bits_groupCounter),
    .out_ffoOutput          (compressUnitResultQueue_enq_bits_ffoOutput),
    .out_compressValid      (_compressUnit_out_compressValid),
    .newInstruction         (instReq_valid),
    .ffoInstruction         (&(instReq_bits_decodeResult_topUop[2:1])),
    .writeData              (_compressUnit_writeData),
    .stageValid             (_compressUnit_stageValid)
  );
  MaskReduce reduceUnit (
    .clock               (clock),
    .reset               (reset),
    .in_ready            (_reduceUnit_in_ready),
    .in_valid            (reduceUnit_in_valid),
    .in_bits_maskType    (instReg_maskType),
    .in_bits_eew         (instReg_sew),
    .in_bits_uop         (instReg_decodeResult_topUop[2:0]),
    .in_bits_readVS1     (readVS1Reg_data),
    .in_bits_source2     (source2),
    .in_bits_sourceValid ({view__in_bits_sourceValid_hi, view__in_bits_sourceValid_lo}),
    .in_bits_lastGroup   (lastGroup),
    .in_bits_vxrm        (instReg_vxrm),
    .in_bits_aluUop      (instReg_decodeResult_uop),
    .in_bits_sign        (~instReg_decodeResult_unsigned1),
    .out_valid           (_reduceUnit_out_valid),
    .out_bits_data       (_reduceUnit_out_bits_data),
    .out_bits_mask       (_reduceUnit_out_bits_mask),
    .firstGroup          (~readVS1Reg_sendToExecution & _view__firstGroup_T_1),
    .newInstruction      (instReq_valid),
    .validInst           (|instReg_vl),
    .pop                 (instReg_decodeResult_popCount)
  );
  MaskExtend extendUnit (
    .in_eew          (instReg_sew),
    .in_uop          (instReg_decodeResult_topUop[2:0]),
    .in_source2      (source2),
    .in_groupCounter (extendGroupCount[4:0]),
    .out             (_extendUnit_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_0_enq_ready & writeQueue_0_enq_valid)),
    .pop_req_n    (~(writeQueue_0_deq_ready & ~_writeQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn),
    .empty        (_writeQueue_fifo_empty),
    .almost_empty (writeQueue_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_0_almostFull),
    .full         (_writeQueue_fifo_full),
    .error        (_writeQueue_fifo_error),
    .data_out     (_writeQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_1_enq_ready & writeQueue_1_enq_valid)),
    .pop_req_n    (~(writeQueue_1_deq_ready & ~_writeQueue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_1),
    .empty        (_writeQueue_fifo_1_empty),
    .almost_empty (writeQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_1_almostFull),
    .full         (_writeQueue_fifo_1_full),
    .error        (_writeQueue_fifo_1_error),
    .data_out     (_writeQueue_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_2_enq_ready & writeQueue_2_enq_valid)),
    .pop_req_n    (~(writeQueue_2_deq_ready & ~_writeQueue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_2),
    .empty        (_writeQueue_fifo_2_empty),
    .almost_empty (writeQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_2_almostFull),
    .full         (_writeQueue_fifo_2_full),
    .error        (_writeQueue_fifo_2_error),
    .data_out     (_writeQueue_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_3_enq_ready & writeQueue_3_enq_valid)),
    .pop_req_n    (~(writeQueue_3_deq_ready & ~_writeQueue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_3),
    .empty        (_writeQueue_fifo_3_empty),
    .almost_empty (writeQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_3_almostFull),
    .full         (_writeQueue_fifo_3_full),
    .error        (_writeQueue_fifo_3_error),
    .data_out     (_writeQueue_fifo_3_data_out)
  );
  assign exeResp_0_valid = exeResp_0_valid_0;
  assign exeResp_0_bits_vd = exeResp_0_bits_vd_0;
  assign exeResp_0_bits_offset = exeResp_0_bits_offset_0;
  assign exeResp_0_bits_mask = exeResp_0_bits_mask_0;
  assign exeResp_0_bits_data = exeResp_0_bits_data_0;
  assign exeResp_0_bits_instructionIndex = exeResp_0_bits_instructionIndex_0;
  assign exeResp_1_valid = exeResp_1_valid_0;
  assign exeResp_1_bits_vd = exeResp_1_bits_vd_0;
  assign exeResp_1_bits_offset = exeResp_1_bits_offset_0;
  assign exeResp_1_bits_mask = exeResp_1_bits_mask_0;
  assign exeResp_1_bits_data = exeResp_1_bits_data_0;
  assign exeResp_1_bits_instructionIndex = exeResp_1_bits_instructionIndex_0;
  assign exeResp_2_valid = exeResp_2_valid_0;
  assign exeResp_2_bits_vd = exeResp_2_bits_vd_0;
  assign exeResp_2_bits_offset = exeResp_2_bits_offset_0;
  assign exeResp_2_bits_mask = exeResp_2_bits_mask_0;
  assign exeResp_2_bits_data = exeResp_2_bits_data_0;
  assign exeResp_2_bits_instructionIndex = exeResp_2_bits_instructionIndex_0;
  assign exeResp_3_valid = exeResp_3_valid_0;
  assign exeResp_3_bits_vd = exeResp_3_bits_vd_0;
  assign exeResp_3_bits_offset = exeResp_3_bits_offset_0;
  assign exeResp_3_bits_mask = exeResp_3_bits_mask_0;
  assign exeResp_3_bits_data = exeResp_3_bits_data_0;
  assign exeResp_3_bits_instructionIndex = exeResp_3_bits_instructionIndex_0;
  assign tokenIO_0_maskRequestRelease = tokenIO_0_maskRequestRelease_0;
  assign tokenIO_1_maskRequestRelease = tokenIO_1_maskRequestRelease_0;
  assign tokenIO_2_maskRequestRelease = tokenIO_2_maskRequestRelease_0;
  assign tokenIO_3_maskRequestRelease = tokenIO_3_maskRequestRelease_0;
  assign readChannel_0_valid = readChannel_0_valid_0;
  assign readChannel_0_bits_vs = readChannel_0_bits_vs_0;
  assign readChannel_0_bits_offset = readChannel_0_bits_offset_0;
  assign readChannel_0_bits_instructionIndex = readChannel_0_bits_instructionIndex_0;
  assign readChannel_1_valid = readChannel_1_valid_0;
  assign readChannel_1_bits_vs = readChannel_1_bits_vs_0;
  assign readChannel_1_bits_offset = readChannel_1_bits_offset_0;
  assign readChannel_1_bits_instructionIndex = readChannel_1_bits_instructionIndex_0;
  assign readChannel_2_valid = readChannel_2_valid_0;
  assign readChannel_2_bits_vs = readChannel_2_bits_vs_0;
  assign readChannel_2_bits_offset = readChannel_2_bits_offset_0;
  assign readChannel_2_bits_instructionIndex = readChannel_2_bits_instructionIndex_0;
  assign readChannel_3_valid = readChannel_3_valid_0;
  assign readChannel_3_bits_vs = readChannel_3_bits_vs_0;
  assign readChannel_3_bits_offset = readChannel_3_bits_offset_0;
  assign readChannel_3_bits_instructionIndex = readChannel_3_bits_instructionIndex_0;
  assign lastReport = _lastReport_output;
  assign laneMaskInput_0 = laneMaskSelect_0[0] ? v0SelectBySew[63:32] : v0SelectBySew[31:0];
  assign laneMaskInput_1 = laneMaskSelect_1[0] ? v0SelectBySew_1[63:32] : v0SelectBySew_1[31:0];
  assign laneMaskInput_2 = laneMaskSelect_2[0] ? v0SelectBySew_2[63:32] : v0SelectBySew_2[31:0];
  assign laneMaskInput_3 = laneMaskSelect_3[0] ? v0SelectBySew_3[63:32] : v0SelectBySew_3[31:0];
  assign writeRDData = instReg_decodeResult_popCount ? _reduceUnit_out_bits_data : _compressUnit_writeData;
  assign gatherData_valid = gatherData_valid_0;
  assign gatherData_bits = gatherData_bits_0;
endmodule

