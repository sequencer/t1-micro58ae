
// Include register initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for register randomization.

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_
module LSU(
  input          clock,
                 reset,
  output         request_ready,
  input          request_valid,
  input  [2:0]   request_bits_instructionInformation_nf,
  input          request_bits_instructionInformation_mew,
  input  [1:0]   request_bits_instructionInformation_mop,
  input  [4:0]   request_bits_instructionInformation_lumop,
  input  [1:0]   request_bits_instructionInformation_eew,
  input  [4:0]   request_bits_instructionInformation_vs3,
  input          request_bits_instructionInformation_isStore,
                 request_bits_instructionInformation_maskedLoadStore,
  input  [31:0]  request_bits_rs1Data,
                 request_bits_rs2Data,
  input  [2:0]   request_bits_instructionIndex,
  input          v0UpdateVec_0_valid,
  input  [31:0]  v0UpdateVec_0_bits_data,
  input  [8:0]   v0UpdateVec_0_bits_offset,
  input  [3:0]   v0UpdateVec_0_bits_mask,
  input          v0UpdateVec_1_valid,
  input  [31:0]  v0UpdateVec_1_bits_data,
  input  [8:0]   v0UpdateVec_1_bits_offset,
  input  [3:0]   v0UpdateVec_1_bits_mask,
  input          v0UpdateVec_2_valid,
  input  [31:0]  v0UpdateVec_2_bits_data,
  input  [8:0]   v0UpdateVec_2_bits_offset,
  input  [3:0]   v0UpdateVec_2_bits_mask,
  input          v0UpdateVec_3_valid,
  input  [31:0]  v0UpdateVec_3_bits_data,
  input  [8:0]   v0UpdateVec_3_bits_offset,
  input  [3:0]   v0UpdateVec_3_bits_mask,
  input          axi4Port_aw_ready,
  output         axi4Port_aw_valid,
  output [1:0]   axi4Port_aw_bits_id,
  output [31:0]  axi4Port_aw_bits_addr,
  input          axi4Port_w_ready,
  output         axi4Port_w_valid,
  output [127:0] axi4Port_w_bits_data,
  output [15:0]  axi4Port_w_bits_strb,
  input          axi4Port_b_valid,
  input  [1:0]   axi4Port_b_bits_id,
                 axi4Port_b_bits_resp,
  input          axi4Port_ar_ready,
  output         axi4Port_ar_valid,
  output [31:0]  axi4Port_ar_bits_addr,
  output         axi4Port_r_ready,
  input          axi4Port_r_valid,
  input  [1:0]   axi4Port_r_bits_id,
  input  [127:0] axi4Port_r_bits_data,
  input  [1:0]   axi4Port_r_bits_resp,
  input          axi4Port_r_bits_last,
                 simpleAccessPorts_aw_ready,
  output         simpleAccessPorts_aw_valid,
  output [1:0]   simpleAccessPorts_aw_bits_id,
  output [31:0]  simpleAccessPorts_aw_bits_addr,
  output [2:0]   simpleAccessPorts_aw_bits_size,
  input          simpleAccessPorts_w_ready,
  output         simpleAccessPorts_w_valid,
  output [31:0]  simpleAccessPorts_w_bits_data,
  output [3:0]   simpleAccessPorts_w_bits_strb,
  input          simpleAccessPorts_b_valid,
  input  [1:0]   simpleAccessPorts_b_bits_id,
                 simpleAccessPorts_b_bits_resp,
  input          simpleAccessPorts_ar_ready,
  output         simpleAccessPorts_ar_valid,
  output [31:0]  simpleAccessPorts_ar_bits_addr,
  output         simpleAccessPorts_r_ready,
  input          simpleAccessPorts_r_valid,
  input  [1:0]   simpleAccessPorts_r_bits_id,
  input  [31:0]  simpleAccessPorts_r_bits_data,
  input  [1:0]   simpleAccessPorts_r_bits_resp,
  input          simpleAccessPorts_r_bits_last,
                 vrfReadDataPorts_0_ready,
  output         vrfReadDataPorts_0_valid,
  output [4:0]   vrfReadDataPorts_0_bits_vs,
  output [8:0]   vrfReadDataPorts_0_bits_offset,
  output [2:0]   vrfReadDataPorts_0_bits_instructionIndex,
  input          vrfReadDataPorts_1_ready,
  output         vrfReadDataPorts_1_valid,
  output [4:0]   vrfReadDataPorts_1_bits_vs,
  output [8:0]   vrfReadDataPorts_1_bits_offset,
  output [2:0]   vrfReadDataPorts_1_bits_instructionIndex,
  input          vrfReadDataPorts_2_ready,
  output         vrfReadDataPorts_2_valid,
  output [4:0]   vrfReadDataPorts_2_bits_vs,
  output [8:0]   vrfReadDataPorts_2_bits_offset,
  output [2:0]   vrfReadDataPorts_2_bits_instructionIndex,
  input          vrfReadDataPorts_3_ready,
  output         vrfReadDataPorts_3_valid,
  output [4:0]   vrfReadDataPorts_3_bits_vs,
  output [8:0]   vrfReadDataPorts_3_bits_offset,
  output [2:0]   vrfReadDataPorts_3_bits_instructionIndex,
  input          vrfReadResults_0_valid,
  input  [31:0]  vrfReadResults_0_bits,
  input          vrfReadResults_1_valid,
  input  [31:0]  vrfReadResults_1_bits,
  input          vrfReadResults_2_valid,
  input  [31:0]  vrfReadResults_2_bits,
  input          vrfReadResults_3_valid,
  input  [31:0]  vrfReadResults_3_bits,
  input          vrfWritePort_0_ready,
  output         vrfWritePort_0_valid,
  output [4:0]   vrfWritePort_0_bits_vd,
  output [8:0]   vrfWritePort_0_bits_offset,
  output [3:0]   vrfWritePort_0_bits_mask,
  output [31:0]  vrfWritePort_0_bits_data,
  output         vrfWritePort_0_bits_last,
  output [2:0]   vrfWritePort_0_bits_instructionIndex,
  input          vrfWritePort_1_ready,
  output         vrfWritePort_1_valid,
  output [4:0]   vrfWritePort_1_bits_vd,
  output [8:0]   vrfWritePort_1_bits_offset,
  output [3:0]   vrfWritePort_1_bits_mask,
  output [31:0]  vrfWritePort_1_bits_data,
  output         vrfWritePort_1_bits_last,
  output [2:0]   vrfWritePort_1_bits_instructionIndex,
  input          vrfWritePort_2_ready,
  output         vrfWritePort_2_valid,
  output [4:0]   vrfWritePort_2_bits_vd,
  output [8:0]   vrfWritePort_2_bits_offset,
  output [3:0]   vrfWritePort_2_bits_mask,
  output [31:0]  vrfWritePort_2_bits_data,
  output         vrfWritePort_2_bits_last,
  output [2:0]   vrfWritePort_2_bits_instructionIndex,
  input          vrfWritePort_3_ready,
  output         vrfWritePort_3_valid,
  output [4:0]   vrfWritePort_3_bits_vd,
  output [8:0]   vrfWritePort_3_bits_offset,
  output [3:0]   vrfWritePort_3_bits_mask,
  output [31:0]  vrfWritePort_3_bits_data,
  output         vrfWritePort_3_bits_last,
  output [2:0]   vrfWritePort_3_bits_instructionIndex,
  input          writeRelease_0,
                 writeRelease_1,
                 writeRelease_2,
                 writeRelease_3,
  output [7:0]   dataInWriteQueue_0,
                 dataInWriteQueue_1,
                 dataInWriteQueue_2,
                 dataInWriteQueue_3,
  input  [16:0]  csrInterface_vl,
                 csrInterface_vStart,
  input  [2:0]   csrInterface_vlmul,
  input  [1:0]   csrInterface_vSew,
                 csrInterface_vxrm,
  input          csrInterface_vta,
                 csrInterface_vma,
                 offsetReadResult_0_valid,
  input  [31:0]  offsetReadResult_0_bits,
  input          offsetReadResult_1_valid,
  input  [31:0]  offsetReadResult_1_bits,
  input          offsetReadResult_2_valid,
  input  [31:0]  offsetReadResult_2_bits,
  input          offsetReadResult_3_valid,
  input  [31:0]  offsetReadResult_3_bits,
  output [7:0]   lastReport,
  output [3:0]   tokenIO_offsetGroupRelease
);

  wire                _simpleDataQueue_fifo_empty;
  wire                _simpleDataQueue_fifo_full;
  wire                _simpleDataQueue_fifo_error;
  wire [77:0]         _simpleDataQueue_fifo_data_out;
  wire                _simpleSourceQueue_fifo_empty;
  wire                _simpleSourceQueue_fifo_full;
  wire                _simpleSourceQueue_fifo_error;
  wire                _dataQueue_fifo_empty;
  wire                _dataQueue_fifo_full;
  wire                _dataQueue_fifo_error;
  wire [188:0]        _dataQueue_fifo_data_out;
  wire                _sourceQueue_fifo_empty;
  wire                _sourceQueue_fifo_full;
  wire                _sourceQueue_fifo_error;
  wire                _writeIndexQueue_fifo_3_empty;
  wire                _writeIndexQueue_fifo_3_full;
  wire                _writeIndexQueue_fifo_3_error;
  wire                _writeIndexQueue_fifo_2_empty;
  wire                _writeIndexQueue_fifo_2_full;
  wire                _writeIndexQueue_fifo_2_error;
  wire                _writeIndexQueue_fifo_1_empty;
  wire                _writeIndexQueue_fifo_1_full;
  wire                _writeIndexQueue_fifo_1_error;
  wire                _writeIndexQueue_fifo_empty;
  wire                _writeIndexQueue_fifo_full;
  wire                _writeIndexQueue_fifo_error;
  wire                _otherUnitDataQueueVec_fifo_3_empty;
  wire                _otherUnitDataQueueVec_fifo_3_full;
  wire                _otherUnitDataQueueVec_fifo_3_error;
  wire [31:0]         _otherUnitDataQueueVec_fifo_3_data_out;
  wire                _otherUnitDataQueueVec_fifo_2_empty;
  wire                _otherUnitDataQueueVec_fifo_2_full;
  wire                _otherUnitDataQueueVec_fifo_2_error;
  wire [31:0]         _otherUnitDataQueueVec_fifo_2_data_out;
  wire                _otherUnitDataQueueVec_fifo_1_empty;
  wire                _otherUnitDataQueueVec_fifo_1_full;
  wire                _otherUnitDataQueueVec_fifo_1_error;
  wire [31:0]         _otherUnitDataQueueVec_fifo_1_data_out;
  wire                _otherUnitDataQueueVec_fifo_empty;
  wire                _otherUnitDataQueueVec_fifo_full;
  wire                _otherUnitDataQueueVec_fifo_error;
  wire [31:0]         _otherUnitDataQueueVec_fifo_data_out;
  wire                _otherUnitTargetQueue_fifo_empty;
  wire                _otherUnitTargetQueue_fifo_full;
  wire                _otherUnitTargetQueue_fifo_error;
  wire                _writeQueueVec_fifo_3_empty;
  wire                _writeQueueVec_fifo_3_full;
  wire                _writeQueueVec_fifo_3_error;
  wire [57:0]         _writeQueueVec_fifo_3_data_out;
  wire                _writeQueueVec_fifo_2_empty;
  wire                _writeQueueVec_fifo_2_full;
  wire                _writeQueueVec_fifo_2_error;
  wire [57:0]         _writeQueueVec_fifo_2_data_out;
  wire                _writeQueueVec_fifo_1_empty;
  wire                _writeQueueVec_fifo_1_full;
  wire                _writeQueueVec_fifo_1_error;
  wire [57:0]         _writeQueueVec_fifo_1_data_out;
  wire                _writeQueueVec_fifo_empty;
  wire                _writeQueueVec_fifo_full;
  wire                _writeQueueVec_fifo_error;
  wire [57:0]         _writeQueueVec_fifo_data_out;
  wire                _otherUnit_vrfReadDataPorts_valid;
  wire [4:0]          _otherUnit_vrfReadDataPorts_bits_vs;
  wire [8:0]          _otherUnit_vrfReadDataPorts_bits_offset;
  wire [2:0]          _otherUnit_vrfReadDataPorts_bits_instructionIndex;
  wire                _otherUnit_maskSelect_valid;
  wire [11:0]         _otherUnit_maskSelect_bits;
  wire                _otherUnit_memReadRequest_valid;
  wire                _otherUnit_memWriteRequest_valid;
  wire [7:0]          _otherUnit_memWriteRequest_bits_source;
  wire [31:0]         _otherUnit_memWriteRequest_bits_address;
  wire [1:0]          _otherUnit_memWriteRequest_bits_size;
  wire                _otherUnit_vrfWritePort_valid;
  wire [4:0]          _otherUnit_vrfWritePort_bits_vd;
  wire [8:0]          _otherUnit_vrfWritePort_bits_offset;
  wire [3:0]          _otherUnit_vrfWritePort_bits_mask;
  wire [31:0]         _otherUnit_vrfWritePort_bits_data;
  wire                _otherUnit_vrfWritePort_bits_last;
  wire [2:0]          _otherUnit_vrfWritePort_bits_instructionIndex;
  wire                _otherUnit_status_idle;
  wire                _otherUnit_status_last;
  wire [2:0]          _otherUnit_status_instructionIndex;
  wire [3:0]          _otherUnit_status_targetLane;
  wire                _otherUnit_status_isStore;
  wire                _otherUnit_offsetRelease_0;
  wire                _otherUnit_offsetRelease_1;
  wire                _otherUnit_offsetRelease_2;
  wire                _otherUnit_offsetRelease_3;
  wire                _storeUnit_maskSelect_valid;
  wire [11:0]         _storeUnit_maskSelect_bits;
  wire                _storeUnit_memRequest_valid;
  wire [12:0]         _storeUnit_memRequest_bits_index;
  wire [31:0]         _storeUnit_memRequest_bits_address;
  wire                _storeUnit_status_idle;
  wire                _storeUnit_status_last;
  wire [2:0]          _storeUnit_status_instructionIndex;
  wire [31:0]         _storeUnit_status_startAddress;
  wire [31:0]         _storeUnit_status_endAddress;
  wire                _storeUnit_vrfReadDataPorts_0_valid;
  wire [4:0]          _storeUnit_vrfReadDataPorts_0_bits_vs;
  wire [8:0]          _storeUnit_vrfReadDataPorts_0_bits_offset;
  wire [2:0]          _storeUnit_vrfReadDataPorts_0_bits_instructionIndex;
  wire                _storeUnit_vrfReadDataPorts_1_valid;
  wire [4:0]          _storeUnit_vrfReadDataPorts_1_bits_vs;
  wire [8:0]          _storeUnit_vrfReadDataPorts_1_bits_offset;
  wire [2:0]          _storeUnit_vrfReadDataPorts_1_bits_instructionIndex;
  wire                _storeUnit_vrfReadDataPorts_2_valid;
  wire [4:0]          _storeUnit_vrfReadDataPorts_2_bits_vs;
  wire [8:0]          _storeUnit_vrfReadDataPorts_2_bits_offset;
  wire [2:0]          _storeUnit_vrfReadDataPorts_2_bits_instructionIndex;
  wire                _storeUnit_vrfReadDataPorts_3_valid;
  wire [4:0]          _storeUnit_vrfReadDataPorts_3_bits_vs;
  wire [8:0]          _storeUnit_vrfReadDataPorts_3_bits_offset;
  wire [2:0]          _storeUnit_vrfReadDataPorts_3_bits_instructionIndex;
  wire                _loadUnit_maskSelect_valid;
  wire [11:0]         _loadUnit_maskSelect_bits;
  wire                _loadUnit_memRequest_valid;
  wire                _loadUnit_status_idle;
  wire                _loadUnit_status_last;
  wire [2:0]          _loadUnit_status_instructionIndex;
  wire [31:0]         _loadUnit_status_startAddress;
  wire [31:0]         _loadUnit_status_endAddress;
  wire                _loadUnit_vrfWritePort_0_valid;
  wire [4:0]          _loadUnit_vrfWritePort_0_bits_vd;
  wire [8:0]          _loadUnit_vrfWritePort_0_bits_offset;
  wire [3:0]          _loadUnit_vrfWritePort_0_bits_mask;
  wire [31:0]         _loadUnit_vrfWritePort_0_bits_data;
  wire [2:0]          _loadUnit_vrfWritePort_0_bits_instructionIndex;
  wire                _loadUnit_vrfWritePort_1_valid;
  wire [4:0]          _loadUnit_vrfWritePort_1_bits_vd;
  wire [8:0]          _loadUnit_vrfWritePort_1_bits_offset;
  wire [3:0]          _loadUnit_vrfWritePort_1_bits_mask;
  wire [31:0]         _loadUnit_vrfWritePort_1_bits_data;
  wire [2:0]          _loadUnit_vrfWritePort_1_bits_instructionIndex;
  wire                _loadUnit_vrfWritePort_2_valid;
  wire [4:0]          _loadUnit_vrfWritePort_2_bits_vd;
  wire [8:0]          _loadUnit_vrfWritePort_2_bits_offset;
  wire [3:0]          _loadUnit_vrfWritePort_2_bits_mask;
  wire [31:0]         _loadUnit_vrfWritePort_2_bits_data;
  wire [2:0]          _loadUnit_vrfWritePort_2_bits_instructionIndex;
  wire                _loadUnit_vrfWritePort_3_valid;
  wire [4:0]          _loadUnit_vrfWritePort_3_bits_vd;
  wire [8:0]          _loadUnit_vrfWritePort_3_bits_offset;
  wire [3:0]          _loadUnit_vrfWritePort_3_bits_mask;
  wire [31:0]         _loadUnit_vrfWritePort_3_bits_data;
  wire [2:0]          _loadUnit_vrfWritePort_3_bits_instructionIndex;
  wire                simpleDataQueue_almostFull;
  wire                simpleDataQueue_almostEmpty;
  wire                simpleSourceQueue_almostFull;
  wire                simpleSourceQueue_almostEmpty;
  wire                dataQueue_almostFull;
  wire                dataQueue_almostEmpty;
  wire                sourceQueue_almostFull;
  wire                sourceQueue_almostEmpty;
  wire                writeIndexQueue_3_almostFull;
  wire                writeIndexQueue_3_almostEmpty;
  wire                writeIndexQueue_2_almostFull;
  wire                writeIndexQueue_2_almostEmpty;
  wire                writeIndexQueue_1_almostFull;
  wire                writeIndexQueue_1_almostEmpty;
  wire                writeIndexQueue_almostFull;
  wire                writeIndexQueue_almostEmpty;
  wire                otherUnitDataQueueVec_3_almostFull;
  wire                otherUnitDataQueueVec_3_almostEmpty;
  wire                otherUnitDataQueueVec_2_almostFull;
  wire                otherUnitDataQueueVec_2_almostEmpty;
  wire                otherUnitDataQueueVec_1_almostFull;
  wire                otherUnitDataQueueVec_1_almostEmpty;
  wire                otherUnitDataQueueVec_0_almostFull;
  wire                otherUnitDataQueueVec_0_almostEmpty;
  wire                otherUnitTargetQueue_almostFull;
  wire                otherUnitTargetQueue_almostEmpty;
  wire                writeQueueVec_3_almostFull;
  wire                writeQueueVec_3_almostEmpty;
  wire                writeQueueVec_2_almostFull;
  wire                writeQueueVec_2_almostEmpty;
  wire                writeQueueVec_1_almostFull;
  wire                writeQueueVec_1_almostEmpty;
  wire                writeQueueVec_0_almostFull;
  wire                writeQueueVec_0_almostEmpty;
  wire [6:0]          simpleSourceQueue_enq_bits;
  wire [31:0]         simpleAccessPorts_ar_bits_addr_0;
  wire [12:0]         sourceQueue_enq_bits;
  wire [31:0]         axi4Port_ar_bits_addr_0;
  wire                request_valid_0 = request_valid;
  wire [2:0]          request_bits_instructionInformation_nf_0 = request_bits_instructionInformation_nf;
  wire                request_bits_instructionInformation_mew_0 = request_bits_instructionInformation_mew;
  wire [1:0]          request_bits_instructionInformation_mop_0 = request_bits_instructionInformation_mop;
  wire [4:0]          request_bits_instructionInformation_lumop_0 = request_bits_instructionInformation_lumop;
  wire [1:0]          request_bits_instructionInformation_eew_0 = request_bits_instructionInformation_eew;
  wire [4:0]          request_bits_instructionInformation_vs3_0 = request_bits_instructionInformation_vs3;
  wire                request_bits_instructionInformation_isStore_0 = request_bits_instructionInformation_isStore;
  wire                request_bits_instructionInformation_maskedLoadStore_0 = request_bits_instructionInformation_maskedLoadStore;
  wire [31:0]         request_bits_rs1Data_0 = request_bits_rs1Data;
  wire [31:0]         request_bits_rs2Data_0 = request_bits_rs2Data;
  wire [2:0]          request_bits_instructionIndex_0 = request_bits_instructionIndex;
  wire                axi4Port_aw_ready_0 = axi4Port_aw_ready;
  wire                axi4Port_w_ready_0 = axi4Port_w_ready;
  wire                axi4Port_b_valid_0 = axi4Port_b_valid;
  wire [1:0]          axi4Port_b_bits_id_0 = axi4Port_b_bits_id;
  wire [1:0]          axi4Port_b_bits_resp_0 = axi4Port_b_bits_resp;
  wire                axi4Port_ar_ready_0 = axi4Port_ar_ready;
  wire                axi4Port_r_valid_0 = axi4Port_r_valid;
  wire [1:0]          axi4Port_r_bits_id_0 = axi4Port_r_bits_id;
  wire [127:0]        axi4Port_r_bits_data_0 = axi4Port_r_bits_data;
  wire [1:0]          axi4Port_r_bits_resp_0 = axi4Port_r_bits_resp;
  wire                axi4Port_r_bits_last_0 = axi4Port_r_bits_last;
  wire                simpleAccessPorts_aw_ready_0 = simpleAccessPorts_aw_ready;
  wire                simpleAccessPorts_w_ready_0 = simpleAccessPorts_w_ready;
  wire                simpleAccessPorts_b_valid_0 = simpleAccessPorts_b_valid;
  wire [1:0]          simpleAccessPorts_b_bits_id_0 = simpleAccessPorts_b_bits_id;
  wire [1:0]          simpleAccessPorts_b_bits_resp_0 = simpleAccessPorts_b_bits_resp;
  wire                simpleAccessPorts_ar_ready_0 = simpleAccessPorts_ar_ready;
  wire                simpleAccessPorts_r_valid_0 = simpleAccessPorts_r_valid;
  wire [1:0]          simpleAccessPorts_r_bits_id_0 = simpleAccessPorts_r_bits_id;
  wire [31:0]         simpleAccessPorts_r_bits_data_0 = simpleAccessPorts_r_bits_data;
  wire [1:0]          simpleAccessPorts_r_bits_resp_0 = simpleAccessPorts_r_bits_resp;
  wire                simpleAccessPorts_r_bits_last_0 = simpleAccessPorts_r_bits_last;
  wire                vrfReadDataPorts_0_ready_0 = vrfReadDataPorts_0_ready;
  wire                vrfReadDataPorts_1_ready_0 = vrfReadDataPorts_1_ready;
  wire                vrfReadDataPorts_2_ready_0 = vrfReadDataPorts_2_ready;
  wire                vrfReadDataPorts_3_ready_0 = vrfReadDataPorts_3_ready;
  wire                vrfWritePort_0_ready_0 = vrfWritePort_0_ready;
  wire                vrfWritePort_1_ready_0 = vrfWritePort_1_ready;
  wire                vrfWritePort_2_ready_0 = vrfWritePort_2_ready;
  wire                vrfWritePort_3_ready_0 = vrfWritePort_3_ready;
  wire [31:0]         otherUnitDataQueueVec_0_enq_bits = vrfReadResults_0_bits;
  wire [31:0]         otherUnitDataQueueVec_1_enq_bits = vrfReadResults_1_bits;
  wire [31:0]         otherUnitDataQueueVec_2_enq_bits = vrfReadResults_2_bits;
  wire [31:0]         otherUnitDataQueueVec_3_enq_bits = vrfReadResults_3_bits;
  wire                writeIndexQueue_deq_ready = writeRelease_0;
  wire                writeIndexQueue_1_deq_ready = writeRelease_1;
  wire                writeIndexQueue_2_deq_ready = writeRelease_2;
  wire                writeIndexQueue_3_deq_ready = writeRelease_3;
  wire [1:0]          vrfReadDataPorts_0_bits_readSource = 2'h2;
  wire [1:0]          vrfReadDataPorts_1_bits_readSource = 2'h2;
  wire [1:0]          vrfReadDataPorts_2_bits_readSource = 2'h2;
  wire [1:0]          vrfReadDataPorts_3_bits_readSource = 2'h2;
  wire [1:0]          axi4Port_ar_bits_id = 2'h0;
  wire [1:0]          simpleAccessPorts_ar_bits_id = 2'h0;
  wire [1:0]          axi4Port_aw_bits_burst = 2'h1;
  wire [1:0]          axi4Port_ar_bits_burst = 2'h1;
  wire [1:0]          simpleAccessPorts_aw_bits_burst = 2'h1;
  wire [1:0]          simpleAccessPorts_ar_bits_burst = 2'h1;
  wire [3:0]          writeQueueVec_0_enq_bits_targetLane = 4'h1;
  wire [3:0]          writeQueueVec_1_enq_bits_targetLane = 4'h2;
  wire [3:0]          writeQueueVec_2_enq_bits_targetLane = 4'h4;
  wire [3:0]          writeQueueVec_3_enq_bits_targetLane = 4'h8;
  wire [7:0]          axi4Port_aw_bits_len = 8'h0;
  wire [7:0]          axi4Port_ar_bits_len = 8'h0;
  wire [7:0]          simpleAccessPorts_aw_bits_len = 8'h0;
  wire [7:0]          simpleAccessPorts_ar_bits_len = 8'h0;
  wire [2:0]          axi4Port_aw_bits_size = 3'h4;
  wire [2:0]          axi4Port_ar_bits_size = 3'h4;
  wire                axi4Port_aw_bits_lock = 1'h0;
  wire                axi4Port_ar_bits_lock = 1'h0;
  wire                simpleAccessPorts_aw_bits_lock = 1'h0;
  wire                simpleAccessPorts_ar_bits_lock = 1'h0;
  wire [3:0]          axi4Port_aw_bits_cache = 4'h0;
  wire [3:0]          axi4Port_aw_bits_qos = 4'h0;
  wire [3:0]          axi4Port_aw_bits_region = 4'h0;
  wire [3:0]          axi4Port_ar_bits_cache = 4'h0;
  wire [3:0]          axi4Port_ar_bits_qos = 4'h0;
  wire [3:0]          axi4Port_ar_bits_region = 4'h0;
  wire [3:0]          simpleAccessPorts_aw_bits_cache = 4'h0;
  wire [3:0]          simpleAccessPorts_aw_bits_qos = 4'h0;
  wire [3:0]          simpleAccessPorts_aw_bits_region = 4'h0;
  wire [3:0]          simpleAccessPorts_ar_bits_cache = 4'h0;
  wire [3:0]          simpleAccessPorts_ar_bits_qos = 4'h0;
  wire [3:0]          simpleAccessPorts_ar_bits_region = 4'h0;
  wire [2:0]          axi4Port_aw_bits_prot = 3'h0;
  wire [2:0]          axi4Port_ar_bits_prot = 3'h0;
  wire [2:0]          simpleAccessPorts_aw_bits_prot = 3'h0;
  wire [2:0]          simpleAccessPorts_ar_bits_prot = 3'h0;
  wire                axi4Port_w_bits_last = 1'h1;
  wire                axi4Port_b_ready = 1'h1;
  wire                simpleAccessPorts_w_bits_last = 1'h1;
  wire                simpleAccessPorts_b_ready = 1'h1;
  wire [2:0]          simpleAccessPorts_ar_bits_size = 3'h2;
  wire                dataQueue_deq_ready = axi4Port_w_ready_0;
  wire                dataQueue_deq_valid;
  wire [127:0]        dataQueue_deq_bits_data;
  wire [15:0]         dataQueue_deq_bits_mask;
  wire                simpleDataQueue_deq_ready = simpleAccessPorts_w_ready_0;
  wire                simpleDataQueue_deq_valid;
  wire [31:0]         simpleDataQueue_deq_bits_data;
  wire [3:0]          simpleDataQueue_deq_bits_mask;
  wire                writeQueueVec_0_deq_ready = vrfWritePort_0_ready_0;
  wire                writeQueueVec_0_deq_valid;
  wire [4:0]          writeQueueVec_0_deq_bits_data_vd;
  wire [8:0]          writeQueueVec_0_deq_bits_data_offset;
  wire [3:0]          writeQueueVec_0_deq_bits_data_mask;
  wire [31:0]         writeQueueVec_0_deq_bits_data_data;
  wire                writeQueueVec_0_deq_bits_data_last;
  wire [2:0]          writeQueueVec_0_deq_bits_data_instructionIndex;
  wire                writeQueueVec_1_deq_ready = vrfWritePort_1_ready_0;
  wire                writeQueueVec_1_deq_valid;
  wire [4:0]          writeQueueVec_1_deq_bits_data_vd;
  wire [8:0]          writeQueueVec_1_deq_bits_data_offset;
  wire [3:0]          writeQueueVec_1_deq_bits_data_mask;
  wire [31:0]         writeQueueVec_1_deq_bits_data_data;
  wire                writeQueueVec_1_deq_bits_data_last;
  wire [2:0]          writeQueueVec_1_deq_bits_data_instructionIndex;
  wire                writeQueueVec_2_deq_ready = vrfWritePort_2_ready_0;
  wire                writeQueueVec_2_deq_valid;
  wire [4:0]          writeQueueVec_2_deq_bits_data_vd;
  wire [8:0]          writeQueueVec_2_deq_bits_data_offset;
  wire [3:0]          writeQueueVec_2_deq_bits_data_mask;
  wire [31:0]         writeQueueVec_2_deq_bits_data_data;
  wire                writeQueueVec_2_deq_bits_data_last;
  wire [2:0]          writeQueueVec_2_deq_bits_data_instructionIndex;
  wire                writeQueueVec_3_deq_ready = vrfWritePort_3_ready_0;
  wire                writeQueueVec_3_deq_valid;
  wire [4:0]          writeQueueVec_3_deq_bits_data_vd;
  wire [8:0]          writeQueueVec_3_deq_bits_data_offset;
  wire [3:0]          writeQueueVec_3_deq_bits_data_mask;
  wire [31:0]         writeQueueVec_3_deq_bits_data_data;
  wire                writeQueueVec_3_deq_bits_data_last;
  wire [2:0]          writeQueueVec_3_deq_bits_data_instructionIndex;
  reg  [31:0]         v0_0;
  reg  [31:0]         v0_1;
  reg  [31:0]         v0_2;
  reg  [31:0]         v0_3;
  reg  [31:0]         v0_4;
  reg  [31:0]         v0_5;
  reg  [31:0]         v0_6;
  reg  [31:0]         v0_7;
  reg  [31:0]         v0_8;
  reg  [31:0]         v0_9;
  reg  [31:0]         v0_10;
  reg  [31:0]         v0_11;
  reg  [31:0]         v0_12;
  reg  [31:0]         v0_13;
  reg  [31:0]         v0_14;
  reg  [31:0]         v0_15;
  reg  [31:0]         v0_16;
  reg  [31:0]         v0_17;
  reg  [31:0]         v0_18;
  reg  [31:0]         v0_19;
  reg  [31:0]         v0_20;
  reg  [31:0]         v0_21;
  reg  [31:0]         v0_22;
  reg  [31:0]         v0_23;
  reg  [31:0]         v0_24;
  reg  [31:0]         v0_25;
  reg  [31:0]         v0_26;
  reg  [31:0]         v0_27;
  reg  [31:0]         v0_28;
  reg  [31:0]         v0_29;
  reg  [31:0]         v0_30;
  reg  [31:0]         v0_31;
  reg  [31:0]         v0_32;
  reg  [31:0]         v0_33;
  reg  [31:0]         v0_34;
  reg  [31:0]         v0_35;
  reg  [31:0]         v0_36;
  reg  [31:0]         v0_37;
  reg  [31:0]         v0_38;
  reg  [31:0]         v0_39;
  reg  [31:0]         v0_40;
  reg  [31:0]         v0_41;
  reg  [31:0]         v0_42;
  reg  [31:0]         v0_43;
  reg  [31:0]         v0_44;
  reg  [31:0]         v0_45;
  reg  [31:0]         v0_46;
  reg  [31:0]         v0_47;
  reg  [31:0]         v0_48;
  reg  [31:0]         v0_49;
  reg  [31:0]         v0_50;
  reg  [31:0]         v0_51;
  reg  [31:0]         v0_52;
  reg  [31:0]         v0_53;
  reg  [31:0]         v0_54;
  reg  [31:0]         v0_55;
  reg  [31:0]         v0_56;
  reg  [31:0]         v0_57;
  reg  [31:0]         v0_58;
  reg  [31:0]         v0_59;
  reg  [31:0]         v0_60;
  reg  [31:0]         v0_61;
  reg  [31:0]         v0_62;
  reg  [31:0]         v0_63;
  reg  [31:0]         v0_64;
  reg  [31:0]         v0_65;
  reg  [31:0]         v0_66;
  reg  [31:0]         v0_67;
  reg  [31:0]         v0_68;
  reg  [31:0]         v0_69;
  reg  [31:0]         v0_70;
  reg  [31:0]         v0_71;
  reg  [31:0]         v0_72;
  reg  [31:0]         v0_73;
  reg  [31:0]         v0_74;
  reg  [31:0]         v0_75;
  reg  [31:0]         v0_76;
  reg  [31:0]         v0_77;
  reg  [31:0]         v0_78;
  reg  [31:0]         v0_79;
  reg  [31:0]         v0_80;
  reg  [31:0]         v0_81;
  reg  [31:0]         v0_82;
  reg  [31:0]         v0_83;
  reg  [31:0]         v0_84;
  reg  [31:0]         v0_85;
  reg  [31:0]         v0_86;
  reg  [31:0]         v0_87;
  reg  [31:0]         v0_88;
  reg  [31:0]         v0_89;
  reg  [31:0]         v0_90;
  reg  [31:0]         v0_91;
  reg  [31:0]         v0_92;
  reg  [31:0]         v0_93;
  reg  [31:0]         v0_94;
  reg  [31:0]         v0_95;
  reg  [31:0]         v0_96;
  reg  [31:0]         v0_97;
  reg  [31:0]         v0_98;
  reg  [31:0]         v0_99;
  reg  [31:0]         v0_100;
  reg  [31:0]         v0_101;
  reg  [31:0]         v0_102;
  reg  [31:0]         v0_103;
  reg  [31:0]         v0_104;
  reg  [31:0]         v0_105;
  reg  [31:0]         v0_106;
  reg  [31:0]         v0_107;
  reg  [31:0]         v0_108;
  reg  [31:0]         v0_109;
  reg  [31:0]         v0_110;
  reg  [31:0]         v0_111;
  reg  [31:0]         v0_112;
  reg  [31:0]         v0_113;
  reg  [31:0]         v0_114;
  reg  [31:0]         v0_115;
  reg  [31:0]         v0_116;
  reg  [31:0]         v0_117;
  reg  [31:0]         v0_118;
  reg  [31:0]         v0_119;
  reg  [31:0]         v0_120;
  reg  [31:0]         v0_121;
  reg  [31:0]         v0_122;
  reg  [31:0]         v0_123;
  reg  [31:0]         v0_124;
  reg  [31:0]         v0_125;
  reg  [31:0]         v0_126;
  reg  [31:0]         v0_127;
  reg  [31:0]         v0_128;
  reg  [31:0]         v0_129;
  reg  [31:0]         v0_130;
  reg  [31:0]         v0_131;
  reg  [31:0]         v0_132;
  reg  [31:0]         v0_133;
  reg  [31:0]         v0_134;
  reg  [31:0]         v0_135;
  reg  [31:0]         v0_136;
  reg  [31:0]         v0_137;
  reg  [31:0]         v0_138;
  reg  [31:0]         v0_139;
  reg  [31:0]         v0_140;
  reg  [31:0]         v0_141;
  reg  [31:0]         v0_142;
  reg  [31:0]         v0_143;
  reg  [31:0]         v0_144;
  reg  [31:0]         v0_145;
  reg  [31:0]         v0_146;
  reg  [31:0]         v0_147;
  reg  [31:0]         v0_148;
  reg  [31:0]         v0_149;
  reg  [31:0]         v0_150;
  reg  [31:0]         v0_151;
  reg  [31:0]         v0_152;
  reg  [31:0]         v0_153;
  reg  [31:0]         v0_154;
  reg  [31:0]         v0_155;
  reg  [31:0]         v0_156;
  reg  [31:0]         v0_157;
  reg  [31:0]         v0_158;
  reg  [31:0]         v0_159;
  reg  [31:0]         v0_160;
  reg  [31:0]         v0_161;
  reg  [31:0]         v0_162;
  reg  [31:0]         v0_163;
  reg  [31:0]         v0_164;
  reg  [31:0]         v0_165;
  reg  [31:0]         v0_166;
  reg  [31:0]         v0_167;
  reg  [31:0]         v0_168;
  reg  [31:0]         v0_169;
  reg  [31:0]         v0_170;
  reg  [31:0]         v0_171;
  reg  [31:0]         v0_172;
  reg  [31:0]         v0_173;
  reg  [31:0]         v0_174;
  reg  [31:0]         v0_175;
  reg  [31:0]         v0_176;
  reg  [31:0]         v0_177;
  reg  [31:0]         v0_178;
  reg  [31:0]         v0_179;
  reg  [31:0]         v0_180;
  reg  [31:0]         v0_181;
  reg  [31:0]         v0_182;
  reg  [31:0]         v0_183;
  reg  [31:0]         v0_184;
  reg  [31:0]         v0_185;
  reg  [31:0]         v0_186;
  reg  [31:0]         v0_187;
  reg  [31:0]         v0_188;
  reg  [31:0]         v0_189;
  reg  [31:0]         v0_190;
  reg  [31:0]         v0_191;
  reg  [31:0]         v0_192;
  reg  [31:0]         v0_193;
  reg  [31:0]         v0_194;
  reg  [31:0]         v0_195;
  reg  [31:0]         v0_196;
  reg  [31:0]         v0_197;
  reg  [31:0]         v0_198;
  reg  [31:0]         v0_199;
  reg  [31:0]         v0_200;
  reg  [31:0]         v0_201;
  reg  [31:0]         v0_202;
  reg  [31:0]         v0_203;
  reg  [31:0]         v0_204;
  reg  [31:0]         v0_205;
  reg  [31:0]         v0_206;
  reg  [31:0]         v0_207;
  reg  [31:0]         v0_208;
  reg  [31:0]         v0_209;
  reg  [31:0]         v0_210;
  reg  [31:0]         v0_211;
  reg  [31:0]         v0_212;
  reg  [31:0]         v0_213;
  reg  [31:0]         v0_214;
  reg  [31:0]         v0_215;
  reg  [31:0]         v0_216;
  reg  [31:0]         v0_217;
  reg  [31:0]         v0_218;
  reg  [31:0]         v0_219;
  reg  [31:0]         v0_220;
  reg  [31:0]         v0_221;
  reg  [31:0]         v0_222;
  reg  [31:0]         v0_223;
  reg  [31:0]         v0_224;
  reg  [31:0]         v0_225;
  reg  [31:0]         v0_226;
  reg  [31:0]         v0_227;
  reg  [31:0]         v0_228;
  reg  [31:0]         v0_229;
  reg  [31:0]         v0_230;
  reg  [31:0]         v0_231;
  reg  [31:0]         v0_232;
  reg  [31:0]         v0_233;
  reg  [31:0]         v0_234;
  reg  [31:0]         v0_235;
  reg  [31:0]         v0_236;
  reg  [31:0]         v0_237;
  reg  [31:0]         v0_238;
  reg  [31:0]         v0_239;
  reg  [31:0]         v0_240;
  reg  [31:0]         v0_241;
  reg  [31:0]         v0_242;
  reg  [31:0]         v0_243;
  reg  [31:0]         v0_244;
  reg  [31:0]         v0_245;
  reg  [31:0]         v0_246;
  reg  [31:0]         v0_247;
  reg  [31:0]         v0_248;
  reg  [31:0]         v0_249;
  reg  [31:0]         v0_250;
  reg  [31:0]         v0_251;
  reg  [31:0]         v0_252;
  reg  [31:0]         v0_253;
  reg  [31:0]         v0_254;
  reg  [31:0]         v0_255;
  reg  [31:0]         v0_256;
  reg  [31:0]         v0_257;
  reg  [31:0]         v0_258;
  reg  [31:0]         v0_259;
  reg  [31:0]         v0_260;
  reg  [31:0]         v0_261;
  reg  [31:0]         v0_262;
  reg  [31:0]         v0_263;
  reg  [31:0]         v0_264;
  reg  [31:0]         v0_265;
  reg  [31:0]         v0_266;
  reg  [31:0]         v0_267;
  reg  [31:0]         v0_268;
  reg  [31:0]         v0_269;
  reg  [31:0]         v0_270;
  reg  [31:0]         v0_271;
  reg  [31:0]         v0_272;
  reg  [31:0]         v0_273;
  reg  [31:0]         v0_274;
  reg  [31:0]         v0_275;
  reg  [31:0]         v0_276;
  reg  [31:0]         v0_277;
  reg  [31:0]         v0_278;
  reg  [31:0]         v0_279;
  reg  [31:0]         v0_280;
  reg  [31:0]         v0_281;
  reg  [31:0]         v0_282;
  reg  [31:0]         v0_283;
  reg  [31:0]         v0_284;
  reg  [31:0]         v0_285;
  reg  [31:0]         v0_286;
  reg  [31:0]         v0_287;
  reg  [31:0]         v0_288;
  reg  [31:0]         v0_289;
  reg  [31:0]         v0_290;
  reg  [31:0]         v0_291;
  reg  [31:0]         v0_292;
  reg  [31:0]         v0_293;
  reg  [31:0]         v0_294;
  reg  [31:0]         v0_295;
  reg  [31:0]         v0_296;
  reg  [31:0]         v0_297;
  reg  [31:0]         v0_298;
  reg  [31:0]         v0_299;
  reg  [31:0]         v0_300;
  reg  [31:0]         v0_301;
  reg  [31:0]         v0_302;
  reg  [31:0]         v0_303;
  reg  [31:0]         v0_304;
  reg  [31:0]         v0_305;
  reg  [31:0]         v0_306;
  reg  [31:0]         v0_307;
  reg  [31:0]         v0_308;
  reg  [31:0]         v0_309;
  reg  [31:0]         v0_310;
  reg  [31:0]         v0_311;
  reg  [31:0]         v0_312;
  reg  [31:0]         v0_313;
  reg  [31:0]         v0_314;
  reg  [31:0]         v0_315;
  reg  [31:0]         v0_316;
  reg  [31:0]         v0_317;
  reg  [31:0]         v0_318;
  reg  [31:0]         v0_319;
  reg  [31:0]         v0_320;
  reg  [31:0]         v0_321;
  reg  [31:0]         v0_322;
  reg  [31:0]         v0_323;
  reg  [31:0]         v0_324;
  reg  [31:0]         v0_325;
  reg  [31:0]         v0_326;
  reg  [31:0]         v0_327;
  reg  [31:0]         v0_328;
  reg  [31:0]         v0_329;
  reg  [31:0]         v0_330;
  reg  [31:0]         v0_331;
  reg  [31:0]         v0_332;
  reg  [31:0]         v0_333;
  reg  [31:0]         v0_334;
  reg  [31:0]         v0_335;
  reg  [31:0]         v0_336;
  reg  [31:0]         v0_337;
  reg  [31:0]         v0_338;
  reg  [31:0]         v0_339;
  reg  [31:0]         v0_340;
  reg  [31:0]         v0_341;
  reg  [31:0]         v0_342;
  reg  [31:0]         v0_343;
  reg  [31:0]         v0_344;
  reg  [31:0]         v0_345;
  reg  [31:0]         v0_346;
  reg  [31:0]         v0_347;
  reg  [31:0]         v0_348;
  reg  [31:0]         v0_349;
  reg  [31:0]         v0_350;
  reg  [31:0]         v0_351;
  reg  [31:0]         v0_352;
  reg  [31:0]         v0_353;
  reg  [31:0]         v0_354;
  reg  [31:0]         v0_355;
  reg  [31:0]         v0_356;
  reg  [31:0]         v0_357;
  reg  [31:0]         v0_358;
  reg  [31:0]         v0_359;
  reg  [31:0]         v0_360;
  reg  [31:0]         v0_361;
  reg  [31:0]         v0_362;
  reg  [31:0]         v0_363;
  reg  [31:0]         v0_364;
  reg  [31:0]         v0_365;
  reg  [31:0]         v0_366;
  reg  [31:0]         v0_367;
  reg  [31:0]         v0_368;
  reg  [31:0]         v0_369;
  reg  [31:0]         v0_370;
  reg  [31:0]         v0_371;
  reg  [31:0]         v0_372;
  reg  [31:0]         v0_373;
  reg  [31:0]         v0_374;
  reg  [31:0]         v0_375;
  reg  [31:0]         v0_376;
  reg  [31:0]         v0_377;
  reg  [31:0]         v0_378;
  reg  [31:0]         v0_379;
  reg  [31:0]         v0_380;
  reg  [31:0]         v0_381;
  reg  [31:0]         v0_382;
  reg  [31:0]         v0_383;
  reg  [31:0]         v0_384;
  reg  [31:0]         v0_385;
  reg  [31:0]         v0_386;
  reg  [31:0]         v0_387;
  reg  [31:0]         v0_388;
  reg  [31:0]         v0_389;
  reg  [31:0]         v0_390;
  reg  [31:0]         v0_391;
  reg  [31:0]         v0_392;
  reg  [31:0]         v0_393;
  reg  [31:0]         v0_394;
  reg  [31:0]         v0_395;
  reg  [31:0]         v0_396;
  reg  [31:0]         v0_397;
  reg  [31:0]         v0_398;
  reg  [31:0]         v0_399;
  reg  [31:0]         v0_400;
  reg  [31:0]         v0_401;
  reg  [31:0]         v0_402;
  reg  [31:0]         v0_403;
  reg  [31:0]         v0_404;
  reg  [31:0]         v0_405;
  reg  [31:0]         v0_406;
  reg  [31:0]         v0_407;
  reg  [31:0]         v0_408;
  reg  [31:0]         v0_409;
  reg  [31:0]         v0_410;
  reg  [31:0]         v0_411;
  reg  [31:0]         v0_412;
  reg  [31:0]         v0_413;
  reg  [31:0]         v0_414;
  reg  [31:0]         v0_415;
  reg  [31:0]         v0_416;
  reg  [31:0]         v0_417;
  reg  [31:0]         v0_418;
  reg  [31:0]         v0_419;
  reg  [31:0]         v0_420;
  reg  [31:0]         v0_421;
  reg  [31:0]         v0_422;
  reg  [31:0]         v0_423;
  reg  [31:0]         v0_424;
  reg  [31:0]         v0_425;
  reg  [31:0]         v0_426;
  reg  [31:0]         v0_427;
  reg  [31:0]         v0_428;
  reg  [31:0]         v0_429;
  reg  [31:0]         v0_430;
  reg  [31:0]         v0_431;
  reg  [31:0]         v0_432;
  reg  [31:0]         v0_433;
  reg  [31:0]         v0_434;
  reg  [31:0]         v0_435;
  reg  [31:0]         v0_436;
  reg  [31:0]         v0_437;
  reg  [31:0]         v0_438;
  reg  [31:0]         v0_439;
  reg  [31:0]         v0_440;
  reg  [31:0]         v0_441;
  reg  [31:0]         v0_442;
  reg  [31:0]         v0_443;
  reg  [31:0]         v0_444;
  reg  [31:0]         v0_445;
  reg  [31:0]         v0_446;
  reg  [31:0]         v0_447;
  reg  [31:0]         v0_448;
  reg  [31:0]         v0_449;
  reg  [31:0]         v0_450;
  reg  [31:0]         v0_451;
  reg  [31:0]         v0_452;
  reg  [31:0]         v0_453;
  reg  [31:0]         v0_454;
  reg  [31:0]         v0_455;
  reg  [31:0]         v0_456;
  reg  [31:0]         v0_457;
  reg  [31:0]         v0_458;
  reg  [31:0]         v0_459;
  reg  [31:0]         v0_460;
  reg  [31:0]         v0_461;
  reg  [31:0]         v0_462;
  reg  [31:0]         v0_463;
  reg  [31:0]         v0_464;
  reg  [31:0]         v0_465;
  reg  [31:0]         v0_466;
  reg  [31:0]         v0_467;
  reg  [31:0]         v0_468;
  reg  [31:0]         v0_469;
  reg  [31:0]         v0_470;
  reg  [31:0]         v0_471;
  reg  [31:0]         v0_472;
  reg  [31:0]         v0_473;
  reg  [31:0]         v0_474;
  reg  [31:0]         v0_475;
  reg  [31:0]         v0_476;
  reg  [31:0]         v0_477;
  reg  [31:0]         v0_478;
  reg  [31:0]         v0_479;
  reg  [31:0]         v0_480;
  reg  [31:0]         v0_481;
  reg  [31:0]         v0_482;
  reg  [31:0]         v0_483;
  reg  [31:0]         v0_484;
  reg  [31:0]         v0_485;
  reg  [31:0]         v0_486;
  reg  [31:0]         v0_487;
  reg  [31:0]         v0_488;
  reg  [31:0]         v0_489;
  reg  [31:0]         v0_490;
  reg  [31:0]         v0_491;
  reg  [31:0]         v0_492;
  reg  [31:0]         v0_493;
  reg  [31:0]         v0_494;
  reg  [31:0]         v0_495;
  reg  [31:0]         v0_496;
  reg  [31:0]         v0_497;
  reg  [31:0]         v0_498;
  reg  [31:0]         v0_499;
  reg  [31:0]         v0_500;
  reg  [31:0]         v0_501;
  reg  [31:0]         v0_502;
  reg  [31:0]         v0_503;
  reg  [31:0]         v0_504;
  reg  [31:0]         v0_505;
  reg  [31:0]         v0_506;
  reg  [31:0]         v0_507;
  reg  [31:0]         v0_508;
  reg  [31:0]         v0_509;
  reg  [31:0]         v0_510;
  reg  [31:0]         v0_511;
  reg  [31:0]         v0_512;
  reg  [31:0]         v0_513;
  reg  [31:0]         v0_514;
  reg  [31:0]         v0_515;
  reg  [31:0]         v0_516;
  reg  [31:0]         v0_517;
  reg  [31:0]         v0_518;
  reg  [31:0]         v0_519;
  reg  [31:0]         v0_520;
  reg  [31:0]         v0_521;
  reg  [31:0]         v0_522;
  reg  [31:0]         v0_523;
  reg  [31:0]         v0_524;
  reg  [31:0]         v0_525;
  reg  [31:0]         v0_526;
  reg  [31:0]         v0_527;
  reg  [31:0]         v0_528;
  reg  [31:0]         v0_529;
  reg  [31:0]         v0_530;
  reg  [31:0]         v0_531;
  reg  [31:0]         v0_532;
  reg  [31:0]         v0_533;
  reg  [31:0]         v0_534;
  reg  [31:0]         v0_535;
  reg  [31:0]         v0_536;
  reg  [31:0]         v0_537;
  reg  [31:0]         v0_538;
  reg  [31:0]         v0_539;
  reg  [31:0]         v0_540;
  reg  [31:0]         v0_541;
  reg  [31:0]         v0_542;
  reg  [31:0]         v0_543;
  reg  [31:0]         v0_544;
  reg  [31:0]         v0_545;
  reg  [31:0]         v0_546;
  reg  [31:0]         v0_547;
  reg  [31:0]         v0_548;
  reg  [31:0]         v0_549;
  reg  [31:0]         v0_550;
  reg  [31:0]         v0_551;
  reg  [31:0]         v0_552;
  reg  [31:0]         v0_553;
  reg  [31:0]         v0_554;
  reg  [31:0]         v0_555;
  reg  [31:0]         v0_556;
  reg  [31:0]         v0_557;
  reg  [31:0]         v0_558;
  reg  [31:0]         v0_559;
  reg  [31:0]         v0_560;
  reg  [31:0]         v0_561;
  reg  [31:0]         v0_562;
  reg  [31:0]         v0_563;
  reg  [31:0]         v0_564;
  reg  [31:0]         v0_565;
  reg  [31:0]         v0_566;
  reg  [31:0]         v0_567;
  reg  [31:0]         v0_568;
  reg  [31:0]         v0_569;
  reg  [31:0]         v0_570;
  reg  [31:0]         v0_571;
  reg  [31:0]         v0_572;
  reg  [31:0]         v0_573;
  reg  [31:0]         v0_574;
  reg  [31:0]         v0_575;
  reg  [31:0]         v0_576;
  reg  [31:0]         v0_577;
  reg  [31:0]         v0_578;
  reg  [31:0]         v0_579;
  reg  [31:0]         v0_580;
  reg  [31:0]         v0_581;
  reg  [31:0]         v0_582;
  reg  [31:0]         v0_583;
  reg  [31:0]         v0_584;
  reg  [31:0]         v0_585;
  reg  [31:0]         v0_586;
  reg  [31:0]         v0_587;
  reg  [31:0]         v0_588;
  reg  [31:0]         v0_589;
  reg  [31:0]         v0_590;
  reg  [31:0]         v0_591;
  reg  [31:0]         v0_592;
  reg  [31:0]         v0_593;
  reg  [31:0]         v0_594;
  reg  [31:0]         v0_595;
  reg  [31:0]         v0_596;
  reg  [31:0]         v0_597;
  reg  [31:0]         v0_598;
  reg  [31:0]         v0_599;
  reg  [31:0]         v0_600;
  reg  [31:0]         v0_601;
  reg  [31:0]         v0_602;
  reg  [31:0]         v0_603;
  reg  [31:0]         v0_604;
  reg  [31:0]         v0_605;
  reg  [31:0]         v0_606;
  reg  [31:0]         v0_607;
  reg  [31:0]         v0_608;
  reg  [31:0]         v0_609;
  reg  [31:0]         v0_610;
  reg  [31:0]         v0_611;
  reg  [31:0]         v0_612;
  reg  [31:0]         v0_613;
  reg  [31:0]         v0_614;
  reg  [31:0]         v0_615;
  reg  [31:0]         v0_616;
  reg  [31:0]         v0_617;
  reg  [31:0]         v0_618;
  reg  [31:0]         v0_619;
  reg  [31:0]         v0_620;
  reg  [31:0]         v0_621;
  reg  [31:0]         v0_622;
  reg  [31:0]         v0_623;
  reg  [31:0]         v0_624;
  reg  [31:0]         v0_625;
  reg  [31:0]         v0_626;
  reg  [31:0]         v0_627;
  reg  [31:0]         v0_628;
  reg  [31:0]         v0_629;
  reg  [31:0]         v0_630;
  reg  [31:0]         v0_631;
  reg  [31:0]         v0_632;
  reg  [31:0]         v0_633;
  reg  [31:0]         v0_634;
  reg  [31:0]         v0_635;
  reg  [31:0]         v0_636;
  reg  [31:0]         v0_637;
  reg  [31:0]         v0_638;
  reg  [31:0]         v0_639;
  reg  [31:0]         v0_640;
  reg  [31:0]         v0_641;
  reg  [31:0]         v0_642;
  reg  [31:0]         v0_643;
  reg  [31:0]         v0_644;
  reg  [31:0]         v0_645;
  reg  [31:0]         v0_646;
  reg  [31:0]         v0_647;
  reg  [31:0]         v0_648;
  reg  [31:0]         v0_649;
  reg  [31:0]         v0_650;
  reg  [31:0]         v0_651;
  reg  [31:0]         v0_652;
  reg  [31:0]         v0_653;
  reg  [31:0]         v0_654;
  reg  [31:0]         v0_655;
  reg  [31:0]         v0_656;
  reg  [31:0]         v0_657;
  reg  [31:0]         v0_658;
  reg  [31:0]         v0_659;
  reg  [31:0]         v0_660;
  reg  [31:0]         v0_661;
  reg  [31:0]         v0_662;
  reg  [31:0]         v0_663;
  reg  [31:0]         v0_664;
  reg  [31:0]         v0_665;
  reg  [31:0]         v0_666;
  reg  [31:0]         v0_667;
  reg  [31:0]         v0_668;
  reg  [31:0]         v0_669;
  reg  [31:0]         v0_670;
  reg  [31:0]         v0_671;
  reg  [31:0]         v0_672;
  reg  [31:0]         v0_673;
  reg  [31:0]         v0_674;
  reg  [31:0]         v0_675;
  reg  [31:0]         v0_676;
  reg  [31:0]         v0_677;
  reg  [31:0]         v0_678;
  reg  [31:0]         v0_679;
  reg  [31:0]         v0_680;
  reg  [31:0]         v0_681;
  reg  [31:0]         v0_682;
  reg  [31:0]         v0_683;
  reg  [31:0]         v0_684;
  reg  [31:0]         v0_685;
  reg  [31:0]         v0_686;
  reg  [31:0]         v0_687;
  reg  [31:0]         v0_688;
  reg  [31:0]         v0_689;
  reg  [31:0]         v0_690;
  reg  [31:0]         v0_691;
  reg  [31:0]         v0_692;
  reg  [31:0]         v0_693;
  reg  [31:0]         v0_694;
  reg  [31:0]         v0_695;
  reg  [31:0]         v0_696;
  reg  [31:0]         v0_697;
  reg  [31:0]         v0_698;
  reg  [31:0]         v0_699;
  reg  [31:0]         v0_700;
  reg  [31:0]         v0_701;
  reg  [31:0]         v0_702;
  reg  [31:0]         v0_703;
  reg  [31:0]         v0_704;
  reg  [31:0]         v0_705;
  reg  [31:0]         v0_706;
  reg  [31:0]         v0_707;
  reg  [31:0]         v0_708;
  reg  [31:0]         v0_709;
  reg  [31:0]         v0_710;
  reg  [31:0]         v0_711;
  reg  [31:0]         v0_712;
  reg  [31:0]         v0_713;
  reg  [31:0]         v0_714;
  reg  [31:0]         v0_715;
  reg  [31:0]         v0_716;
  reg  [31:0]         v0_717;
  reg  [31:0]         v0_718;
  reg  [31:0]         v0_719;
  reg  [31:0]         v0_720;
  reg  [31:0]         v0_721;
  reg  [31:0]         v0_722;
  reg  [31:0]         v0_723;
  reg  [31:0]         v0_724;
  reg  [31:0]         v0_725;
  reg  [31:0]         v0_726;
  reg  [31:0]         v0_727;
  reg  [31:0]         v0_728;
  reg  [31:0]         v0_729;
  reg  [31:0]         v0_730;
  reg  [31:0]         v0_731;
  reg  [31:0]         v0_732;
  reg  [31:0]         v0_733;
  reg  [31:0]         v0_734;
  reg  [31:0]         v0_735;
  reg  [31:0]         v0_736;
  reg  [31:0]         v0_737;
  reg  [31:0]         v0_738;
  reg  [31:0]         v0_739;
  reg  [31:0]         v0_740;
  reg  [31:0]         v0_741;
  reg  [31:0]         v0_742;
  reg  [31:0]         v0_743;
  reg  [31:0]         v0_744;
  reg  [31:0]         v0_745;
  reg  [31:0]         v0_746;
  reg  [31:0]         v0_747;
  reg  [31:0]         v0_748;
  reg  [31:0]         v0_749;
  reg  [31:0]         v0_750;
  reg  [31:0]         v0_751;
  reg  [31:0]         v0_752;
  reg  [31:0]         v0_753;
  reg  [31:0]         v0_754;
  reg  [31:0]         v0_755;
  reg  [31:0]         v0_756;
  reg  [31:0]         v0_757;
  reg  [31:0]         v0_758;
  reg  [31:0]         v0_759;
  reg  [31:0]         v0_760;
  reg  [31:0]         v0_761;
  reg  [31:0]         v0_762;
  reg  [31:0]         v0_763;
  reg  [31:0]         v0_764;
  reg  [31:0]         v0_765;
  reg  [31:0]         v0_766;
  reg  [31:0]         v0_767;
  reg  [31:0]         v0_768;
  reg  [31:0]         v0_769;
  reg  [31:0]         v0_770;
  reg  [31:0]         v0_771;
  reg  [31:0]         v0_772;
  reg  [31:0]         v0_773;
  reg  [31:0]         v0_774;
  reg  [31:0]         v0_775;
  reg  [31:0]         v0_776;
  reg  [31:0]         v0_777;
  reg  [31:0]         v0_778;
  reg  [31:0]         v0_779;
  reg  [31:0]         v0_780;
  reg  [31:0]         v0_781;
  reg  [31:0]         v0_782;
  reg  [31:0]         v0_783;
  reg  [31:0]         v0_784;
  reg  [31:0]         v0_785;
  reg  [31:0]         v0_786;
  reg  [31:0]         v0_787;
  reg  [31:0]         v0_788;
  reg  [31:0]         v0_789;
  reg  [31:0]         v0_790;
  reg  [31:0]         v0_791;
  reg  [31:0]         v0_792;
  reg  [31:0]         v0_793;
  reg  [31:0]         v0_794;
  reg  [31:0]         v0_795;
  reg  [31:0]         v0_796;
  reg  [31:0]         v0_797;
  reg  [31:0]         v0_798;
  reg  [31:0]         v0_799;
  reg  [31:0]         v0_800;
  reg  [31:0]         v0_801;
  reg  [31:0]         v0_802;
  reg  [31:0]         v0_803;
  reg  [31:0]         v0_804;
  reg  [31:0]         v0_805;
  reg  [31:0]         v0_806;
  reg  [31:0]         v0_807;
  reg  [31:0]         v0_808;
  reg  [31:0]         v0_809;
  reg  [31:0]         v0_810;
  reg  [31:0]         v0_811;
  reg  [31:0]         v0_812;
  reg  [31:0]         v0_813;
  reg  [31:0]         v0_814;
  reg  [31:0]         v0_815;
  reg  [31:0]         v0_816;
  reg  [31:0]         v0_817;
  reg  [31:0]         v0_818;
  reg  [31:0]         v0_819;
  reg  [31:0]         v0_820;
  reg  [31:0]         v0_821;
  reg  [31:0]         v0_822;
  reg  [31:0]         v0_823;
  reg  [31:0]         v0_824;
  reg  [31:0]         v0_825;
  reg  [31:0]         v0_826;
  reg  [31:0]         v0_827;
  reg  [31:0]         v0_828;
  reg  [31:0]         v0_829;
  reg  [31:0]         v0_830;
  reg  [31:0]         v0_831;
  reg  [31:0]         v0_832;
  reg  [31:0]         v0_833;
  reg  [31:0]         v0_834;
  reg  [31:0]         v0_835;
  reg  [31:0]         v0_836;
  reg  [31:0]         v0_837;
  reg  [31:0]         v0_838;
  reg  [31:0]         v0_839;
  reg  [31:0]         v0_840;
  reg  [31:0]         v0_841;
  reg  [31:0]         v0_842;
  reg  [31:0]         v0_843;
  reg  [31:0]         v0_844;
  reg  [31:0]         v0_845;
  reg  [31:0]         v0_846;
  reg  [31:0]         v0_847;
  reg  [31:0]         v0_848;
  reg  [31:0]         v0_849;
  reg  [31:0]         v0_850;
  reg  [31:0]         v0_851;
  reg  [31:0]         v0_852;
  reg  [31:0]         v0_853;
  reg  [31:0]         v0_854;
  reg  [31:0]         v0_855;
  reg  [31:0]         v0_856;
  reg  [31:0]         v0_857;
  reg  [31:0]         v0_858;
  reg  [31:0]         v0_859;
  reg  [31:0]         v0_860;
  reg  [31:0]         v0_861;
  reg  [31:0]         v0_862;
  reg  [31:0]         v0_863;
  reg  [31:0]         v0_864;
  reg  [31:0]         v0_865;
  reg  [31:0]         v0_866;
  reg  [31:0]         v0_867;
  reg  [31:0]         v0_868;
  reg  [31:0]         v0_869;
  reg  [31:0]         v0_870;
  reg  [31:0]         v0_871;
  reg  [31:0]         v0_872;
  reg  [31:0]         v0_873;
  reg  [31:0]         v0_874;
  reg  [31:0]         v0_875;
  reg  [31:0]         v0_876;
  reg  [31:0]         v0_877;
  reg  [31:0]         v0_878;
  reg  [31:0]         v0_879;
  reg  [31:0]         v0_880;
  reg  [31:0]         v0_881;
  reg  [31:0]         v0_882;
  reg  [31:0]         v0_883;
  reg  [31:0]         v0_884;
  reg  [31:0]         v0_885;
  reg  [31:0]         v0_886;
  reg  [31:0]         v0_887;
  reg  [31:0]         v0_888;
  reg  [31:0]         v0_889;
  reg  [31:0]         v0_890;
  reg  [31:0]         v0_891;
  reg  [31:0]         v0_892;
  reg  [31:0]         v0_893;
  reg  [31:0]         v0_894;
  reg  [31:0]         v0_895;
  reg  [31:0]         v0_896;
  reg  [31:0]         v0_897;
  reg  [31:0]         v0_898;
  reg  [31:0]         v0_899;
  reg  [31:0]         v0_900;
  reg  [31:0]         v0_901;
  reg  [31:0]         v0_902;
  reg  [31:0]         v0_903;
  reg  [31:0]         v0_904;
  reg  [31:0]         v0_905;
  reg  [31:0]         v0_906;
  reg  [31:0]         v0_907;
  reg  [31:0]         v0_908;
  reg  [31:0]         v0_909;
  reg  [31:0]         v0_910;
  reg  [31:0]         v0_911;
  reg  [31:0]         v0_912;
  reg  [31:0]         v0_913;
  reg  [31:0]         v0_914;
  reg  [31:0]         v0_915;
  reg  [31:0]         v0_916;
  reg  [31:0]         v0_917;
  reg  [31:0]         v0_918;
  reg  [31:0]         v0_919;
  reg  [31:0]         v0_920;
  reg  [31:0]         v0_921;
  reg  [31:0]         v0_922;
  reg  [31:0]         v0_923;
  reg  [31:0]         v0_924;
  reg  [31:0]         v0_925;
  reg  [31:0]         v0_926;
  reg  [31:0]         v0_927;
  reg  [31:0]         v0_928;
  reg  [31:0]         v0_929;
  reg  [31:0]         v0_930;
  reg  [31:0]         v0_931;
  reg  [31:0]         v0_932;
  reg  [31:0]         v0_933;
  reg  [31:0]         v0_934;
  reg  [31:0]         v0_935;
  reg  [31:0]         v0_936;
  reg  [31:0]         v0_937;
  reg  [31:0]         v0_938;
  reg  [31:0]         v0_939;
  reg  [31:0]         v0_940;
  reg  [31:0]         v0_941;
  reg  [31:0]         v0_942;
  reg  [31:0]         v0_943;
  reg  [31:0]         v0_944;
  reg  [31:0]         v0_945;
  reg  [31:0]         v0_946;
  reg  [31:0]         v0_947;
  reg  [31:0]         v0_948;
  reg  [31:0]         v0_949;
  reg  [31:0]         v0_950;
  reg  [31:0]         v0_951;
  reg  [31:0]         v0_952;
  reg  [31:0]         v0_953;
  reg  [31:0]         v0_954;
  reg  [31:0]         v0_955;
  reg  [31:0]         v0_956;
  reg  [31:0]         v0_957;
  reg  [31:0]         v0_958;
  reg  [31:0]         v0_959;
  reg  [31:0]         v0_960;
  reg  [31:0]         v0_961;
  reg  [31:0]         v0_962;
  reg  [31:0]         v0_963;
  reg  [31:0]         v0_964;
  reg  [31:0]         v0_965;
  reg  [31:0]         v0_966;
  reg  [31:0]         v0_967;
  reg  [31:0]         v0_968;
  reg  [31:0]         v0_969;
  reg  [31:0]         v0_970;
  reg  [31:0]         v0_971;
  reg  [31:0]         v0_972;
  reg  [31:0]         v0_973;
  reg  [31:0]         v0_974;
  reg  [31:0]         v0_975;
  reg  [31:0]         v0_976;
  reg  [31:0]         v0_977;
  reg  [31:0]         v0_978;
  reg  [31:0]         v0_979;
  reg  [31:0]         v0_980;
  reg  [31:0]         v0_981;
  reg  [31:0]         v0_982;
  reg  [31:0]         v0_983;
  reg  [31:0]         v0_984;
  reg  [31:0]         v0_985;
  reg  [31:0]         v0_986;
  reg  [31:0]         v0_987;
  reg  [31:0]         v0_988;
  reg  [31:0]         v0_989;
  reg  [31:0]         v0_990;
  reg  [31:0]         v0_991;
  reg  [31:0]         v0_992;
  reg  [31:0]         v0_993;
  reg  [31:0]         v0_994;
  reg  [31:0]         v0_995;
  reg  [31:0]         v0_996;
  reg  [31:0]         v0_997;
  reg  [31:0]         v0_998;
  reg  [31:0]         v0_999;
  reg  [31:0]         v0_1000;
  reg  [31:0]         v0_1001;
  reg  [31:0]         v0_1002;
  reg  [31:0]         v0_1003;
  reg  [31:0]         v0_1004;
  reg  [31:0]         v0_1005;
  reg  [31:0]         v0_1006;
  reg  [31:0]         v0_1007;
  reg  [31:0]         v0_1008;
  reg  [31:0]         v0_1009;
  reg  [31:0]         v0_1010;
  reg  [31:0]         v0_1011;
  reg  [31:0]         v0_1012;
  reg  [31:0]         v0_1013;
  reg  [31:0]         v0_1014;
  reg  [31:0]         v0_1015;
  reg  [31:0]         v0_1016;
  reg  [31:0]         v0_1017;
  reg  [31:0]         v0_1018;
  reg  [31:0]         v0_1019;
  reg  [31:0]         v0_1020;
  reg  [31:0]         v0_1021;
  reg  [31:0]         v0_1022;
  reg  [31:0]         v0_1023;
  reg  [31:0]         v0_1024;
  reg  [31:0]         v0_1025;
  reg  [31:0]         v0_1026;
  reg  [31:0]         v0_1027;
  reg  [31:0]         v0_1028;
  reg  [31:0]         v0_1029;
  reg  [31:0]         v0_1030;
  reg  [31:0]         v0_1031;
  reg  [31:0]         v0_1032;
  reg  [31:0]         v0_1033;
  reg  [31:0]         v0_1034;
  reg  [31:0]         v0_1035;
  reg  [31:0]         v0_1036;
  reg  [31:0]         v0_1037;
  reg  [31:0]         v0_1038;
  reg  [31:0]         v0_1039;
  reg  [31:0]         v0_1040;
  reg  [31:0]         v0_1041;
  reg  [31:0]         v0_1042;
  reg  [31:0]         v0_1043;
  reg  [31:0]         v0_1044;
  reg  [31:0]         v0_1045;
  reg  [31:0]         v0_1046;
  reg  [31:0]         v0_1047;
  reg  [31:0]         v0_1048;
  reg  [31:0]         v0_1049;
  reg  [31:0]         v0_1050;
  reg  [31:0]         v0_1051;
  reg  [31:0]         v0_1052;
  reg  [31:0]         v0_1053;
  reg  [31:0]         v0_1054;
  reg  [31:0]         v0_1055;
  reg  [31:0]         v0_1056;
  reg  [31:0]         v0_1057;
  reg  [31:0]         v0_1058;
  reg  [31:0]         v0_1059;
  reg  [31:0]         v0_1060;
  reg  [31:0]         v0_1061;
  reg  [31:0]         v0_1062;
  reg  [31:0]         v0_1063;
  reg  [31:0]         v0_1064;
  reg  [31:0]         v0_1065;
  reg  [31:0]         v0_1066;
  reg  [31:0]         v0_1067;
  reg  [31:0]         v0_1068;
  reg  [31:0]         v0_1069;
  reg  [31:0]         v0_1070;
  reg  [31:0]         v0_1071;
  reg  [31:0]         v0_1072;
  reg  [31:0]         v0_1073;
  reg  [31:0]         v0_1074;
  reg  [31:0]         v0_1075;
  reg  [31:0]         v0_1076;
  reg  [31:0]         v0_1077;
  reg  [31:0]         v0_1078;
  reg  [31:0]         v0_1079;
  reg  [31:0]         v0_1080;
  reg  [31:0]         v0_1081;
  reg  [31:0]         v0_1082;
  reg  [31:0]         v0_1083;
  reg  [31:0]         v0_1084;
  reg  [31:0]         v0_1085;
  reg  [31:0]         v0_1086;
  reg  [31:0]         v0_1087;
  reg  [31:0]         v0_1088;
  reg  [31:0]         v0_1089;
  reg  [31:0]         v0_1090;
  reg  [31:0]         v0_1091;
  reg  [31:0]         v0_1092;
  reg  [31:0]         v0_1093;
  reg  [31:0]         v0_1094;
  reg  [31:0]         v0_1095;
  reg  [31:0]         v0_1096;
  reg  [31:0]         v0_1097;
  reg  [31:0]         v0_1098;
  reg  [31:0]         v0_1099;
  reg  [31:0]         v0_1100;
  reg  [31:0]         v0_1101;
  reg  [31:0]         v0_1102;
  reg  [31:0]         v0_1103;
  reg  [31:0]         v0_1104;
  reg  [31:0]         v0_1105;
  reg  [31:0]         v0_1106;
  reg  [31:0]         v0_1107;
  reg  [31:0]         v0_1108;
  reg  [31:0]         v0_1109;
  reg  [31:0]         v0_1110;
  reg  [31:0]         v0_1111;
  reg  [31:0]         v0_1112;
  reg  [31:0]         v0_1113;
  reg  [31:0]         v0_1114;
  reg  [31:0]         v0_1115;
  reg  [31:0]         v0_1116;
  reg  [31:0]         v0_1117;
  reg  [31:0]         v0_1118;
  reg  [31:0]         v0_1119;
  reg  [31:0]         v0_1120;
  reg  [31:0]         v0_1121;
  reg  [31:0]         v0_1122;
  reg  [31:0]         v0_1123;
  reg  [31:0]         v0_1124;
  reg  [31:0]         v0_1125;
  reg  [31:0]         v0_1126;
  reg  [31:0]         v0_1127;
  reg  [31:0]         v0_1128;
  reg  [31:0]         v0_1129;
  reg  [31:0]         v0_1130;
  reg  [31:0]         v0_1131;
  reg  [31:0]         v0_1132;
  reg  [31:0]         v0_1133;
  reg  [31:0]         v0_1134;
  reg  [31:0]         v0_1135;
  reg  [31:0]         v0_1136;
  reg  [31:0]         v0_1137;
  reg  [31:0]         v0_1138;
  reg  [31:0]         v0_1139;
  reg  [31:0]         v0_1140;
  reg  [31:0]         v0_1141;
  reg  [31:0]         v0_1142;
  reg  [31:0]         v0_1143;
  reg  [31:0]         v0_1144;
  reg  [31:0]         v0_1145;
  reg  [31:0]         v0_1146;
  reg  [31:0]         v0_1147;
  reg  [31:0]         v0_1148;
  reg  [31:0]         v0_1149;
  reg  [31:0]         v0_1150;
  reg  [31:0]         v0_1151;
  reg  [31:0]         v0_1152;
  reg  [31:0]         v0_1153;
  reg  [31:0]         v0_1154;
  reg  [31:0]         v0_1155;
  reg  [31:0]         v0_1156;
  reg  [31:0]         v0_1157;
  reg  [31:0]         v0_1158;
  reg  [31:0]         v0_1159;
  reg  [31:0]         v0_1160;
  reg  [31:0]         v0_1161;
  reg  [31:0]         v0_1162;
  reg  [31:0]         v0_1163;
  reg  [31:0]         v0_1164;
  reg  [31:0]         v0_1165;
  reg  [31:0]         v0_1166;
  reg  [31:0]         v0_1167;
  reg  [31:0]         v0_1168;
  reg  [31:0]         v0_1169;
  reg  [31:0]         v0_1170;
  reg  [31:0]         v0_1171;
  reg  [31:0]         v0_1172;
  reg  [31:0]         v0_1173;
  reg  [31:0]         v0_1174;
  reg  [31:0]         v0_1175;
  reg  [31:0]         v0_1176;
  reg  [31:0]         v0_1177;
  reg  [31:0]         v0_1178;
  reg  [31:0]         v0_1179;
  reg  [31:0]         v0_1180;
  reg  [31:0]         v0_1181;
  reg  [31:0]         v0_1182;
  reg  [31:0]         v0_1183;
  reg  [31:0]         v0_1184;
  reg  [31:0]         v0_1185;
  reg  [31:0]         v0_1186;
  reg  [31:0]         v0_1187;
  reg  [31:0]         v0_1188;
  reg  [31:0]         v0_1189;
  reg  [31:0]         v0_1190;
  reg  [31:0]         v0_1191;
  reg  [31:0]         v0_1192;
  reg  [31:0]         v0_1193;
  reg  [31:0]         v0_1194;
  reg  [31:0]         v0_1195;
  reg  [31:0]         v0_1196;
  reg  [31:0]         v0_1197;
  reg  [31:0]         v0_1198;
  reg  [31:0]         v0_1199;
  reg  [31:0]         v0_1200;
  reg  [31:0]         v0_1201;
  reg  [31:0]         v0_1202;
  reg  [31:0]         v0_1203;
  reg  [31:0]         v0_1204;
  reg  [31:0]         v0_1205;
  reg  [31:0]         v0_1206;
  reg  [31:0]         v0_1207;
  reg  [31:0]         v0_1208;
  reg  [31:0]         v0_1209;
  reg  [31:0]         v0_1210;
  reg  [31:0]         v0_1211;
  reg  [31:0]         v0_1212;
  reg  [31:0]         v0_1213;
  reg  [31:0]         v0_1214;
  reg  [31:0]         v0_1215;
  reg  [31:0]         v0_1216;
  reg  [31:0]         v0_1217;
  reg  [31:0]         v0_1218;
  reg  [31:0]         v0_1219;
  reg  [31:0]         v0_1220;
  reg  [31:0]         v0_1221;
  reg  [31:0]         v0_1222;
  reg  [31:0]         v0_1223;
  reg  [31:0]         v0_1224;
  reg  [31:0]         v0_1225;
  reg  [31:0]         v0_1226;
  reg  [31:0]         v0_1227;
  reg  [31:0]         v0_1228;
  reg  [31:0]         v0_1229;
  reg  [31:0]         v0_1230;
  reg  [31:0]         v0_1231;
  reg  [31:0]         v0_1232;
  reg  [31:0]         v0_1233;
  reg  [31:0]         v0_1234;
  reg  [31:0]         v0_1235;
  reg  [31:0]         v0_1236;
  reg  [31:0]         v0_1237;
  reg  [31:0]         v0_1238;
  reg  [31:0]         v0_1239;
  reg  [31:0]         v0_1240;
  reg  [31:0]         v0_1241;
  reg  [31:0]         v0_1242;
  reg  [31:0]         v0_1243;
  reg  [31:0]         v0_1244;
  reg  [31:0]         v0_1245;
  reg  [31:0]         v0_1246;
  reg  [31:0]         v0_1247;
  reg  [31:0]         v0_1248;
  reg  [31:0]         v0_1249;
  reg  [31:0]         v0_1250;
  reg  [31:0]         v0_1251;
  reg  [31:0]         v0_1252;
  reg  [31:0]         v0_1253;
  reg  [31:0]         v0_1254;
  reg  [31:0]         v0_1255;
  reg  [31:0]         v0_1256;
  reg  [31:0]         v0_1257;
  reg  [31:0]         v0_1258;
  reg  [31:0]         v0_1259;
  reg  [31:0]         v0_1260;
  reg  [31:0]         v0_1261;
  reg  [31:0]         v0_1262;
  reg  [31:0]         v0_1263;
  reg  [31:0]         v0_1264;
  reg  [31:0]         v0_1265;
  reg  [31:0]         v0_1266;
  reg  [31:0]         v0_1267;
  reg  [31:0]         v0_1268;
  reg  [31:0]         v0_1269;
  reg  [31:0]         v0_1270;
  reg  [31:0]         v0_1271;
  reg  [31:0]         v0_1272;
  reg  [31:0]         v0_1273;
  reg  [31:0]         v0_1274;
  reg  [31:0]         v0_1275;
  reg  [31:0]         v0_1276;
  reg  [31:0]         v0_1277;
  reg  [31:0]         v0_1278;
  reg  [31:0]         v0_1279;
  reg  [31:0]         v0_1280;
  reg  [31:0]         v0_1281;
  reg  [31:0]         v0_1282;
  reg  [31:0]         v0_1283;
  reg  [31:0]         v0_1284;
  reg  [31:0]         v0_1285;
  reg  [31:0]         v0_1286;
  reg  [31:0]         v0_1287;
  reg  [31:0]         v0_1288;
  reg  [31:0]         v0_1289;
  reg  [31:0]         v0_1290;
  reg  [31:0]         v0_1291;
  reg  [31:0]         v0_1292;
  reg  [31:0]         v0_1293;
  reg  [31:0]         v0_1294;
  reg  [31:0]         v0_1295;
  reg  [31:0]         v0_1296;
  reg  [31:0]         v0_1297;
  reg  [31:0]         v0_1298;
  reg  [31:0]         v0_1299;
  reg  [31:0]         v0_1300;
  reg  [31:0]         v0_1301;
  reg  [31:0]         v0_1302;
  reg  [31:0]         v0_1303;
  reg  [31:0]         v0_1304;
  reg  [31:0]         v0_1305;
  reg  [31:0]         v0_1306;
  reg  [31:0]         v0_1307;
  reg  [31:0]         v0_1308;
  reg  [31:0]         v0_1309;
  reg  [31:0]         v0_1310;
  reg  [31:0]         v0_1311;
  reg  [31:0]         v0_1312;
  reg  [31:0]         v0_1313;
  reg  [31:0]         v0_1314;
  reg  [31:0]         v0_1315;
  reg  [31:0]         v0_1316;
  reg  [31:0]         v0_1317;
  reg  [31:0]         v0_1318;
  reg  [31:0]         v0_1319;
  reg  [31:0]         v0_1320;
  reg  [31:0]         v0_1321;
  reg  [31:0]         v0_1322;
  reg  [31:0]         v0_1323;
  reg  [31:0]         v0_1324;
  reg  [31:0]         v0_1325;
  reg  [31:0]         v0_1326;
  reg  [31:0]         v0_1327;
  reg  [31:0]         v0_1328;
  reg  [31:0]         v0_1329;
  reg  [31:0]         v0_1330;
  reg  [31:0]         v0_1331;
  reg  [31:0]         v0_1332;
  reg  [31:0]         v0_1333;
  reg  [31:0]         v0_1334;
  reg  [31:0]         v0_1335;
  reg  [31:0]         v0_1336;
  reg  [31:0]         v0_1337;
  reg  [31:0]         v0_1338;
  reg  [31:0]         v0_1339;
  reg  [31:0]         v0_1340;
  reg  [31:0]         v0_1341;
  reg  [31:0]         v0_1342;
  reg  [31:0]         v0_1343;
  reg  [31:0]         v0_1344;
  reg  [31:0]         v0_1345;
  reg  [31:0]         v0_1346;
  reg  [31:0]         v0_1347;
  reg  [31:0]         v0_1348;
  reg  [31:0]         v0_1349;
  reg  [31:0]         v0_1350;
  reg  [31:0]         v0_1351;
  reg  [31:0]         v0_1352;
  reg  [31:0]         v0_1353;
  reg  [31:0]         v0_1354;
  reg  [31:0]         v0_1355;
  reg  [31:0]         v0_1356;
  reg  [31:0]         v0_1357;
  reg  [31:0]         v0_1358;
  reg  [31:0]         v0_1359;
  reg  [31:0]         v0_1360;
  reg  [31:0]         v0_1361;
  reg  [31:0]         v0_1362;
  reg  [31:0]         v0_1363;
  reg  [31:0]         v0_1364;
  reg  [31:0]         v0_1365;
  reg  [31:0]         v0_1366;
  reg  [31:0]         v0_1367;
  reg  [31:0]         v0_1368;
  reg  [31:0]         v0_1369;
  reg  [31:0]         v0_1370;
  reg  [31:0]         v0_1371;
  reg  [31:0]         v0_1372;
  reg  [31:0]         v0_1373;
  reg  [31:0]         v0_1374;
  reg  [31:0]         v0_1375;
  reg  [31:0]         v0_1376;
  reg  [31:0]         v0_1377;
  reg  [31:0]         v0_1378;
  reg  [31:0]         v0_1379;
  reg  [31:0]         v0_1380;
  reg  [31:0]         v0_1381;
  reg  [31:0]         v0_1382;
  reg  [31:0]         v0_1383;
  reg  [31:0]         v0_1384;
  reg  [31:0]         v0_1385;
  reg  [31:0]         v0_1386;
  reg  [31:0]         v0_1387;
  reg  [31:0]         v0_1388;
  reg  [31:0]         v0_1389;
  reg  [31:0]         v0_1390;
  reg  [31:0]         v0_1391;
  reg  [31:0]         v0_1392;
  reg  [31:0]         v0_1393;
  reg  [31:0]         v0_1394;
  reg  [31:0]         v0_1395;
  reg  [31:0]         v0_1396;
  reg  [31:0]         v0_1397;
  reg  [31:0]         v0_1398;
  reg  [31:0]         v0_1399;
  reg  [31:0]         v0_1400;
  reg  [31:0]         v0_1401;
  reg  [31:0]         v0_1402;
  reg  [31:0]         v0_1403;
  reg  [31:0]         v0_1404;
  reg  [31:0]         v0_1405;
  reg  [31:0]         v0_1406;
  reg  [31:0]         v0_1407;
  reg  [31:0]         v0_1408;
  reg  [31:0]         v0_1409;
  reg  [31:0]         v0_1410;
  reg  [31:0]         v0_1411;
  reg  [31:0]         v0_1412;
  reg  [31:0]         v0_1413;
  reg  [31:0]         v0_1414;
  reg  [31:0]         v0_1415;
  reg  [31:0]         v0_1416;
  reg  [31:0]         v0_1417;
  reg  [31:0]         v0_1418;
  reg  [31:0]         v0_1419;
  reg  [31:0]         v0_1420;
  reg  [31:0]         v0_1421;
  reg  [31:0]         v0_1422;
  reg  [31:0]         v0_1423;
  reg  [31:0]         v0_1424;
  reg  [31:0]         v0_1425;
  reg  [31:0]         v0_1426;
  reg  [31:0]         v0_1427;
  reg  [31:0]         v0_1428;
  reg  [31:0]         v0_1429;
  reg  [31:0]         v0_1430;
  reg  [31:0]         v0_1431;
  reg  [31:0]         v0_1432;
  reg  [31:0]         v0_1433;
  reg  [31:0]         v0_1434;
  reg  [31:0]         v0_1435;
  reg  [31:0]         v0_1436;
  reg  [31:0]         v0_1437;
  reg  [31:0]         v0_1438;
  reg  [31:0]         v0_1439;
  reg  [31:0]         v0_1440;
  reg  [31:0]         v0_1441;
  reg  [31:0]         v0_1442;
  reg  [31:0]         v0_1443;
  reg  [31:0]         v0_1444;
  reg  [31:0]         v0_1445;
  reg  [31:0]         v0_1446;
  reg  [31:0]         v0_1447;
  reg  [31:0]         v0_1448;
  reg  [31:0]         v0_1449;
  reg  [31:0]         v0_1450;
  reg  [31:0]         v0_1451;
  reg  [31:0]         v0_1452;
  reg  [31:0]         v0_1453;
  reg  [31:0]         v0_1454;
  reg  [31:0]         v0_1455;
  reg  [31:0]         v0_1456;
  reg  [31:0]         v0_1457;
  reg  [31:0]         v0_1458;
  reg  [31:0]         v0_1459;
  reg  [31:0]         v0_1460;
  reg  [31:0]         v0_1461;
  reg  [31:0]         v0_1462;
  reg  [31:0]         v0_1463;
  reg  [31:0]         v0_1464;
  reg  [31:0]         v0_1465;
  reg  [31:0]         v0_1466;
  reg  [31:0]         v0_1467;
  reg  [31:0]         v0_1468;
  reg  [31:0]         v0_1469;
  reg  [31:0]         v0_1470;
  reg  [31:0]         v0_1471;
  reg  [31:0]         v0_1472;
  reg  [31:0]         v0_1473;
  reg  [31:0]         v0_1474;
  reg  [31:0]         v0_1475;
  reg  [31:0]         v0_1476;
  reg  [31:0]         v0_1477;
  reg  [31:0]         v0_1478;
  reg  [31:0]         v0_1479;
  reg  [31:0]         v0_1480;
  reg  [31:0]         v0_1481;
  reg  [31:0]         v0_1482;
  reg  [31:0]         v0_1483;
  reg  [31:0]         v0_1484;
  reg  [31:0]         v0_1485;
  reg  [31:0]         v0_1486;
  reg  [31:0]         v0_1487;
  reg  [31:0]         v0_1488;
  reg  [31:0]         v0_1489;
  reg  [31:0]         v0_1490;
  reg  [31:0]         v0_1491;
  reg  [31:0]         v0_1492;
  reg  [31:0]         v0_1493;
  reg  [31:0]         v0_1494;
  reg  [31:0]         v0_1495;
  reg  [31:0]         v0_1496;
  reg  [31:0]         v0_1497;
  reg  [31:0]         v0_1498;
  reg  [31:0]         v0_1499;
  reg  [31:0]         v0_1500;
  reg  [31:0]         v0_1501;
  reg  [31:0]         v0_1502;
  reg  [31:0]         v0_1503;
  reg  [31:0]         v0_1504;
  reg  [31:0]         v0_1505;
  reg  [31:0]         v0_1506;
  reg  [31:0]         v0_1507;
  reg  [31:0]         v0_1508;
  reg  [31:0]         v0_1509;
  reg  [31:0]         v0_1510;
  reg  [31:0]         v0_1511;
  reg  [31:0]         v0_1512;
  reg  [31:0]         v0_1513;
  reg  [31:0]         v0_1514;
  reg  [31:0]         v0_1515;
  reg  [31:0]         v0_1516;
  reg  [31:0]         v0_1517;
  reg  [31:0]         v0_1518;
  reg  [31:0]         v0_1519;
  reg  [31:0]         v0_1520;
  reg  [31:0]         v0_1521;
  reg  [31:0]         v0_1522;
  reg  [31:0]         v0_1523;
  reg  [31:0]         v0_1524;
  reg  [31:0]         v0_1525;
  reg  [31:0]         v0_1526;
  reg  [31:0]         v0_1527;
  reg  [31:0]         v0_1528;
  reg  [31:0]         v0_1529;
  reg  [31:0]         v0_1530;
  reg  [31:0]         v0_1531;
  reg  [31:0]         v0_1532;
  reg  [31:0]         v0_1533;
  reg  [31:0]         v0_1534;
  reg  [31:0]         v0_1535;
  reg  [31:0]         v0_1536;
  reg  [31:0]         v0_1537;
  reg  [31:0]         v0_1538;
  reg  [31:0]         v0_1539;
  reg  [31:0]         v0_1540;
  reg  [31:0]         v0_1541;
  reg  [31:0]         v0_1542;
  reg  [31:0]         v0_1543;
  reg  [31:0]         v0_1544;
  reg  [31:0]         v0_1545;
  reg  [31:0]         v0_1546;
  reg  [31:0]         v0_1547;
  reg  [31:0]         v0_1548;
  reg  [31:0]         v0_1549;
  reg  [31:0]         v0_1550;
  reg  [31:0]         v0_1551;
  reg  [31:0]         v0_1552;
  reg  [31:0]         v0_1553;
  reg  [31:0]         v0_1554;
  reg  [31:0]         v0_1555;
  reg  [31:0]         v0_1556;
  reg  [31:0]         v0_1557;
  reg  [31:0]         v0_1558;
  reg  [31:0]         v0_1559;
  reg  [31:0]         v0_1560;
  reg  [31:0]         v0_1561;
  reg  [31:0]         v0_1562;
  reg  [31:0]         v0_1563;
  reg  [31:0]         v0_1564;
  reg  [31:0]         v0_1565;
  reg  [31:0]         v0_1566;
  reg  [31:0]         v0_1567;
  reg  [31:0]         v0_1568;
  reg  [31:0]         v0_1569;
  reg  [31:0]         v0_1570;
  reg  [31:0]         v0_1571;
  reg  [31:0]         v0_1572;
  reg  [31:0]         v0_1573;
  reg  [31:0]         v0_1574;
  reg  [31:0]         v0_1575;
  reg  [31:0]         v0_1576;
  reg  [31:0]         v0_1577;
  reg  [31:0]         v0_1578;
  reg  [31:0]         v0_1579;
  reg  [31:0]         v0_1580;
  reg  [31:0]         v0_1581;
  reg  [31:0]         v0_1582;
  reg  [31:0]         v0_1583;
  reg  [31:0]         v0_1584;
  reg  [31:0]         v0_1585;
  reg  [31:0]         v0_1586;
  reg  [31:0]         v0_1587;
  reg  [31:0]         v0_1588;
  reg  [31:0]         v0_1589;
  reg  [31:0]         v0_1590;
  reg  [31:0]         v0_1591;
  reg  [31:0]         v0_1592;
  reg  [31:0]         v0_1593;
  reg  [31:0]         v0_1594;
  reg  [31:0]         v0_1595;
  reg  [31:0]         v0_1596;
  reg  [31:0]         v0_1597;
  reg  [31:0]         v0_1598;
  reg  [31:0]         v0_1599;
  reg  [31:0]         v0_1600;
  reg  [31:0]         v0_1601;
  reg  [31:0]         v0_1602;
  reg  [31:0]         v0_1603;
  reg  [31:0]         v0_1604;
  reg  [31:0]         v0_1605;
  reg  [31:0]         v0_1606;
  reg  [31:0]         v0_1607;
  reg  [31:0]         v0_1608;
  reg  [31:0]         v0_1609;
  reg  [31:0]         v0_1610;
  reg  [31:0]         v0_1611;
  reg  [31:0]         v0_1612;
  reg  [31:0]         v0_1613;
  reg  [31:0]         v0_1614;
  reg  [31:0]         v0_1615;
  reg  [31:0]         v0_1616;
  reg  [31:0]         v0_1617;
  reg  [31:0]         v0_1618;
  reg  [31:0]         v0_1619;
  reg  [31:0]         v0_1620;
  reg  [31:0]         v0_1621;
  reg  [31:0]         v0_1622;
  reg  [31:0]         v0_1623;
  reg  [31:0]         v0_1624;
  reg  [31:0]         v0_1625;
  reg  [31:0]         v0_1626;
  reg  [31:0]         v0_1627;
  reg  [31:0]         v0_1628;
  reg  [31:0]         v0_1629;
  reg  [31:0]         v0_1630;
  reg  [31:0]         v0_1631;
  reg  [31:0]         v0_1632;
  reg  [31:0]         v0_1633;
  reg  [31:0]         v0_1634;
  reg  [31:0]         v0_1635;
  reg  [31:0]         v0_1636;
  reg  [31:0]         v0_1637;
  reg  [31:0]         v0_1638;
  reg  [31:0]         v0_1639;
  reg  [31:0]         v0_1640;
  reg  [31:0]         v0_1641;
  reg  [31:0]         v0_1642;
  reg  [31:0]         v0_1643;
  reg  [31:0]         v0_1644;
  reg  [31:0]         v0_1645;
  reg  [31:0]         v0_1646;
  reg  [31:0]         v0_1647;
  reg  [31:0]         v0_1648;
  reg  [31:0]         v0_1649;
  reg  [31:0]         v0_1650;
  reg  [31:0]         v0_1651;
  reg  [31:0]         v0_1652;
  reg  [31:0]         v0_1653;
  reg  [31:0]         v0_1654;
  reg  [31:0]         v0_1655;
  reg  [31:0]         v0_1656;
  reg  [31:0]         v0_1657;
  reg  [31:0]         v0_1658;
  reg  [31:0]         v0_1659;
  reg  [31:0]         v0_1660;
  reg  [31:0]         v0_1661;
  reg  [31:0]         v0_1662;
  reg  [31:0]         v0_1663;
  reg  [31:0]         v0_1664;
  reg  [31:0]         v0_1665;
  reg  [31:0]         v0_1666;
  reg  [31:0]         v0_1667;
  reg  [31:0]         v0_1668;
  reg  [31:0]         v0_1669;
  reg  [31:0]         v0_1670;
  reg  [31:0]         v0_1671;
  reg  [31:0]         v0_1672;
  reg  [31:0]         v0_1673;
  reg  [31:0]         v0_1674;
  reg  [31:0]         v0_1675;
  reg  [31:0]         v0_1676;
  reg  [31:0]         v0_1677;
  reg  [31:0]         v0_1678;
  reg  [31:0]         v0_1679;
  reg  [31:0]         v0_1680;
  reg  [31:0]         v0_1681;
  reg  [31:0]         v0_1682;
  reg  [31:0]         v0_1683;
  reg  [31:0]         v0_1684;
  reg  [31:0]         v0_1685;
  reg  [31:0]         v0_1686;
  reg  [31:0]         v0_1687;
  reg  [31:0]         v0_1688;
  reg  [31:0]         v0_1689;
  reg  [31:0]         v0_1690;
  reg  [31:0]         v0_1691;
  reg  [31:0]         v0_1692;
  reg  [31:0]         v0_1693;
  reg  [31:0]         v0_1694;
  reg  [31:0]         v0_1695;
  reg  [31:0]         v0_1696;
  reg  [31:0]         v0_1697;
  reg  [31:0]         v0_1698;
  reg  [31:0]         v0_1699;
  reg  [31:0]         v0_1700;
  reg  [31:0]         v0_1701;
  reg  [31:0]         v0_1702;
  reg  [31:0]         v0_1703;
  reg  [31:0]         v0_1704;
  reg  [31:0]         v0_1705;
  reg  [31:0]         v0_1706;
  reg  [31:0]         v0_1707;
  reg  [31:0]         v0_1708;
  reg  [31:0]         v0_1709;
  reg  [31:0]         v0_1710;
  reg  [31:0]         v0_1711;
  reg  [31:0]         v0_1712;
  reg  [31:0]         v0_1713;
  reg  [31:0]         v0_1714;
  reg  [31:0]         v0_1715;
  reg  [31:0]         v0_1716;
  reg  [31:0]         v0_1717;
  reg  [31:0]         v0_1718;
  reg  [31:0]         v0_1719;
  reg  [31:0]         v0_1720;
  reg  [31:0]         v0_1721;
  reg  [31:0]         v0_1722;
  reg  [31:0]         v0_1723;
  reg  [31:0]         v0_1724;
  reg  [31:0]         v0_1725;
  reg  [31:0]         v0_1726;
  reg  [31:0]         v0_1727;
  reg  [31:0]         v0_1728;
  reg  [31:0]         v0_1729;
  reg  [31:0]         v0_1730;
  reg  [31:0]         v0_1731;
  reg  [31:0]         v0_1732;
  reg  [31:0]         v0_1733;
  reg  [31:0]         v0_1734;
  reg  [31:0]         v0_1735;
  reg  [31:0]         v0_1736;
  reg  [31:0]         v0_1737;
  reg  [31:0]         v0_1738;
  reg  [31:0]         v0_1739;
  reg  [31:0]         v0_1740;
  reg  [31:0]         v0_1741;
  reg  [31:0]         v0_1742;
  reg  [31:0]         v0_1743;
  reg  [31:0]         v0_1744;
  reg  [31:0]         v0_1745;
  reg  [31:0]         v0_1746;
  reg  [31:0]         v0_1747;
  reg  [31:0]         v0_1748;
  reg  [31:0]         v0_1749;
  reg  [31:0]         v0_1750;
  reg  [31:0]         v0_1751;
  reg  [31:0]         v0_1752;
  reg  [31:0]         v0_1753;
  reg  [31:0]         v0_1754;
  reg  [31:0]         v0_1755;
  reg  [31:0]         v0_1756;
  reg  [31:0]         v0_1757;
  reg  [31:0]         v0_1758;
  reg  [31:0]         v0_1759;
  reg  [31:0]         v0_1760;
  reg  [31:0]         v0_1761;
  reg  [31:0]         v0_1762;
  reg  [31:0]         v0_1763;
  reg  [31:0]         v0_1764;
  reg  [31:0]         v0_1765;
  reg  [31:0]         v0_1766;
  reg  [31:0]         v0_1767;
  reg  [31:0]         v0_1768;
  reg  [31:0]         v0_1769;
  reg  [31:0]         v0_1770;
  reg  [31:0]         v0_1771;
  reg  [31:0]         v0_1772;
  reg  [31:0]         v0_1773;
  reg  [31:0]         v0_1774;
  reg  [31:0]         v0_1775;
  reg  [31:0]         v0_1776;
  reg  [31:0]         v0_1777;
  reg  [31:0]         v0_1778;
  reg  [31:0]         v0_1779;
  reg  [31:0]         v0_1780;
  reg  [31:0]         v0_1781;
  reg  [31:0]         v0_1782;
  reg  [31:0]         v0_1783;
  reg  [31:0]         v0_1784;
  reg  [31:0]         v0_1785;
  reg  [31:0]         v0_1786;
  reg  [31:0]         v0_1787;
  reg  [31:0]         v0_1788;
  reg  [31:0]         v0_1789;
  reg  [31:0]         v0_1790;
  reg  [31:0]         v0_1791;
  reg  [31:0]         v0_1792;
  reg  [31:0]         v0_1793;
  reg  [31:0]         v0_1794;
  reg  [31:0]         v0_1795;
  reg  [31:0]         v0_1796;
  reg  [31:0]         v0_1797;
  reg  [31:0]         v0_1798;
  reg  [31:0]         v0_1799;
  reg  [31:0]         v0_1800;
  reg  [31:0]         v0_1801;
  reg  [31:0]         v0_1802;
  reg  [31:0]         v0_1803;
  reg  [31:0]         v0_1804;
  reg  [31:0]         v0_1805;
  reg  [31:0]         v0_1806;
  reg  [31:0]         v0_1807;
  reg  [31:0]         v0_1808;
  reg  [31:0]         v0_1809;
  reg  [31:0]         v0_1810;
  reg  [31:0]         v0_1811;
  reg  [31:0]         v0_1812;
  reg  [31:0]         v0_1813;
  reg  [31:0]         v0_1814;
  reg  [31:0]         v0_1815;
  reg  [31:0]         v0_1816;
  reg  [31:0]         v0_1817;
  reg  [31:0]         v0_1818;
  reg  [31:0]         v0_1819;
  reg  [31:0]         v0_1820;
  reg  [31:0]         v0_1821;
  reg  [31:0]         v0_1822;
  reg  [31:0]         v0_1823;
  reg  [31:0]         v0_1824;
  reg  [31:0]         v0_1825;
  reg  [31:0]         v0_1826;
  reg  [31:0]         v0_1827;
  reg  [31:0]         v0_1828;
  reg  [31:0]         v0_1829;
  reg  [31:0]         v0_1830;
  reg  [31:0]         v0_1831;
  reg  [31:0]         v0_1832;
  reg  [31:0]         v0_1833;
  reg  [31:0]         v0_1834;
  reg  [31:0]         v0_1835;
  reg  [31:0]         v0_1836;
  reg  [31:0]         v0_1837;
  reg  [31:0]         v0_1838;
  reg  [31:0]         v0_1839;
  reg  [31:0]         v0_1840;
  reg  [31:0]         v0_1841;
  reg  [31:0]         v0_1842;
  reg  [31:0]         v0_1843;
  reg  [31:0]         v0_1844;
  reg  [31:0]         v0_1845;
  reg  [31:0]         v0_1846;
  reg  [31:0]         v0_1847;
  reg  [31:0]         v0_1848;
  reg  [31:0]         v0_1849;
  reg  [31:0]         v0_1850;
  reg  [31:0]         v0_1851;
  reg  [31:0]         v0_1852;
  reg  [31:0]         v0_1853;
  reg  [31:0]         v0_1854;
  reg  [31:0]         v0_1855;
  reg  [31:0]         v0_1856;
  reg  [31:0]         v0_1857;
  reg  [31:0]         v0_1858;
  reg  [31:0]         v0_1859;
  reg  [31:0]         v0_1860;
  reg  [31:0]         v0_1861;
  reg  [31:0]         v0_1862;
  reg  [31:0]         v0_1863;
  reg  [31:0]         v0_1864;
  reg  [31:0]         v0_1865;
  reg  [31:0]         v0_1866;
  reg  [31:0]         v0_1867;
  reg  [31:0]         v0_1868;
  reg  [31:0]         v0_1869;
  reg  [31:0]         v0_1870;
  reg  [31:0]         v0_1871;
  reg  [31:0]         v0_1872;
  reg  [31:0]         v0_1873;
  reg  [31:0]         v0_1874;
  reg  [31:0]         v0_1875;
  reg  [31:0]         v0_1876;
  reg  [31:0]         v0_1877;
  reg  [31:0]         v0_1878;
  reg  [31:0]         v0_1879;
  reg  [31:0]         v0_1880;
  reg  [31:0]         v0_1881;
  reg  [31:0]         v0_1882;
  reg  [31:0]         v0_1883;
  reg  [31:0]         v0_1884;
  reg  [31:0]         v0_1885;
  reg  [31:0]         v0_1886;
  reg  [31:0]         v0_1887;
  reg  [31:0]         v0_1888;
  reg  [31:0]         v0_1889;
  reg  [31:0]         v0_1890;
  reg  [31:0]         v0_1891;
  reg  [31:0]         v0_1892;
  reg  [31:0]         v0_1893;
  reg  [31:0]         v0_1894;
  reg  [31:0]         v0_1895;
  reg  [31:0]         v0_1896;
  reg  [31:0]         v0_1897;
  reg  [31:0]         v0_1898;
  reg  [31:0]         v0_1899;
  reg  [31:0]         v0_1900;
  reg  [31:0]         v0_1901;
  reg  [31:0]         v0_1902;
  reg  [31:0]         v0_1903;
  reg  [31:0]         v0_1904;
  reg  [31:0]         v0_1905;
  reg  [31:0]         v0_1906;
  reg  [31:0]         v0_1907;
  reg  [31:0]         v0_1908;
  reg  [31:0]         v0_1909;
  reg  [31:0]         v0_1910;
  reg  [31:0]         v0_1911;
  reg  [31:0]         v0_1912;
  reg  [31:0]         v0_1913;
  reg  [31:0]         v0_1914;
  reg  [31:0]         v0_1915;
  reg  [31:0]         v0_1916;
  reg  [31:0]         v0_1917;
  reg  [31:0]         v0_1918;
  reg  [31:0]         v0_1919;
  reg  [31:0]         v0_1920;
  reg  [31:0]         v0_1921;
  reg  [31:0]         v0_1922;
  reg  [31:0]         v0_1923;
  reg  [31:0]         v0_1924;
  reg  [31:0]         v0_1925;
  reg  [31:0]         v0_1926;
  reg  [31:0]         v0_1927;
  reg  [31:0]         v0_1928;
  reg  [31:0]         v0_1929;
  reg  [31:0]         v0_1930;
  reg  [31:0]         v0_1931;
  reg  [31:0]         v0_1932;
  reg  [31:0]         v0_1933;
  reg  [31:0]         v0_1934;
  reg  [31:0]         v0_1935;
  reg  [31:0]         v0_1936;
  reg  [31:0]         v0_1937;
  reg  [31:0]         v0_1938;
  reg  [31:0]         v0_1939;
  reg  [31:0]         v0_1940;
  reg  [31:0]         v0_1941;
  reg  [31:0]         v0_1942;
  reg  [31:0]         v0_1943;
  reg  [31:0]         v0_1944;
  reg  [31:0]         v0_1945;
  reg  [31:0]         v0_1946;
  reg  [31:0]         v0_1947;
  reg  [31:0]         v0_1948;
  reg  [31:0]         v0_1949;
  reg  [31:0]         v0_1950;
  reg  [31:0]         v0_1951;
  reg  [31:0]         v0_1952;
  reg  [31:0]         v0_1953;
  reg  [31:0]         v0_1954;
  reg  [31:0]         v0_1955;
  reg  [31:0]         v0_1956;
  reg  [31:0]         v0_1957;
  reg  [31:0]         v0_1958;
  reg  [31:0]         v0_1959;
  reg  [31:0]         v0_1960;
  reg  [31:0]         v0_1961;
  reg  [31:0]         v0_1962;
  reg  [31:0]         v0_1963;
  reg  [31:0]         v0_1964;
  reg  [31:0]         v0_1965;
  reg  [31:0]         v0_1966;
  reg  [31:0]         v0_1967;
  reg  [31:0]         v0_1968;
  reg  [31:0]         v0_1969;
  reg  [31:0]         v0_1970;
  reg  [31:0]         v0_1971;
  reg  [31:0]         v0_1972;
  reg  [31:0]         v0_1973;
  reg  [31:0]         v0_1974;
  reg  [31:0]         v0_1975;
  reg  [31:0]         v0_1976;
  reg  [31:0]         v0_1977;
  reg  [31:0]         v0_1978;
  reg  [31:0]         v0_1979;
  reg  [31:0]         v0_1980;
  reg  [31:0]         v0_1981;
  reg  [31:0]         v0_1982;
  reg  [31:0]         v0_1983;
  reg  [31:0]         v0_1984;
  reg  [31:0]         v0_1985;
  reg  [31:0]         v0_1986;
  reg  [31:0]         v0_1987;
  reg  [31:0]         v0_1988;
  reg  [31:0]         v0_1989;
  reg  [31:0]         v0_1990;
  reg  [31:0]         v0_1991;
  reg  [31:0]         v0_1992;
  reg  [31:0]         v0_1993;
  reg  [31:0]         v0_1994;
  reg  [31:0]         v0_1995;
  reg  [31:0]         v0_1996;
  reg  [31:0]         v0_1997;
  reg  [31:0]         v0_1998;
  reg  [31:0]         v0_1999;
  reg  [31:0]         v0_2000;
  reg  [31:0]         v0_2001;
  reg  [31:0]         v0_2002;
  reg  [31:0]         v0_2003;
  reg  [31:0]         v0_2004;
  reg  [31:0]         v0_2005;
  reg  [31:0]         v0_2006;
  reg  [31:0]         v0_2007;
  reg  [31:0]         v0_2008;
  reg  [31:0]         v0_2009;
  reg  [31:0]         v0_2010;
  reg  [31:0]         v0_2011;
  reg  [31:0]         v0_2012;
  reg  [31:0]         v0_2013;
  reg  [31:0]         v0_2014;
  reg  [31:0]         v0_2015;
  reg  [31:0]         v0_2016;
  reg  [31:0]         v0_2017;
  reg  [31:0]         v0_2018;
  reg  [31:0]         v0_2019;
  reg  [31:0]         v0_2020;
  reg  [31:0]         v0_2021;
  reg  [31:0]         v0_2022;
  reg  [31:0]         v0_2023;
  reg  [31:0]         v0_2024;
  reg  [31:0]         v0_2025;
  reg  [31:0]         v0_2026;
  reg  [31:0]         v0_2027;
  reg  [31:0]         v0_2028;
  reg  [31:0]         v0_2029;
  reg  [31:0]         v0_2030;
  reg  [31:0]         v0_2031;
  reg  [31:0]         v0_2032;
  reg  [31:0]         v0_2033;
  reg  [31:0]         v0_2034;
  reg  [31:0]         v0_2035;
  reg  [31:0]         v0_2036;
  reg  [31:0]         v0_2037;
  reg  [31:0]         v0_2038;
  reg  [31:0]         v0_2039;
  reg  [31:0]         v0_2040;
  reg  [31:0]         v0_2041;
  reg  [31:0]         v0_2042;
  reg  [31:0]         v0_2043;
  reg  [31:0]         v0_2044;
  reg  [31:0]         v0_2045;
  reg  [31:0]         v0_2046;
  reg  [31:0]         v0_2047;
  wire [15:0]         maskExt_lo = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt = {maskExt_hi, maskExt_lo};
  wire [15:0]         maskExt_lo_1 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1 = {maskExt_hi_1, maskExt_lo_1};
  wire [15:0]         maskExt_lo_2 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_2 = {maskExt_hi_2, maskExt_lo_2};
  wire [15:0]         maskExt_lo_3 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_3 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_3 = {maskExt_hi_3, maskExt_lo_3};
  wire [15:0]         maskExt_lo_4 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_4 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_4 = {maskExt_hi_4, maskExt_lo_4};
  wire [15:0]         maskExt_lo_5 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_5 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_5 = {maskExt_hi_5, maskExt_lo_5};
  wire [15:0]         maskExt_lo_6 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_6 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_6 = {maskExt_hi_6, maskExt_lo_6};
  wire [15:0]         maskExt_lo_7 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_7 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_7 = {maskExt_hi_7, maskExt_lo_7};
  wire [15:0]         maskExt_lo_8 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_8 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_8 = {maskExt_hi_8, maskExt_lo_8};
  wire [15:0]         maskExt_lo_9 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_9 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_9 = {maskExt_hi_9, maskExt_lo_9};
  wire [15:0]         maskExt_lo_10 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_10 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_10 = {maskExt_hi_10, maskExt_lo_10};
  wire [15:0]         maskExt_lo_11 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_11 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_11 = {maskExt_hi_11, maskExt_lo_11};
  wire [15:0]         maskExt_lo_12 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_12 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_12 = {maskExt_hi_12, maskExt_lo_12};
  wire [15:0]         maskExt_lo_13 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_13 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_13 = {maskExt_hi_13, maskExt_lo_13};
  wire [15:0]         maskExt_lo_14 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_14 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_14 = {maskExt_hi_14, maskExt_lo_14};
  wire [15:0]         maskExt_lo_15 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_15 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_15 = {maskExt_hi_15, maskExt_lo_15};
  wire [15:0]         maskExt_lo_16 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_16 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_16 = {maskExt_hi_16, maskExt_lo_16};
  wire [15:0]         maskExt_lo_17 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_17 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_17 = {maskExt_hi_17, maskExt_lo_17};
  wire [15:0]         maskExt_lo_18 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_18 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_18 = {maskExt_hi_18, maskExt_lo_18};
  wire [15:0]         maskExt_lo_19 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_19 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_19 = {maskExt_hi_19, maskExt_lo_19};
  wire [15:0]         maskExt_lo_20 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_20 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_20 = {maskExt_hi_20, maskExt_lo_20};
  wire [15:0]         maskExt_lo_21 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_21 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_21 = {maskExt_hi_21, maskExt_lo_21};
  wire [15:0]         maskExt_lo_22 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_22 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_22 = {maskExt_hi_22, maskExt_lo_22};
  wire [15:0]         maskExt_lo_23 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_23 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_23 = {maskExt_hi_23, maskExt_lo_23};
  wire [15:0]         maskExt_lo_24 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_24 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_24 = {maskExt_hi_24, maskExt_lo_24};
  wire [15:0]         maskExt_lo_25 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_25 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_25 = {maskExt_hi_25, maskExt_lo_25};
  wire [15:0]         maskExt_lo_26 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_26 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_26 = {maskExt_hi_26, maskExt_lo_26};
  wire [15:0]         maskExt_lo_27 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_27 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_27 = {maskExt_hi_27, maskExt_lo_27};
  wire [15:0]         maskExt_lo_28 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_28 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_28 = {maskExt_hi_28, maskExt_lo_28};
  wire [15:0]         maskExt_lo_29 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_29 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_29 = {maskExt_hi_29, maskExt_lo_29};
  wire [15:0]         maskExt_lo_30 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_30 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_30 = {maskExt_hi_30, maskExt_lo_30};
  wire [15:0]         maskExt_lo_31 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_31 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_31 = {maskExt_hi_31, maskExt_lo_31};
  wire [15:0]         maskExt_lo_32 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_32 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_32 = {maskExt_hi_32, maskExt_lo_32};
  wire [15:0]         maskExt_lo_33 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_33 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_33 = {maskExt_hi_33, maskExt_lo_33};
  wire [15:0]         maskExt_lo_34 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_34 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_34 = {maskExt_hi_34, maskExt_lo_34};
  wire [15:0]         maskExt_lo_35 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_35 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_35 = {maskExt_hi_35, maskExt_lo_35};
  wire [15:0]         maskExt_lo_36 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_36 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_36 = {maskExt_hi_36, maskExt_lo_36};
  wire [15:0]         maskExt_lo_37 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_37 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_37 = {maskExt_hi_37, maskExt_lo_37};
  wire [15:0]         maskExt_lo_38 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_38 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_38 = {maskExt_hi_38, maskExt_lo_38};
  wire [15:0]         maskExt_lo_39 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_39 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_39 = {maskExt_hi_39, maskExt_lo_39};
  wire [15:0]         maskExt_lo_40 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_40 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_40 = {maskExt_hi_40, maskExt_lo_40};
  wire [15:0]         maskExt_lo_41 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_41 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_41 = {maskExt_hi_41, maskExt_lo_41};
  wire [15:0]         maskExt_lo_42 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_42 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_42 = {maskExt_hi_42, maskExt_lo_42};
  wire [15:0]         maskExt_lo_43 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_43 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_43 = {maskExt_hi_43, maskExt_lo_43};
  wire [15:0]         maskExt_lo_44 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_44 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_44 = {maskExt_hi_44, maskExt_lo_44};
  wire [15:0]         maskExt_lo_45 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_45 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_45 = {maskExt_hi_45, maskExt_lo_45};
  wire [15:0]         maskExt_lo_46 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_46 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_46 = {maskExt_hi_46, maskExt_lo_46};
  wire [15:0]         maskExt_lo_47 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_47 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_47 = {maskExt_hi_47, maskExt_lo_47};
  wire [15:0]         maskExt_lo_48 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_48 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_48 = {maskExt_hi_48, maskExt_lo_48};
  wire [15:0]         maskExt_lo_49 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_49 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_49 = {maskExt_hi_49, maskExt_lo_49};
  wire [15:0]         maskExt_lo_50 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_50 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_50 = {maskExt_hi_50, maskExt_lo_50};
  wire [15:0]         maskExt_lo_51 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_51 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_51 = {maskExt_hi_51, maskExt_lo_51};
  wire [15:0]         maskExt_lo_52 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_52 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_52 = {maskExt_hi_52, maskExt_lo_52};
  wire [15:0]         maskExt_lo_53 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_53 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_53 = {maskExt_hi_53, maskExt_lo_53};
  wire [15:0]         maskExt_lo_54 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_54 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_54 = {maskExt_hi_54, maskExt_lo_54};
  wire [15:0]         maskExt_lo_55 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_55 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_55 = {maskExt_hi_55, maskExt_lo_55};
  wire [15:0]         maskExt_lo_56 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_56 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_56 = {maskExt_hi_56, maskExt_lo_56};
  wire [15:0]         maskExt_lo_57 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_57 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_57 = {maskExt_hi_57, maskExt_lo_57};
  wire [15:0]         maskExt_lo_58 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_58 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_58 = {maskExt_hi_58, maskExt_lo_58};
  wire [15:0]         maskExt_lo_59 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_59 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_59 = {maskExt_hi_59, maskExt_lo_59};
  wire [15:0]         maskExt_lo_60 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_60 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_60 = {maskExt_hi_60, maskExt_lo_60};
  wire [15:0]         maskExt_lo_61 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_61 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_61 = {maskExt_hi_61, maskExt_lo_61};
  wire [15:0]         maskExt_lo_62 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_62 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_62 = {maskExt_hi_62, maskExt_lo_62};
  wire [15:0]         maskExt_lo_63 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_63 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_63 = {maskExt_hi_63, maskExt_lo_63};
  wire [15:0]         maskExt_lo_64 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_64 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_64 = {maskExt_hi_64, maskExt_lo_64};
  wire [15:0]         maskExt_lo_65 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_65 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_65 = {maskExt_hi_65, maskExt_lo_65};
  wire [15:0]         maskExt_lo_66 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_66 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_66 = {maskExt_hi_66, maskExt_lo_66};
  wire [15:0]         maskExt_lo_67 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_67 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_67 = {maskExt_hi_67, maskExt_lo_67};
  wire [15:0]         maskExt_lo_68 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_68 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_68 = {maskExt_hi_68, maskExt_lo_68};
  wire [15:0]         maskExt_lo_69 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_69 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_69 = {maskExt_hi_69, maskExt_lo_69};
  wire [15:0]         maskExt_lo_70 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_70 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_70 = {maskExt_hi_70, maskExt_lo_70};
  wire [15:0]         maskExt_lo_71 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_71 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_71 = {maskExt_hi_71, maskExt_lo_71};
  wire [15:0]         maskExt_lo_72 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_72 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_72 = {maskExt_hi_72, maskExt_lo_72};
  wire [15:0]         maskExt_lo_73 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_73 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_73 = {maskExt_hi_73, maskExt_lo_73};
  wire [15:0]         maskExt_lo_74 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_74 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_74 = {maskExt_hi_74, maskExt_lo_74};
  wire [15:0]         maskExt_lo_75 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_75 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_75 = {maskExt_hi_75, maskExt_lo_75};
  wire [15:0]         maskExt_lo_76 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_76 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_76 = {maskExt_hi_76, maskExt_lo_76};
  wire [15:0]         maskExt_lo_77 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_77 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_77 = {maskExt_hi_77, maskExt_lo_77};
  wire [15:0]         maskExt_lo_78 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_78 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_78 = {maskExt_hi_78, maskExt_lo_78};
  wire [15:0]         maskExt_lo_79 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_79 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_79 = {maskExt_hi_79, maskExt_lo_79};
  wire [15:0]         maskExt_lo_80 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_80 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_80 = {maskExt_hi_80, maskExt_lo_80};
  wire [15:0]         maskExt_lo_81 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_81 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_81 = {maskExt_hi_81, maskExt_lo_81};
  wire [15:0]         maskExt_lo_82 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_82 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_82 = {maskExt_hi_82, maskExt_lo_82};
  wire [15:0]         maskExt_lo_83 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_83 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_83 = {maskExt_hi_83, maskExt_lo_83};
  wire [15:0]         maskExt_lo_84 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_84 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_84 = {maskExt_hi_84, maskExt_lo_84};
  wire [15:0]         maskExt_lo_85 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_85 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_85 = {maskExt_hi_85, maskExt_lo_85};
  wire [15:0]         maskExt_lo_86 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_86 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_86 = {maskExt_hi_86, maskExt_lo_86};
  wire [15:0]         maskExt_lo_87 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_87 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_87 = {maskExt_hi_87, maskExt_lo_87};
  wire [15:0]         maskExt_lo_88 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_88 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_88 = {maskExt_hi_88, maskExt_lo_88};
  wire [15:0]         maskExt_lo_89 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_89 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_89 = {maskExt_hi_89, maskExt_lo_89};
  wire [15:0]         maskExt_lo_90 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_90 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_90 = {maskExt_hi_90, maskExt_lo_90};
  wire [15:0]         maskExt_lo_91 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_91 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_91 = {maskExt_hi_91, maskExt_lo_91};
  wire [15:0]         maskExt_lo_92 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_92 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_92 = {maskExt_hi_92, maskExt_lo_92};
  wire [15:0]         maskExt_lo_93 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_93 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_93 = {maskExt_hi_93, maskExt_lo_93};
  wire [15:0]         maskExt_lo_94 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_94 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_94 = {maskExt_hi_94, maskExt_lo_94};
  wire [15:0]         maskExt_lo_95 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_95 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_95 = {maskExt_hi_95, maskExt_lo_95};
  wire [15:0]         maskExt_lo_96 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_96 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_96 = {maskExt_hi_96, maskExt_lo_96};
  wire [15:0]         maskExt_lo_97 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_97 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_97 = {maskExt_hi_97, maskExt_lo_97};
  wire [15:0]         maskExt_lo_98 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_98 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_98 = {maskExt_hi_98, maskExt_lo_98};
  wire [15:0]         maskExt_lo_99 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_99 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_99 = {maskExt_hi_99, maskExt_lo_99};
  wire [15:0]         maskExt_lo_100 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_100 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_100 = {maskExt_hi_100, maskExt_lo_100};
  wire [15:0]         maskExt_lo_101 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_101 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_101 = {maskExt_hi_101, maskExt_lo_101};
  wire [15:0]         maskExt_lo_102 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_102 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_102 = {maskExt_hi_102, maskExt_lo_102};
  wire [15:0]         maskExt_lo_103 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_103 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_103 = {maskExt_hi_103, maskExt_lo_103};
  wire [15:0]         maskExt_lo_104 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_104 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_104 = {maskExt_hi_104, maskExt_lo_104};
  wire [15:0]         maskExt_lo_105 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_105 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_105 = {maskExt_hi_105, maskExt_lo_105};
  wire [15:0]         maskExt_lo_106 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_106 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_106 = {maskExt_hi_106, maskExt_lo_106};
  wire [15:0]         maskExt_lo_107 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_107 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_107 = {maskExt_hi_107, maskExt_lo_107};
  wire [15:0]         maskExt_lo_108 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_108 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_108 = {maskExt_hi_108, maskExt_lo_108};
  wire [15:0]         maskExt_lo_109 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_109 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_109 = {maskExt_hi_109, maskExt_lo_109};
  wire [15:0]         maskExt_lo_110 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_110 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_110 = {maskExt_hi_110, maskExt_lo_110};
  wire [15:0]         maskExt_lo_111 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_111 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_111 = {maskExt_hi_111, maskExt_lo_111};
  wire [15:0]         maskExt_lo_112 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_112 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_112 = {maskExt_hi_112, maskExt_lo_112};
  wire [15:0]         maskExt_lo_113 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_113 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_113 = {maskExt_hi_113, maskExt_lo_113};
  wire [15:0]         maskExt_lo_114 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_114 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_114 = {maskExt_hi_114, maskExt_lo_114};
  wire [15:0]         maskExt_lo_115 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_115 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_115 = {maskExt_hi_115, maskExt_lo_115};
  wire [15:0]         maskExt_lo_116 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_116 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_116 = {maskExt_hi_116, maskExt_lo_116};
  wire [15:0]         maskExt_lo_117 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_117 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_117 = {maskExt_hi_117, maskExt_lo_117};
  wire [15:0]         maskExt_lo_118 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_118 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_118 = {maskExt_hi_118, maskExt_lo_118};
  wire [15:0]         maskExt_lo_119 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_119 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_119 = {maskExt_hi_119, maskExt_lo_119};
  wire [15:0]         maskExt_lo_120 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_120 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_120 = {maskExt_hi_120, maskExt_lo_120};
  wire [15:0]         maskExt_lo_121 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_121 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_121 = {maskExt_hi_121, maskExt_lo_121};
  wire [15:0]         maskExt_lo_122 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_122 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_122 = {maskExt_hi_122, maskExt_lo_122};
  wire [15:0]         maskExt_lo_123 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_123 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_123 = {maskExt_hi_123, maskExt_lo_123};
  wire [15:0]         maskExt_lo_124 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_124 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_124 = {maskExt_hi_124, maskExt_lo_124};
  wire [15:0]         maskExt_lo_125 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_125 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_125 = {maskExt_hi_125, maskExt_lo_125};
  wire [15:0]         maskExt_lo_126 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_126 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_126 = {maskExt_hi_126, maskExt_lo_126};
  wire [15:0]         maskExt_lo_127 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_127 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_127 = {maskExt_hi_127, maskExt_lo_127};
  wire [15:0]         maskExt_lo_128 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_128 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_128 = {maskExt_hi_128, maskExt_lo_128};
  wire [15:0]         maskExt_lo_129 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_129 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_129 = {maskExt_hi_129, maskExt_lo_129};
  wire [15:0]         maskExt_lo_130 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_130 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_130 = {maskExt_hi_130, maskExt_lo_130};
  wire [15:0]         maskExt_lo_131 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_131 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_131 = {maskExt_hi_131, maskExt_lo_131};
  wire [15:0]         maskExt_lo_132 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_132 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_132 = {maskExt_hi_132, maskExt_lo_132};
  wire [15:0]         maskExt_lo_133 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_133 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_133 = {maskExt_hi_133, maskExt_lo_133};
  wire [15:0]         maskExt_lo_134 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_134 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_134 = {maskExt_hi_134, maskExt_lo_134};
  wire [15:0]         maskExt_lo_135 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_135 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_135 = {maskExt_hi_135, maskExt_lo_135};
  wire [15:0]         maskExt_lo_136 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_136 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_136 = {maskExt_hi_136, maskExt_lo_136};
  wire [15:0]         maskExt_lo_137 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_137 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_137 = {maskExt_hi_137, maskExt_lo_137};
  wire [15:0]         maskExt_lo_138 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_138 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_138 = {maskExt_hi_138, maskExt_lo_138};
  wire [15:0]         maskExt_lo_139 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_139 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_139 = {maskExt_hi_139, maskExt_lo_139};
  wire [15:0]         maskExt_lo_140 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_140 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_140 = {maskExt_hi_140, maskExt_lo_140};
  wire [15:0]         maskExt_lo_141 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_141 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_141 = {maskExt_hi_141, maskExt_lo_141};
  wire [15:0]         maskExt_lo_142 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_142 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_142 = {maskExt_hi_142, maskExt_lo_142};
  wire [15:0]         maskExt_lo_143 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_143 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_143 = {maskExt_hi_143, maskExt_lo_143};
  wire [15:0]         maskExt_lo_144 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_144 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_144 = {maskExt_hi_144, maskExt_lo_144};
  wire [15:0]         maskExt_lo_145 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_145 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_145 = {maskExt_hi_145, maskExt_lo_145};
  wire [15:0]         maskExt_lo_146 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_146 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_146 = {maskExt_hi_146, maskExt_lo_146};
  wire [15:0]         maskExt_lo_147 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_147 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_147 = {maskExt_hi_147, maskExt_lo_147};
  wire [15:0]         maskExt_lo_148 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_148 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_148 = {maskExt_hi_148, maskExt_lo_148};
  wire [15:0]         maskExt_lo_149 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_149 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_149 = {maskExt_hi_149, maskExt_lo_149};
  wire [15:0]         maskExt_lo_150 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_150 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_150 = {maskExt_hi_150, maskExt_lo_150};
  wire [15:0]         maskExt_lo_151 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_151 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_151 = {maskExt_hi_151, maskExt_lo_151};
  wire [15:0]         maskExt_lo_152 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_152 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_152 = {maskExt_hi_152, maskExt_lo_152};
  wire [15:0]         maskExt_lo_153 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_153 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_153 = {maskExt_hi_153, maskExt_lo_153};
  wire [15:0]         maskExt_lo_154 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_154 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_154 = {maskExt_hi_154, maskExt_lo_154};
  wire [15:0]         maskExt_lo_155 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_155 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_155 = {maskExt_hi_155, maskExt_lo_155};
  wire [15:0]         maskExt_lo_156 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_156 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_156 = {maskExt_hi_156, maskExt_lo_156};
  wire [15:0]         maskExt_lo_157 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_157 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_157 = {maskExt_hi_157, maskExt_lo_157};
  wire [15:0]         maskExt_lo_158 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_158 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_158 = {maskExt_hi_158, maskExt_lo_158};
  wire [15:0]         maskExt_lo_159 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_159 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_159 = {maskExt_hi_159, maskExt_lo_159};
  wire [15:0]         maskExt_lo_160 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_160 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_160 = {maskExt_hi_160, maskExt_lo_160};
  wire [15:0]         maskExt_lo_161 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_161 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_161 = {maskExt_hi_161, maskExt_lo_161};
  wire [15:0]         maskExt_lo_162 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_162 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_162 = {maskExt_hi_162, maskExt_lo_162};
  wire [15:0]         maskExt_lo_163 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_163 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_163 = {maskExt_hi_163, maskExt_lo_163};
  wire [15:0]         maskExt_lo_164 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_164 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_164 = {maskExt_hi_164, maskExt_lo_164};
  wire [15:0]         maskExt_lo_165 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_165 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_165 = {maskExt_hi_165, maskExt_lo_165};
  wire [15:0]         maskExt_lo_166 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_166 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_166 = {maskExt_hi_166, maskExt_lo_166};
  wire [15:0]         maskExt_lo_167 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_167 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_167 = {maskExt_hi_167, maskExt_lo_167};
  wire [15:0]         maskExt_lo_168 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_168 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_168 = {maskExt_hi_168, maskExt_lo_168};
  wire [15:0]         maskExt_lo_169 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_169 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_169 = {maskExt_hi_169, maskExt_lo_169};
  wire [15:0]         maskExt_lo_170 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_170 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_170 = {maskExt_hi_170, maskExt_lo_170};
  wire [15:0]         maskExt_lo_171 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_171 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_171 = {maskExt_hi_171, maskExt_lo_171};
  wire [15:0]         maskExt_lo_172 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_172 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_172 = {maskExt_hi_172, maskExt_lo_172};
  wire [15:0]         maskExt_lo_173 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_173 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_173 = {maskExt_hi_173, maskExt_lo_173};
  wire [15:0]         maskExt_lo_174 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_174 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_174 = {maskExt_hi_174, maskExt_lo_174};
  wire [15:0]         maskExt_lo_175 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_175 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_175 = {maskExt_hi_175, maskExt_lo_175};
  wire [15:0]         maskExt_lo_176 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_176 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_176 = {maskExt_hi_176, maskExt_lo_176};
  wire [15:0]         maskExt_lo_177 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_177 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_177 = {maskExt_hi_177, maskExt_lo_177};
  wire [15:0]         maskExt_lo_178 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_178 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_178 = {maskExt_hi_178, maskExt_lo_178};
  wire [15:0]         maskExt_lo_179 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_179 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_179 = {maskExt_hi_179, maskExt_lo_179};
  wire [15:0]         maskExt_lo_180 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_180 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_180 = {maskExt_hi_180, maskExt_lo_180};
  wire [15:0]         maskExt_lo_181 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_181 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_181 = {maskExt_hi_181, maskExt_lo_181};
  wire [15:0]         maskExt_lo_182 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_182 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_182 = {maskExt_hi_182, maskExt_lo_182};
  wire [15:0]         maskExt_lo_183 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_183 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_183 = {maskExt_hi_183, maskExt_lo_183};
  wire [15:0]         maskExt_lo_184 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_184 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_184 = {maskExt_hi_184, maskExt_lo_184};
  wire [15:0]         maskExt_lo_185 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_185 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_185 = {maskExt_hi_185, maskExt_lo_185};
  wire [15:0]         maskExt_lo_186 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_186 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_186 = {maskExt_hi_186, maskExt_lo_186};
  wire [15:0]         maskExt_lo_187 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_187 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_187 = {maskExt_hi_187, maskExt_lo_187};
  wire [15:0]         maskExt_lo_188 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_188 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_188 = {maskExt_hi_188, maskExt_lo_188};
  wire [15:0]         maskExt_lo_189 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_189 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_189 = {maskExt_hi_189, maskExt_lo_189};
  wire [15:0]         maskExt_lo_190 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_190 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_190 = {maskExt_hi_190, maskExt_lo_190};
  wire [15:0]         maskExt_lo_191 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_191 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_191 = {maskExt_hi_191, maskExt_lo_191};
  wire [15:0]         maskExt_lo_192 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_192 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_192 = {maskExt_hi_192, maskExt_lo_192};
  wire [15:0]         maskExt_lo_193 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_193 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_193 = {maskExt_hi_193, maskExt_lo_193};
  wire [15:0]         maskExt_lo_194 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_194 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_194 = {maskExt_hi_194, maskExt_lo_194};
  wire [15:0]         maskExt_lo_195 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_195 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_195 = {maskExt_hi_195, maskExt_lo_195};
  wire [15:0]         maskExt_lo_196 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_196 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_196 = {maskExt_hi_196, maskExt_lo_196};
  wire [15:0]         maskExt_lo_197 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_197 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_197 = {maskExt_hi_197, maskExt_lo_197};
  wire [15:0]         maskExt_lo_198 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_198 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_198 = {maskExt_hi_198, maskExt_lo_198};
  wire [15:0]         maskExt_lo_199 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_199 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_199 = {maskExt_hi_199, maskExt_lo_199};
  wire [15:0]         maskExt_lo_200 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_200 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_200 = {maskExt_hi_200, maskExt_lo_200};
  wire [15:0]         maskExt_lo_201 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_201 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_201 = {maskExt_hi_201, maskExt_lo_201};
  wire [15:0]         maskExt_lo_202 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_202 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_202 = {maskExt_hi_202, maskExt_lo_202};
  wire [15:0]         maskExt_lo_203 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_203 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_203 = {maskExt_hi_203, maskExt_lo_203};
  wire [15:0]         maskExt_lo_204 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_204 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_204 = {maskExt_hi_204, maskExt_lo_204};
  wire [15:0]         maskExt_lo_205 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_205 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_205 = {maskExt_hi_205, maskExt_lo_205};
  wire [15:0]         maskExt_lo_206 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_206 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_206 = {maskExt_hi_206, maskExt_lo_206};
  wire [15:0]         maskExt_lo_207 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_207 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_207 = {maskExt_hi_207, maskExt_lo_207};
  wire [15:0]         maskExt_lo_208 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_208 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_208 = {maskExt_hi_208, maskExt_lo_208};
  wire [15:0]         maskExt_lo_209 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_209 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_209 = {maskExt_hi_209, maskExt_lo_209};
  wire [15:0]         maskExt_lo_210 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_210 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_210 = {maskExt_hi_210, maskExt_lo_210};
  wire [15:0]         maskExt_lo_211 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_211 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_211 = {maskExt_hi_211, maskExt_lo_211};
  wire [15:0]         maskExt_lo_212 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_212 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_212 = {maskExt_hi_212, maskExt_lo_212};
  wire [15:0]         maskExt_lo_213 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_213 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_213 = {maskExt_hi_213, maskExt_lo_213};
  wire [15:0]         maskExt_lo_214 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_214 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_214 = {maskExt_hi_214, maskExt_lo_214};
  wire [15:0]         maskExt_lo_215 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_215 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_215 = {maskExt_hi_215, maskExt_lo_215};
  wire [15:0]         maskExt_lo_216 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_216 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_216 = {maskExt_hi_216, maskExt_lo_216};
  wire [15:0]         maskExt_lo_217 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_217 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_217 = {maskExt_hi_217, maskExt_lo_217};
  wire [15:0]         maskExt_lo_218 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_218 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_218 = {maskExt_hi_218, maskExt_lo_218};
  wire [15:0]         maskExt_lo_219 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_219 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_219 = {maskExt_hi_219, maskExt_lo_219};
  wire [15:0]         maskExt_lo_220 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_220 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_220 = {maskExt_hi_220, maskExt_lo_220};
  wire [15:0]         maskExt_lo_221 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_221 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_221 = {maskExt_hi_221, maskExt_lo_221};
  wire [15:0]         maskExt_lo_222 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_222 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_222 = {maskExt_hi_222, maskExt_lo_222};
  wire [15:0]         maskExt_lo_223 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_223 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_223 = {maskExt_hi_223, maskExt_lo_223};
  wire [15:0]         maskExt_lo_224 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_224 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_224 = {maskExt_hi_224, maskExt_lo_224};
  wire [15:0]         maskExt_lo_225 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_225 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_225 = {maskExt_hi_225, maskExt_lo_225};
  wire [15:0]         maskExt_lo_226 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_226 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_226 = {maskExt_hi_226, maskExt_lo_226};
  wire [15:0]         maskExt_lo_227 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_227 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_227 = {maskExt_hi_227, maskExt_lo_227};
  wire [15:0]         maskExt_lo_228 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_228 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_228 = {maskExt_hi_228, maskExt_lo_228};
  wire [15:0]         maskExt_lo_229 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_229 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_229 = {maskExt_hi_229, maskExt_lo_229};
  wire [15:0]         maskExt_lo_230 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_230 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_230 = {maskExt_hi_230, maskExt_lo_230};
  wire [15:0]         maskExt_lo_231 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_231 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_231 = {maskExt_hi_231, maskExt_lo_231};
  wire [15:0]         maskExt_lo_232 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_232 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_232 = {maskExt_hi_232, maskExt_lo_232};
  wire [15:0]         maskExt_lo_233 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_233 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_233 = {maskExt_hi_233, maskExt_lo_233};
  wire [15:0]         maskExt_lo_234 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_234 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_234 = {maskExt_hi_234, maskExt_lo_234};
  wire [15:0]         maskExt_lo_235 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_235 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_235 = {maskExt_hi_235, maskExt_lo_235};
  wire [15:0]         maskExt_lo_236 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_236 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_236 = {maskExt_hi_236, maskExt_lo_236};
  wire [15:0]         maskExt_lo_237 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_237 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_237 = {maskExt_hi_237, maskExt_lo_237};
  wire [15:0]         maskExt_lo_238 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_238 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_238 = {maskExt_hi_238, maskExt_lo_238};
  wire [15:0]         maskExt_lo_239 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_239 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_239 = {maskExt_hi_239, maskExt_lo_239};
  wire [15:0]         maskExt_lo_240 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_240 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_240 = {maskExt_hi_240, maskExt_lo_240};
  wire [15:0]         maskExt_lo_241 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_241 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_241 = {maskExt_hi_241, maskExt_lo_241};
  wire [15:0]         maskExt_lo_242 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_242 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_242 = {maskExt_hi_242, maskExt_lo_242};
  wire [15:0]         maskExt_lo_243 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_243 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_243 = {maskExt_hi_243, maskExt_lo_243};
  wire [15:0]         maskExt_lo_244 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_244 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_244 = {maskExt_hi_244, maskExt_lo_244};
  wire [15:0]         maskExt_lo_245 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_245 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_245 = {maskExt_hi_245, maskExt_lo_245};
  wire [15:0]         maskExt_lo_246 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_246 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_246 = {maskExt_hi_246, maskExt_lo_246};
  wire [15:0]         maskExt_lo_247 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_247 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_247 = {maskExt_hi_247, maskExt_lo_247};
  wire [15:0]         maskExt_lo_248 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_248 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_248 = {maskExt_hi_248, maskExt_lo_248};
  wire [15:0]         maskExt_lo_249 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_249 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_249 = {maskExt_hi_249, maskExt_lo_249};
  wire [15:0]         maskExt_lo_250 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_250 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_250 = {maskExt_hi_250, maskExt_lo_250};
  wire [15:0]         maskExt_lo_251 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_251 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_251 = {maskExt_hi_251, maskExt_lo_251};
  wire [15:0]         maskExt_lo_252 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_252 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_252 = {maskExt_hi_252, maskExt_lo_252};
  wire [15:0]         maskExt_lo_253 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_253 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_253 = {maskExt_hi_253, maskExt_lo_253};
  wire [15:0]         maskExt_lo_254 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_254 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_254 = {maskExt_hi_254, maskExt_lo_254};
  wire [15:0]         maskExt_lo_255 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_255 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_255 = {maskExt_hi_255, maskExt_lo_255};
  wire [15:0]         maskExt_lo_256 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_256 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_256 = {maskExt_hi_256, maskExt_lo_256};
  wire [15:0]         maskExt_lo_257 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_257 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_257 = {maskExt_hi_257, maskExt_lo_257};
  wire [15:0]         maskExt_lo_258 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_258 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_258 = {maskExt_hi_258, maskExt_lo_258};
  wire [15:0]         maskExt_lo_259 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_259 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_259 = {maskExt_hi_259, maskExt_lo_259};
  wire [15:0]         maskExt_lo_260 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_260 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_260 = {maskExt_hi_260, maskExt_lo_260};
  wire [15:0]         maskExt_lo_261 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_261 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_261 = {maskExt_hi_261, maskExt_lo_261};
  wire [15:0]         maskExt_lo_262 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_262 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_262 = {maskExt_hi_262, maskExt_lo_262};
  wire [15:0]         maskExt_lo_263 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_263 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_263 = {maskExt_hi_263, maskExt_lo_263};
  wire [15:0]         maskExt_lo_264 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_264 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_264 = {maskExt_hi_264, maskExt_lo_264};
  wire [15:0]         maskExt_lo_265 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_265 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_265 = {maskExt_hi_265, maskExt_lo_265};
  wire [15:0]         maskExt_lo_266 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_266 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_266 = {maskExt_hi_266, maskExt_lo_266};
  wire [15:0]         maskExt_lo_267 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_267 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_267 = {maskExt_hi_267, maskExt_lo_267};
  wire [15:0]         maskExt_lo_268 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_268 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_268 = {maskExt_hi_268, maskExt_lo_268};
  wire [15:0]         maskExt_lo_269 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_269 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_269 = {maskExt_hi_269, maskExt_lo_269};
  wire [15:0]         maskExt_lo_270 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_270 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_270 = {maskExt_hi_270, maskExt_lo_270};
  wire [15:0]         maskExt_lo_271 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_271 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_271 = {maskExt_hi_271, maskExt_lo_271};
  wire [15:0]         maskExt_lo_272 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_272 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_272 = {maskExt_hi_272, maskExt_lo_272};
  wire [15:0]         maskExt_lo_273 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_273 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_273 = {maskExt_hi_273, maskExt_lo_273};
  wire [15:0]         maskExt_lo_274 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_274 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_274 = {maskExt_hi_274, maskExt_lo_274};
  wire [15:0]         maskExt_lo_275 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_275 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_275 = {maskExt_hi_275, maskExt_lo_275};
  wire [15:0]         maskExt_lo_276 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_276 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_276 = {maskExt_hi_276, maskExt_lo_276};
  wire [15:0]         maskExt_lo_277 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_277 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_277 = {maskExt_hi_277, maskExt_lo_277};
  wire [15:0]         maskExt_lo_278 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_278 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_278 = {maskExt_hi_278, maskExt_lo_278};
  wire [15:0]         maskExt_lo_279 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_279 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_279 = {maskExt_hi_279, maskExt_lo_279};
  wire [15:0]         maskExt_lo_280 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_280 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_280 = {maskExt_hi_280, maskExt_lo_280};
  wire [15:0]         maskExt_lo_281 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_281 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_281 = {maskExt_hi_281, maskExt_lo_281};
  wire [15:0]         maskExt_lo_282 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_282 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_282 = {maskExt_hi_282, maskExt_lo_282};
  wire [15:0]         maskExt_lo_283 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_283 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_283 = {maskExt_hi_283, maskExt_lo_283};
  wire [15:0]         maskExt_lo_284 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_284 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_284 = {maskExt_hi_284, maskExt_lo_284};
  wire [15:0]         maskExt_lo_285 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_285 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_285 = {maskExt_hi_285, maskExt_lo_285};
  wire [15:0]         maskExt_lo_286 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_286 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_286 = {maskExt_hi_286, maskExt_lo_286};
  wire [15:0]         maskExt_lo_287 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_287 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_287 = {maskExt_hi_287, maskExt_lo_287};
  wire [15:0]         maskExt_lo_288 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_288 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_288 = {maskExt_hi_288, maskExt_lo_288};
  wire [15:0]         maskExt_lo_289 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_289 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_289 = {maskExt_hi_289, maskExt_lo_289};
  wire [15:0]         maskExt_lo_290 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_290 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_290 = {maskExt_hi_290, maskExt_lo_290};
  wire [15:0]         maskExt_lo_291 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_291 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_291 = {maskExt_hi_291, maskExt_lo_291};
  wire [15:0]         maskExt_lo_292 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_292 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_292 = {maskExt_hi_292, maskExt_lo_292};
  wire [15:0]         maskExt_lo_293 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_293 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_293 = {maskExt_hi_293, maskExt_lo_293};
  wire [15:0]         maskExt_lo_294 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_294 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_294 = {maskExt_hi_294, maskExt_lo_294};
  wire [15:0]         maskExt_lo_295 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_295 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_295 = {maskExt_hi_295, maskExt_lo_295};
  wire [15:0]         maskExt_lo_296 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_296 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_296 = {maskExt_hi_296, maskExt_lo_296};
  wire [15:0]         maskExt_lo_297 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_297 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_297 = {maskExt_hi_297, maskExt_lo_297};
  wire [15:0]         maskExt_lo_298 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_298 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_298 = {maskExt_hi_298, maskExt_lo_298};
  wire [15:0]         maskExt_lo_299 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_299 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_299 = {maskExt_hi_299, maskExt_lo_299};
  wire [15:0]         maskExt_lo_300 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_300 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_300 = {maskExt_hi_300, maskExt_lo_300};
  wire [15:0]         maskExt_lo_301 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_301 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_301 = {maskExt_hi_301, maskExt_lo_301};
  wire [15:0]         maskExt_lo_302 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_302 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_302 = {maskExt_hi_302, maskExt_lo_302};
  wire [15:0]         maskExt_lo_303 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_303 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_303 = {maskExt_hi_303, maskExt_lo_303};
  wire [15:0]         maskExt_lo_304 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_304 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_304 = {maskExt_hi_304, maskExt_lo_304};
  wire [15:0]         maskExt_lo_305 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_305 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_305 = {maskExt_hi_305, maskExt_lo_305};
  wire [15:0]         maskExt_lo_306 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_306 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_306 = {maskExt_hi_306, maskExt_lo_306};
  wire [15:0]         maskExt_lo_307 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_307 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_307 = {maskExt_hi_307, maskExt_lo_307};
  wire [15:0]         maskExt_lo_308 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_308 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_308 = {maskExt_hi_308, maskExt_lo_308};
  wire [15:0]         maskExt_lo_309 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_309 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_309 = {maskExt_hi_309, maskExt_lo_309};
  wire [15:0]         maskExt_lo_310 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_310 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_310 = {maskExt_hi_310, maskExt_lo_310};
  wire [15:0]         maskExt_lo_311 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_311 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_311 = {maskExt_hi_311, maskExt_lo_311};
  wire [15:0]         maskExt_lo_312 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_312 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_312 = {maskExt_hi_312, maskExt_lo_312};
  wire [15:0]         maskExt_lo_313 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_313 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_313 = {maskExt_hi_313, maskExt_lo_313};
  wire [15:0]         maskExt_lo_314 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_314 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_314 = {maskExt_hi_314, maskExt_lo_314};
  wire [15:0]         maskExt_lo_315 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_315 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_315 = {maskExt_hi_315, maskExt_lo_315};
  wire [15:0]         maskExt_lo_316 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_316 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_316 = {maskExt_hi_316, maskExt_lo_316};
  wire [15:0]         maskExt_lo_317 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_317 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_317 = {maskExt_hi_317, maskExt_lo_317};
  wire [15:0]         maskExt_lo_318 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_318 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_318 = {maskExt_hi_318, maskExt_lo_318};
  wire [15:0]         maskExt_lo_319 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_319 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_319 = {maskExt_hi_319, maskExt_lo_319};
  wire [15:0]         maskExt_lo_320 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_320 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_320 = {maskExt_hi_320, maskExt_lo_320};
  wire [15:0]         maskExt_lo_321 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_321 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_321 = {maskExt_hi_321, maskExt_lo_321};
  wire [15:0]         maskExt_lo_322 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_322 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_322 = {maskExt_hi_322, maskExt_lo_322};
  wire [15:0]         maskExt_lo_323 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_323 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_323 = {maskExt_hi_323, maskExt_lo_323};
  wire [15:0]         maskExt_lo_324 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_324 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_324 = {maskExt_hi_324, maskExt_lo_324};
  wire [15:0]         maskExt_lo_325 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_325 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_325 = {maskExt_hi_325, maskExt_lo_325};
  wire [15:0]         maskExt_lo_326 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_326 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_326 = {maskExt_hi_326, maskExt_lo_326};
  wire [15:0]         maskExt_lo_327 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_327 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_327 = {maskExt_hi_327, maskExt_lo_327};
  wire [15:0]         maskExt_lo_328 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_328 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_328 = {maskExt_hi_328, maskExt_lo_328};
  wire [15:0]         maskExt_lo_329 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_329 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_329 = {maskExt_hi_329, maskExt_lo_329};
  wire [15:0]         maskExt_lo_330 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_330 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_330 = {maskExt_hi_330, maskExt_lo_330};
  wire [15:0]         maskExt_lo_331 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_331 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_331 = {maskExt_hi_331, maskExt_lo_331};
  wire [15:0]         maskExt_lo_332 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_332 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_332 = {maskExt_hi_332, maskExt_lo_332};
  wire [15:0]         maskExt_lo_333 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_333 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_333 = {maskExt_hi_333, maskExt_lo_333};
  wire [15:0]         maskExt_lo_334 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_334 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_334 = {maskExt_hi_334, maskExt_lo_334};
  wire [15:0]         maskExt_lo_335 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_335 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_335 = {maskExt_hi_335, maskExt_lo_335};
  wire [15:0]         maskExt_lo_336 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_336 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_336 = {maskExt_hi_336, maskExt_lo_336};
  wire [15:0]         maskExt_lo_337 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_337 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_337 = {maskExt_hi_337, maskExt_lo_337};
  wire [15:0]         maskExt_lo_338 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_338 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_338 = {maskExt_hi_338, maskExt_lo_338};
  wire [15:0]         maskExt_lo_339 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_339 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_339 = {maskExt_hi_339, maskExt_lo_339};
  wire [15:0]         maskExt_lo_340 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_340 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_340 = {maskExt_hi_340, maskExt_lo_340};
  wire [15:0]         maskExt_lo_341 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_341 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_341 = {maskExt_hi_341, maskExt_lo_341};
  wire [15:0]         maskExt_lo_342 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_342 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_342 = {maskExt_hi_342, maskExt_lo_342};
  wire [15:0]         maskExt_lo_343 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_343 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_343 = {maskExt_hi_343, maskExt_lo_343};
  wire [15:0]         maskExt_lo_344 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_344 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_344 = {maskExt_hi_344, maskExt_lo_344};
  wire [15:0]         maskExt_lo_345 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_345 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_345 = {maskExt_hi_345, maskExt_lo_345};
  wire [15:0]         maskExt_lo_346 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_346 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_346 = {maskExt_hi_346, maskExt_lo_346};
  wire [15:0]         maskExt_lo_347 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_347 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_347 = {maskExt_hi_347, maskExt_lo_347};
  wire [15:0]         maskExt_lo_348 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_348 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_348 = {maskExt_hi_348, maskExt_lo_348};
  wire [15:0]         maskExt_lo_349 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_349 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_349 = {maskExt_hi_349, maskExt_lo_349};
  wire [15:0]         maskExt_lo_350 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_350 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_350 = {maskExt_hi_350, maskExt_lo_350};
  wire [15:0]         maskExt_lo_351 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_351 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_351 = {maskExt_hi_351, maskExt_lo_351};
  wire [15:0]         maskExt_lo_352 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_352 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_352 = {maskExt_hi_352, maskExt_lo_352};
  wire [15:0]         maskExt_lo_353 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_353 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_353 = {maskExt_hi_353, maskExt_lo_353};
  wire [15:0]         maskExt_lo_354 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_354 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_354 = {maskExt_hi_354, maskExt_lo_354};
  wire [15:0]         maskExt_lo_355 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_355 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_355 = {maskExt_hi_355, maskExt_lo_355};
  wire [15:0]         maskExt_lo_356 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_356 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_356 = {maskExt_hi_356, maskExt_lo_356};
  wire [15:0]         maskExt_lo_357 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_357 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_357 = {maskExt_hi_357, maskExt_lo_357};
  wire [15:0]         maskExt_lo_358 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_358 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_358 = {maskExt_hi_358, maskExt_lo_358};
  wire [15:0]         maskExt_lo_359 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_359 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_359 = {maskExt_hi_359, maskExt_lo_359};
  wire [15:0]         maskExt_lo_360 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_360 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_360 = {maskExt_hi_360, maskExt_lo_360};
  wire [15:0]         maskExt_lo_361 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_361 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_361 = {maskExt_hi_361, maskExt_lo_361};
  wire [15:0]         maskExt_lo_362 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_362 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_362 = {maskExt_hi_362, maskExt_lo_362};
  wire [15:0]         maskExt_lo_363 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_363 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_363 = {maskExt_hi_363, maskExt_lo_363};
  wire [15:0]         maskExt_lo_364 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_364 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_364 = {maskExt_hi_364, maskExt_lo_364};
  wire [15:0]         maskExt_lo_365 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_365 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_365 = {maskExt_hi_365, maskExt_lo_365};
  wire [15:0]         maskExt_lo_366 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_366 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_366 = {maskExt_hi_366, maskExt_lo_366};
  wire [15:0]         maskExt_lo_367 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_367 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_367 = {maskExt_hi_367, maskExt_lo_367};
  wire [15:0]         maskExt_lo_368 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_368 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_368 = {maskExt_hi_368, maskExt_lo_368};
  wire [15:0]         maskExt_lo_369 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_369 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_369 = {maskExt_hi_369, maskExt_lo_369};
  wire [15:0]         maskExt_lo_370 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_370 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_370 = {maskExt_hi_370, maskExt_lo_370};
  wire [15:0]         maskExt_lo_371 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_371 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_371 = {maskExt_hi_371, maskExt_lo_371};
  wire [15:0]         maskExt_lo_372 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_372 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_372 = {maskExt_hi_372, maskExt_lo_372};
  wire [15:0]         maskExt_lo_373 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_373 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_373 = {maskExt_hi_373, maskExt_lo_373};
  wire [15:0]         maskExt_lo_374 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_374 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_374 = {maskExt_hi_374, maskExt_lo_374};
  wire [15:0]         maskExt_lo_375 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_375 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_375 = {maskExt_hi_375, maskExt_lo_375};
  wire [15:0]         maskExt_lo_376 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_376 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_376 = {maskExt_hi_376, maskExt_lo_376};
  wire [15:0]         maskExt_lo_377 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_377 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_377 = {maskExt_hi_377, maskExt_lo_377};
  wire [15:0]         maskExt_lo_378 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_378 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_378 = {maskExt_hi_378, maskExt_lo_378};
  wire [15:0]         maskExt_lo_379 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_379 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_379 = {maskExt_hi_379, maskExt_lo_379};
  wire [15:0]         maskExt_lo_380 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_380 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_380 = {maskExt_hi_380, maskExt_lo_380};
  wire [15:0]         maskExt_lo_381 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_381 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_381 = {maskExt_hi_381, maskExt_lo_381};
  wire [15:0]         maskExt_lo_382 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_382 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_382 = {maskExt_hi_382, maskExt_lo_382};
  wire [15:0]         maskExt_lo_383 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_383 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_383 = {maskExt_hi_383, maskExt_lo_383};
  wire [15:0]         maskExt_lo_384 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_384 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_384 = {maskExt_hi_384, maskExt_lo_384};
  wire [15:0]         maskExt_lo_385 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_385 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_385 = {maskExt_hi_385, maskExt_lo_385};
  wire [15:0]         maskExt_lo_386 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_386 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_386 = {maskExt_hi_386, maskExt_lo_386};
  wire [15:0]         maskExt_lo_387 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_387 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_387 = {maskExt_hi_387, maskExt_lo_387};
  wire [15:0]         maskExt_lo_388 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_388 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_388 = {maskExt_hi_388, maskExt_lo_388};
  wire [15:0]         maskExt_lo_389 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_389 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_389 = {maskExt_hi_389, maskExt_lo_389};
  wire [15:0]         maskExt_lo_390 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_390 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_390 = {maskExt_hi_390, maskExt_lo_390};
  wire [15:0]         maskExt_lo_391 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_391 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_391 = {maskExt_hi_391, maskExt_lo_391};
  wire [15:0]         maskExt_lo_392 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_392 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_392 = {maskExt_hi_392, maskExt_lo_392};
  wire [15:0]         maskExt_lo_393 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_393 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_393 = {maskExt_hi_393, maskExt_lo_393};
  wire [15:0]         maskExt_lo_394 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_394 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_394 = {maskExt_hi_394, maskExt_lo_394};
  wire [15:0]         maskExt_lo_395 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_395 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_395 = {maskExt_hi_395, maskExt_lo_395};
  wire [15:0]         maskExt_lo_396 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_396 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_396 = {maskExt_hi_396, maskExt_lo_396};
  wire [15:0]         maskExt_lo_397 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_397 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_397 = {maskExt_hi_397, maskExt_lo_397};
  wire [15:0]         maskExt_lo_398 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_398 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_398 = {maskExt_hi_398, maskExt_lo_398};
  wire [15:0]         maskExt_lo_399 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_399 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_399 = {maskExt_hi_399, maskExt_lo_399};
  wire [15:0]         maskExt_lo_400 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_400 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_400 = {maskExt_hi_400, maskExt_lo_400};
  wire [15:0]         maskExt_lo_401 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_401 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_401 = {maskExt_hi_401, maskExt_lo_401};
  wire [15:0]         maskExt_lo_402 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_402 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_402 = {maskExt_hi_402, maskExt_lo_402};
  wire [15:0]         maskExt_lo_403 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_403 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_403 = {maskExt_hi_403, maskExt_lo_403};
  wire [15:0]         maskExt_lo_404 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_404 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_404 = {maskExt_hi_404, maskExt_lo_404};
  wire [15:0]         maskExt_lo_405 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_405 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_405 = {maskExt_hi_405, maskExt_lo_405};
  wire [15:0]         maskExt_lo_406 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_406 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_406 = {maskExt_hi_406, maskExt_lo_406};
  wire [15:0]         maskExt_lo_407 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_407 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_407 = {maskExt_hi_407, maskExt_lo_407};
  wire [15:0]         maskExt_lo_408 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_408 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_408 = {maskExt_hi_408, maskExt_lo_408};
  wire [15:0]         maskExt_lo_409 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_409 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_409 = {maskExt_hi_409, maskExt_lo_409};
  wire [15:0]         maskExt_lo_410 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_410 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_410 = {maskExt_hi_410, maskExt_lo_410};
  wire [15:0]         maskExt_lo_411 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_411 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_411 = {maskExt_hi_411, maskExt_lo_411};
  wire [15:0]         maskExt_lo_412 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_412 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_412 = {maskExt_hi_412, maskExt_lo_412};
  wire [15:0]         maskExt_lo_413 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_413 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_413 = {maskExt_hi_413, maskExt_lo_413};
  wire [15:0]         maskExt_lo_414 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_414 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_414 = {maskExt_hi_414, maskExt_lo_414};
  wire [15:0]         maskExt_lo_415 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_415 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_415 = {maskExt_hi_415, maskExt_lo_415};
  wire [15:0]         maskExt_lo_416 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_416 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_416 = {maskExt_hi_416, maskExt_lo_416};
  wire [15:0]         maskExt_lo_417 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_417 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_417 = {maskExt_hi_417, maskExt_lo_417};
  wire [15:0]         maskExt_lo_418 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_418 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_418 = {maskExt_hi_418, maskExt_lo_418};
  wire [15:0]         maskExt_lo_419 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_419 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_419 = {maskExt_hi_419, maskExt_lo_419};
  wire [15:0]         maskExt_lo_420 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_420 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_420 = {maskExt_hi_420, maskExt_lo_420};
  wire [15:0]         maskExt_lo_421 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_421 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_421 = {maskExt_hi_421, maskExt_lo_421};
  wire [15:0]         maskExt_lo_422 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_422 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_422 = {maskExt_hi_422, maskExt_lo_422};
  wire [15:0]         maskExt_lo_423 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_423 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_423 = {maskExt_hi_423, maskExt_lo_423};
  wire [15:0]         maskExt_lo_424 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_424 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_424 = {maskExt_hi_424, maskExt_lo_424};
  wire [15:0]         maskExt_lo_425 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_425 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_425 = {maskExt_hi_425, maskExt_lo_425};
  wire [15:0]         maskExt_lo_426 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_426 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_426 = {maskExt_hi_426, maskExt_lo_426};
  wire [15:0]         maskExt_lo_427 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_427 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_427 = {maskExt_hi_427, maskExt_lo_427};
  wire [15:0]         maskExt_lo_428 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_428 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_428 = {maskExt_hi_428, maskExt_lo_428};
  wire [15:0]         maskExt_lo_429 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_429 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_429 = {maskExt_hi_429, maskExt_lo_429};
  wire [15:0]         maskExt_lo_430 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_430 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_430 = {maskExt_hi_430, maskExt_lo_430};
  wire [15:0]         maskExt_lo_431 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_431 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_431 = {maskExt_hi_431, maskExt_lo_431};
  wire [15:0]         maskExt_lo_432 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_432 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_432 = {maskExt_hi_432, maskExt_lo_432};
  wire [15:0]         maskExt_lo_433 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_433 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_433 = {maskExt_hi_433, maskExt_lo_433};
  wire [15:0]         maskExt_lo_434 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_434 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_434 = {maskExt_hi_434, maskExt_lo_434};
  wire [15:0]         maskExt_lo_435 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_435 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_435 = {maskExt_hi_435, maskExt_lo_435};
  wire [15:0]         maskExt_lo_436 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_436 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_436 = {maskExt_hi_436, maskExt_lo_436};
  wire [15:0]         maskExt_lo_437 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_437 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_437 = {maskExt_hi_437, maskExt_lo_437};
  wire [15:0]         maskExt_lo_438 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_438 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_438 = {maskExt_hi_438, maskExt_lo_438};
  wire [15:0]         maskExt_lo_439 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_439 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_439 = {maskExt_hi_439, maskExt_lo_439};
  wire [15:0]         maskExt_lo_440 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_440 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_440 = {maskExt_hi_440, maskExt_lo_440};
  wire [15:0]         maskExt_lo_441 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_441 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_441 = {maskExt_hi_441, maskExt_lo_441};
  wire [15:0]         maskExt_lo_442 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_442 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_442 = {maskExt_hi_442, maskExt_lo_442};
  wire [15:0]         maskExt_lo_443 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_443 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_443 = {maskExt_hi_443, maskExt_lo_443};
  wire [15:0]         maskExt_lo_444 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_444 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_444 = {maskExt_hi_444, maskExt_lo_444};
  wire [15:0]         maskExt_lo_445 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_445 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_445 = {maskExt_hi_445, maskExt_lo_445};
  wire [15:0]         maskExt_lo_446 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_446 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_446 = {maskExt_hi_446, maskExt_lo_446};
  wire [15:0]         maskExt_lo_447 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_447 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_447 = {maskExt_hi_447, maskExt_lo_447};
  wire [15:0]         maskExt_lo_448 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_448 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_448 = {maskExt_hi_448, maskExt_lo_448};
  wire [15:0]         maskExt_lo_449 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_449 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_449 = {maskExt_hi_449, maskExt_lo_449};
  wire [15:0]         maskExt_lo_450 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_450 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_450 = {maskExt_hi_450, maskExt_lo_450};
  wire [15:0]         maskExt_lo_451 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_451 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_451 = {maskExt_hi_451, maskExt_lo_451};
  wire [15:0]         maskExt_lo_452 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_452 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_452 = {maskExt_hi_452, maskExt_lo_452};
  wire [15:0]         maskExt_lo_453 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_453 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_453 = {maskExt_hi_453, maskExt_lo_453};
  wire [15:0]         maskExt_lo_454 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_454 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_454 = {maskExt_hi_454, maskExt_lo_454};
  wire [15:0]         maskExt_lo_455 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_455 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_455 = {maskExt_hi_455, maskExt_lo_455};
  wire [15:0]         maskExt_lo_456 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_456 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_456 = {maskExt_hi_456, maskExt_lo_456};
  wire [15:0]         maskExt_lo_457 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_457 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_457 = {maskExt_hi_457, maskExt_lo_457};
  wire [15:0]         maskExt_lo_458 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_458 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_458 = {maskExt_hi_458, maskExt_lo_458};
  wire [15:0]         maskExt_lo_459 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_459 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_459 = {maskExt_hi_459, maskExt_lo_459};
  wire [15:0]         maskExt_lo_460 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_460 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_460 = {maskExt_hi_460, maskExt_lo_460};
  wire [15:0]         maskExt_lo_461 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_461 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_461 = {maskExt_hi_461, maskExt_lo_461};
  wire [15:0]         maskExt_lo_462 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_462 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_462 = {maskExt_hi_462, maskExt_lo_462};
  wire [15:0]         maskExt_lo_463 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_463 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_463 = {maskExt_hi_463, maskExt_lo_463};
  wire [15:0]         maskExt_lo_464 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_464 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_464 = {maskExt_hi_464, maskExt_lo_464};
  wire [15:0]         maskExt_lo_465 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_465 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_465 = {maskExt_hi_465, maskExt_lo_465};
  wire [15:0]         maskExt_lo_466 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_466 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_466 = {maskExt_hi_466, maskExt_lo_466};
  wire [15:0]         maskExt_lo_467 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_467 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_467 = {maskExt_hi_467, maskExt_lo_467};
  wire [15:0]         maskExt_lo_468 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_468 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_468 = {maskExt_hi_468, maskExt_lo_468};
  wire [15:0]         maskExt_lo_469 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_469 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_469 = {maskExt_hi_469, maskExt_lo_469};
  wire [15:0]         maskExt_lo_470 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_470 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_470 = {maskExt_hi_470, maskExt_lo_470};
  wire [15:0]         maskExt_lo_471 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_471 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_471 = {maskExt_hi_471, maskExt_lo_471};
  wire [15:0]         maskExt_lo_472 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_472 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_472 = {maskExt_hi_472, maskExt_lo_472};
  wire [15:0]         maskExt_lo_473 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_473 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_473 = {maskExt_hi_473, maskExt_lo_473};
  wire [15:0]         maskExt_lo_474 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_474 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_474 = {maskExt_hi_474, maskExt_lo_474};
  wire [15:0]         maskExt_lo_475 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_475 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_475 = {maskExt_hi_475, maskExt_lo_475};
  wire [15:0]         maskExt_lo_476 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_476 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_476 = {maskExt_hi_476, maskExt_lo_476};
  wire [15:0]         maskExt_lo_477 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_477 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_477 = {maskExt_hi_477, maskExt_lo_477};
  wire [15:0]         maskExt_lo_478 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_478 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_478 = {maskExt_hi_478, maskExt_lo_478};
  wire [15:0]         maskExt_lo_479 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_479 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_479 = {maskExt_hi_479, maskExt_lo_479};
  wire [15:0]         maskExt_lo_480 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_480 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_480 = {maskExt_hi_480, maskExt_lo_480};
  wire [15:0]         maskExt_lo_481 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_481 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_481 = {maskExt_hi_481, maskExt_lo_481};
  wire [15:0]         maskExt_lo_482 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_482 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_482 = {maskExt_hi_482, maskExt_lo_482};
  wire [15:0]         maskExt_lo_483 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_483 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_483 = {maskExt_hi_483, maskExt_lo_483};
  wire [15:0]         maskExt_lo_484 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_484 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_484 = {maskExt_hi_484, maskExt_lo_484};
  wire [15:0]         maskExt_lo_485 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_485 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_485 = {maskExt_hi_485, maskExt_lo_485};
  wire [15:0]         maskExt_lo_486 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_486 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_486 = {maskExt_hi_486, maskExt_lo_486};
  wire [15:0]         maskExt_lo_487 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_487 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_487 = {maskExt_hi_487, maskExt_lo_487};
  wire [15:0]         maskExt_lo_488 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_488 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_488 = {maskExt_hi_488, maskExt_lo_488};
  wire [15:0]         maskExt_lo_489 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_489 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_489 = {maskExt_hi_489, maskExt_lo_489};
  wire [15:0]         maskExt_lo_490 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_490 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_490 = {maskExt_hi_490, maskExt_lo_490};
  wire [15:0]         maskExt_lo_491 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_491 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_491 = {maskExt_hi_491, maskExt_lo_491};
  wire [15:0]         maskExt_lo_492 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_492 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_492 = {maskExt_hi_492, maskExt_lo_492};
  wire [15:0]         maskExt_lo_493 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_493 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_493 = {maskExt_hi_493, maskExt_lo_493};
  wire [15:0]         maskExt_lo_494 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_494 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_494 = {maskExt_hi_494, maskExt_lo_494};
  wire [15:0]         maskExt_lo_495 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_495 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_495 = {maskExt_hi_495, maskExt_lo_495};
  wire [15:0]         maskExt_lo_496 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_496 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_496 = {maskExt_hi_496, maskExt_lo_496};
  wire [15:0]         maskExt_lo_497 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_497 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_497 = {maskExt_hi_497, maskExt_lo_497};
  wire [15:0]         maskExt_lo_498 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_498 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_498 = {maskExt_hi_498, maskExt_lo_498};
  wire [15:0]         maskExt_lo_499 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_499 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_499 = {maskExt_hi_499, maskExt_lo_499};
  wire [15:0]         maskExt_lo_500 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_500 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_500 = {maskExt_hi_500, maskExt_lo_500};
  wire [15:0]         maskExt_lo_501 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_501 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_501 = {maskExt_hi_501, maskExt_lo_501};
  wire [15:0]         maskExt_lo_502 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_502 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_502 = {maskExt_hi_502, maskExt_lo_502};
  wire [15:0]         maskExt_lo_503 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_503 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_503 = {maskExt_hi_503, maskExt_lo_503};
  wire [15:0]         maskExt_lo_504 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_504 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_504 = {maskExt_hi_504, maskExt_lo_504};
  wire [15:0]         maskExt_lo_505 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_505 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_505 = {maskExt_hi_505, maskExt_lo_505};
  wire [15:0]         maskExt_lo_506 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_506 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_506 = {maskExt_hi_506, maskExt_lo_506};
  wire [15:0]         maskExt_lo_507 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_507 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_507 = {maskExt_hi_507, maskExt_lo_507};
  wire [15:0]         maskExt_lo_508 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_508 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_508 = {maskExt_hi_508, maskExt_lo_508};
  wire [15:0]         maskExt_lo_509 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_509 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_509 = {maskExt_hi_509, maskExt_lo_509};
  wire [15:0]         maskExt_lo_510 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_510 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_510 = {maskExt_hi_510, maskExt_lo_510};
  wire [15:0]         maskExt_lo_511 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_511 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_511 = {maskExt_hi_511, maskExt_lo_511};
  wire [15:0]         maskExt_lo_512 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_512 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_512 = {maskExt_hi_512, maskExt_lo_512};
  wire [15:0]         maskExt_lo_513 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_513 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_513 = {maskExt_hi_513, maskExt_lo_513};
  wire [15:0]         maskExt_lo_514 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_514 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_514 = {maskExt_hi_514, maskExt_lo_514};
  wire [15:0]         maskExt_lo_515 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_515 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_515 = {maskExt_hi_515, maskExt_lo_515};
  wire [15:0]         maskExt_lo_516 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_516 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_516 = {maskExt_hi_516, maskExt_lo_516};
  wire [15:0]         maskExt_lo_517 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_517 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_517 = {maskExt_hi_517, maskExt_lo_517};
  wire [15:0]         maskExt_lo_518 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_518 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_518 = {maskExt_hi_518, maskExt_lo_518};
  wire [15:0]         maskExt_lo_519 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_519 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_519 = {maskExt_hi_519, maskExt_lo_519};
  wire [15:0]         maskExt_lo_520 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_520 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_520 = {maskExt_hi_520, maskExt_lo_520};
  wire [15:0]         maskExt_lo_521 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_521 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_521 = {maskExt_hi_521, maskExt_lo_521};
  wire [15:0]         maskExt_lo_522 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_522 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_522 = {maskExt_hi_522, maskExt_lo_522};
  wire [15:0]         maskExt_lo_523 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_523 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_523 = {maskExt_hi_523, maskExt_lo_523};
  wire [15:0]         maskExt_lo_524 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_524 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_524 = {maskExt_hi_524, maskExt_lo_524};
  wire [15:0]         maskExt_lo_525 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_525 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_525 = {maskExt_hi_525, maskExt_lo_525};
  wire [15:0]         maskExt_lo_526 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_526 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_526 = {maskExt_hi_526, maskExt_lo_526};
  wire [15:0]         maskExt_lo_527 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_527 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_527 = {maskExt_hi_527, maskExt_lo_527};
  wire [15:0]         maskExt_lo_528 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_528 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_528 = {maskExt_hi_528, maskExt_lo_528};
  wire [15:0]         maskExt_lo_529 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_529 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_529 = {maskExt_hi_529, maskExt_lo_529};
  wire [15:0]         maskExt_lo_530 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_530 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_530 = {maskExt_hi_530, maskExt_lo_530};
  wire [15:0]         maskExt_lo_531 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_531 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_531 = {maskExt_hi_531, maskExt_lo_531};
  wire [15:0]         maskExt_lo_532 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_532 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_532 = {maskExt_hi_532, maskExt_lo_532};
  wire [15:0]         maskExt_lo_533 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_533 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_533 = {maskExt_hi_533, maskExt_lo_533};
  wire [15:0]         maskExt_lo_534 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_534 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_534 = {maskExt_hi_534, maskExt_lo_534};
  wire [15:0]         maskExt_lo_535 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_535 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_535 = {maskExt_hi_535, maskExt_lo_535};
  wire [15:0]         maskExt_lo_536 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_536 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_536 = {maskExt_hi_536, maskExt_lo_536};
  wire [15:0]         maskExt_lo_537 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_537 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_537 = {maskExt_hi_537, maskExt_lo_537};
  wire [15:0]         maskExt_lo_538 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_538 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_538 = {maskExt_hi_538, maskExt_lo_538};
  wire [15:0]         maskExt_lo_539 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_539 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_539 = {maskExt_hi_539, maskExt_lo_539};
  wire [15:0]         maskExt_lo_540 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_540 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_540 = {maskExt_hi_540, maskExt_lo_540};
  wire [15:0]         maskExt_lo_541 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_541 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_541 = {maskExt_hi_541, maskExt_lo_541};
  wire [15:0]         maskExt_lo_542 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_542 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_542 = {maskExt_hi_542, maskExt_lo_542};
  wire [15:0]         maskExt_lo_543 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_543 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_543 = {maskExt_hi_543, maskExt_lo_543};
  wire [15:0]         maskExt_lo_544 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_544 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_544 = {maskExt_hi_544, maskExt_lo_544};
  wire [15:0]         maskExt_lo_545 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_545 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_545 = {maskExt_hi_545, maskExt_lo_545};
  wire [15:0]         maskExt_lo_546 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_546 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_546 = {maskExt_hi_546, maskExt_lo_546};
  wire [15:0]         maskExt_lo_547 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_547 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_547 = {maskExt_hi_547, maskExt_lo_547};
  wire [15:0]         maskExt_lo_548 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_548 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_548 = {maskExt_hi_548, maskExt_lo_548};
  wire [15:0]         maskExt_lo_549 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_549 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_549 = {maskExt_hi_549, maskExt_lo_549};
  wire [15:0]         maskExt_lo_550 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_550 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_550 = {maskExt_hi_550, maskExt_lo_550};
  wire [15:0]         maskExt_lo_551 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_551 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_551 = {maskExt_hi_551, maskExt_lo_551};
  wire [15:0]         maskExt_lo_552 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_552 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_552 = {maskExt_hi_552, maskExt_lo_552};
  wire [15:0]         maskExt_lo_553 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_553 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_553 = {maskExt_hi_553, maskExt_lo_553};
  wire [15:0]         maskExt_lo_554 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_554 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_554 = {maskExt_hi_554, maskExt_lo_554};
  wire [15:0]         maskExt_lo_555 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_555 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_555 = {maskExt_hi_555, maskExt_lo_555};
  wire [15:0]         maskExt_lo_556 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_556 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_556 = {maskExt_hi_556, maskExt_lo_556};
  wire [15:0]         maskExt_lo_557 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_557 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_557 = {maskExt_hi_557, maskExt_lo_557};
  wire [15:0]         maskExt_lo_558 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_558 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_558 = {maskExt_hi_558, maskExt_lo_558};
  wire [15:0]         maskExt_lo_559 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_559 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_559 = {maskExt_hi_559, maskExt_lo_559};
  wire [15:0]         maskExt_lo_560 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_560 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_560 = {maskExt_hi_560, maskExt_lo_560};
  wire [15:0]         maskExt_lo_561 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_561 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_561 = {maskExt_hi_561, maskExt_lo_561};
  wire [15:0]         maskExt_lo_562 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_562 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_562 = {maskExt_hi_562, maskExt_lo_562};
  wire [15:0]         maskExt_lo_563 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_563 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_563 = {maskExt_hi_563, maskExt_lo_563};
  wire [15:0]         maskExt_lo_564 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_564 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_564 = {maskExt_hi_564, maskExt_lo_564};
  wire [15:0]         maskExt_lo_565 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_565 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_565 = {maskExt_hi_565, maskExt_lo_565};
  wire [15:0]         maskExt_lo_566 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_566 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_566 = {maskExt_hi_566, maskExt_lo_566};
  wire [15:0]         maskExt_lo_567 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_567 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_567 = {maskExt_hi_567, maskExt_lo_567};
  wire [15:0]         maskExt_lo_568 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_568 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_568 = {maskExt_hi_568, maskExt_lo_568};
  wire [15:0]         maskExt_lo_569 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_569 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_569 = {maskExt_hi_569, maskExt_lo_569};
  wire [15:0]         maskExt_lo_570 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_570 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_570 = {maskExt_hi_570, maskExt_lo_570};
  wire [15:0]         maskExt_lo_571 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_571 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_571 = {maskExt_hi_571, maskExt_lo_571};
  wire [15:0]         maskExt_lo_572 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_572 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_572 = {maskExt_hi_572, maskExt_lo_572};
  wire [15:0]         maskExt_lo_573 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_573 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_573 = {maskExt_hi_573, maskExt_lo_573};
  wire [15:0]         maskExt_lo_574 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_574 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_574 = {maskExt_hi_574, maskExt_lo_574};
  wire [15:0]         maskExt_lo_575 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_575 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_575 = {maskExt_hi_575, maskExt_lo_575};
  wire [15:0]         maskExt_lo_576 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_576 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_576 = {maskExt_hi_576, maskExt_lo_576};
  wire [15:0]         maskExt_lo_577 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_577 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_577 = {maskExt_hi_577, maskExt_lo_577};
  wire [15:0]         maskExt_lo_578 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_578 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_578 = {maskExt_hi_578, maskExt_lo_578};
  wire [15:0]         maskExt_lo_579 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_579 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_579 = {maskExt_hi_579, maskExt_lo_579};
  wire [15:0]         maskExt_lo_580 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_580 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_580 = {maskExt_hi_580, maskExt_lo_580};
  wire [15:0]         maskExt_lo_581 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_581 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_581 = {maskExt_hi_581, maskExt_lo_581};
  wire [15:0]         maskExt_lo_582 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_582 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_582 = {maskExt_hi_582, maskExt_lo_582};
  wire [15:0]         maskExt_lo_583 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_583 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_583 = {maskExt_hi_583, maskExt_lo_583};
  wire [15:0]         maskExt_lo_584 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_584 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_584 = {maskExt_hi_584, maskExt_lo_584};
  wire [15:0]         maskExt_lo_585 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_585 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_585 = {maskExt_hi_585, maskExt_lo_585};
  wire [15:0]         maskExt_lo_586 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_586 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_586 = {maskExt_hi_586, maskExt_lo_586};
  wire [15:0]         maskExt_lo_587 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_587 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_587 = {maskExt_hi_587, maskExt_lo_587};
  wire [15:0]         maskExt_lo_588 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_588 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_588 = {maskExt_hi_588, maskExt_lo_588};
  wire [15:0]         maskExt_lo_589 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_589 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_589 = {maskExt_hi_589, maskExt_lo_589};
  wire [15:0]         maskExt_lo_590 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_590 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_590 = {maskExt_hi_590, maskExt_lo_590};
  wire [15:0]         maskExt_lo_591 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_591 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_591 = {maskExt_hi_591, maskExt_lo_591};
  wire [15:0]         maskExt_lo_592 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_592 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_592 = {maskExt_hi_592, maskExt_lo_592};
  wire [15:0]         maskExt_lo_593 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_593 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_593 = {maskExt_hi_593, maskExt_lo_593};
  wire [15:0]         maskExt_lo_594 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_594 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_594 = {maskExt_hi_594, maskExt_lo_594};
  wire [15:0]         maskExt_lo_595 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_595 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_595 = {maskExt_hi_595, maskExt_lo_595};
  wire [15:0]         maskExt_lo_596 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_596 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_596 = {maskExt_hi_596, maskExt_lo_596};
  wire [15:0]         maskExt_lo_597 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_597 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_597 = {maskExt_hi_597, maskExt_lo_597};
  wire [15:0]         maskExt_lo_598 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_598 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_598 = {maskExt_hi_598, maskExt_lo_598};
  wire [15:0]         maskExt_lo_599 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_599 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_599 = {maskExt_hi_599, maskExt_lo_599};
  wire [15:0]         maskExt_lo_600 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_600 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_600 = {maskExt_hi_600, maskExt_lo_600};
  wire [15:0]         maskExt_lo_601 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_601 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_601 = {maskExt_hi_601, maskExt_lo_601};
  wire [15:0]         maskExt_lo_602 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_602 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_602 = {maskExt_hi_602, maskExt_lo_602};
  wire [15:0]         maskExt_lo_603 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_603 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_603 = {maskExt_hi_603, maskExt_lo_603};
  wire [15:0]         maskExt_lo_604 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_604 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_604 = {maskExt_hi_604, maskExt_lo_604};
  wire [15:0]         maskExt_lo_605 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_605 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_605 = {maskExt_hi_605, maskExt_lo_605};
  wire [15:0]         maskExt_lo_606 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_606 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_606 = {maskExt_hi_606, maskExt_lo_606};
  wire [15:0]         maskExt_lo_607 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_607 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_607 = {maskExt_hi_607, maskExt_lo_607};
  wire [15:0]         maskExt_lo_608 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_608 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_608 = {maskExt_hi_608, maskExt_lo_608};
  wire [15:0]         maskExt_lo_609 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_609 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_609 = {maskExt_hi_609, maskExt_lo_609};
  wire [15:0]         maskExt_lo_610 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_610 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_610 = {maskExt_hi_610, maskExt_lo_610};
  wire [15:0]         maskExt_lo_611 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_611 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_611 = {maskExt_hi_611, maskExt_lo_611};
  wire [15:0]         maskExt_lo_612 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_612 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_612 = {maskExt_hi_612, maskExt_lo_612};
  wire [15:0]         maskExt_lo_613 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_613 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_613 = {maskExt_hi_613, maskExt_lo_613};
  wire [15:0]         maskExt_lo_614 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_614 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_614 = {maskExt_hi_614, maskExt_lo_614};
  wire [15:0]         maskExt_lo_615 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_615 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_615 = {maskExt_hi_615, maskExt_lo_615};
  wire [15:0]         maskExt_lo_616 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_616 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_616 = {maskExt_hi_616, maskExt_lo_616};
  wire [15:0]         maskExt_lo_617 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_617 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_617 = {maskExt_hi_617, maskExt_lo_617};
  wire [15:0]         maskExt_lo_618 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_618 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_618 = {maskExt_hi_618, maskExt_lo_618};
  wire [15:0]         maskExt_lo_619 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_619 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_619 = {maskExt_hi_619, maskExt_lo_619};
  wire [15:0]         maskExt_lo_620 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_620 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_620 = {maskExt_hi_620, maskExt_lo_620};
  wire [15:0]         maskExt_lo_621 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_621 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_621 = {maskExt_hi_621, maskExt_lo_621};
  wire [15:0]         maskExt_lo_622 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_622 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_622 = {maskExt_hi_622, maskExt_lo_622};
  wire [15:0]         maskExt_lo_623 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_623 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_623 = {maskExt_hi_623, maskExt_lo_623};
  wire [15:0]         maskExt_lo_624 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_624 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_624 = {maskExt_hi_624, maskExt_lo_624};
  wire [15:0]         maskExt_lo_625 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_625 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_625 = {maskExt_hi_625, maskExt_lo_625};
  wire [15:0]         maskExt_lo_626 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_626 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_626 = {maskExt_hi_626, maskExt_lo_626};
  wire [15:0]         maskExt_lo_627 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_627 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_627 = {maskExt_hi_627, maskExt_lo_627};
  wire [15:0]         maskExt_lo_628 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_628 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_628 = {maskExt_hi_628, maskExt_lo_628};
  wire [15:0]         maskExt_lo_629 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_629 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_629 = {maskExt_hi_629, maskExt_lo_629};
  wire [15:0]         maskExt_lo_630 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_630 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_630 = {maskExt_hi_630, maskExt_lo_630};
  wire [15:0]         maskExt_lo_631 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_631 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_631 = {maskExt_hi_631, maskExt_lo_631};
  wire [15:0]         maskExt_lo_632 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_632 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_632 = {maskExt_hi_632, maskExt_lo_632};
  wire [15:0]         maskExt_lo_633 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_633 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_633 = {maskExt_hi_633, maskExt_lo_633};
  wire [15:0]         maskExt_lo_634 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_634 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_634 = {maskExt_hi_634, maskExt_lo_634};
  wire [15:0]         maskExt_lo_635 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_635 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_635 = {maskExt_hi_635, maskExt_lo_635};
  wire [15:0]         maskExt_lo_636 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_636 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_636 = {maskExt_hi_636, maskExt_lo_636};
  wire [15:0]         maskExt_lo_637 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_637 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_637 = {maskExt_hi_637, maskExt_lo_637};
  wire [15:0]         maskExt_lo_638 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_638 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_638 = {maskExt_hi_638, maskExt_lo_638};
  wire [15:0]         maskExt_lo_639 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_639 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_639 = {maskExt_hi_639, maskExt_lo_639};
  wire [15:0]         maskExt_lo_640 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_640 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_640 = {maskExt_hi_640, maskExt_lo_640};
  wire [15:0]         maskExt_lo_641 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_641 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_641 = {maskExt_hi_641, maskExt_lo_641};
  wire [15:0]         maskExt_lo_642 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_642 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_642 = {maskExt_hi_642, maskExt_lo_642};
  wire [15:0]         maskExt_lo_643 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_643 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_643 = {maskExt_hi_643, maskExt_lo_643};
  wire [15:0]         maskExt_lo_644 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_644 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_644 = {maskExt_hi_644, maskExt_lo_644};
  wire [15:0]         maskExt_lo_645 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_645 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_645 = {maskExt_hi_645, maskExt_lo_645};
  wire [15:0]         maskExt_lo_646 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_646 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_646 = {maskExt_hi_646, maskExt_lo_646};
  wire [15:0]         maskExt_lo_647 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_647 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_647 = {maskExt_hi_647, maskExt_lo_647};
  wire [15:0]         maskExt_lo_648 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_648 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_648 = {maskExt_hi_648, maskExt_lo_648};
  wire [15:0]         maskExt_lo_649 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_649 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_649 = {maskExt_hi_649, maskExt_lo_649};
  wire [15:0]         maskExt_lo_650 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_650 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_650 = {maskExt_hi_650, maskExt_lo_650};
  wire [15:0]         maskExt_lo_651 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_651 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_651 = {maskExt_hi_651, maskExt_lo_651};
  wire [15:0]         maskExt_lo_652 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_652 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_652 = {maskExt_hi_652, maskExt_lo_652};
  wire [15:0]         maskExt_lo_653 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_653 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_653 = {maskExt_hi_653, maskExt_lo_653};
  wire [15:0]         maskExt_lo_654 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_654 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_654 = {maskExt_hi_654, maskExt_lo_654};
  wire [15:0]         maskExt_lo_655 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_655 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_655 = {maskExt_hi_655, maskExt_lo_655};
  wire [15:0]         maskExt_lo_656 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_656 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_656 = {maskExt_hi_656, maskExt_lo_656};
  wire [15:0]         maskExt_lo_657 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_657 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_657 = {maskExt_hi_657, maskExt_lo_657};
  wire [15:0]         maskExt_lo_658 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_658 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_658 = {maskExt_hi_658, maskExt_lo_658};
  wire [15:0]         maskExt_lo_659 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_659 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_659 = {maskExt_hi_659, maskExt_lo_659};
  wire [15:0]         maskExt_lo_660 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_660 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_660 = {maskExt_hi_660, maskExt_lo_660};
  wire [15:0]         maskExt_lo_661 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_661 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_661 = {maskExt_hi_661, maskExt_lo_661};
  wire [15:0]         maskExt_lo_662 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_662 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_662 = {maskExt_hi_662, maskExt_lo_662};
  wire [15:0]         maskExt_lo_663 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_663 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_663 = {maskExt_hi_663, maskExt_lo_663};
  wire [15:0]         maskExt_lo_664 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_664 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_664 = {maskExt_hi_664, maskExt_lo_664};
  wire [15:0]         maskExt_lo_665 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_665 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_665 = {maskExt_hi_665, maskExt_lo_665};
  wire [15:0]         maskExt_lo_666 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_666 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_666 = {maskExt_hi_666, maskExt_lo_666};
  wire [15:0]         maskExt_lo_667 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_667 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_667 = {maskExt_hi_667, maskExt_lo_667};
  wire [15:0]         maskExt_lo_668 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_668 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_668 = {maskExt_hi_668, maskExt_lo_668};
  wire [15:0]         maskExt_lo_669 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_669 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_669 = {maskExt_hi_669, maskExt_lo_669};
  wire [15:0]         maskExt_lo_670 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_670 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_670 = {maskExt_hi_670, maskExt_lo_670};
  wire [15:0]         maskExt_lo_671 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_671 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_671 = {maskExt_hi_671, maskExt_lo_671};
  wire [15:0]         maskExt_lo_672 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_672 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_672 = {maskExt_hi_672, maskExt_lo_672};
  wire [15:0]         maskExt_lo_673 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_673 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_673 = {maskExt_hi_673, maskExt_lo_673};
  wire [15:0]         maskExt_lo_674 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_674 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_674 = {maskExt_hi_674, maskExt_lo_674};
  wire [15:0]         maskExt_lo_675 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_675 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_675 = {maskExt_hi_675, maskExt_lo_675};
  wire [15:0]         maskExt_lo_676 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_676 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_676 = {maskExt_hi_676, maskExt_lo_676};
  wire [15:0]         maskExt_lo_677 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_677 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_677 = {maskExt_hi_677, maskExt_lo_677};
  wire [15:0]         maskExt_lo_678 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_678 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_678 = {maskExt_hi_678, maskExt_lo_678};
  wire [15:0]         maskExt_lo_679 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_679 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_679 = {maskExt_hi_679, maskExt_lo_679};
  wire [15:0]         maskExt_lo_680 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_680 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_680 = {maskExt_hi_680, maskExt_lo_680};
  wire [15:0]         maskExt_lo_681 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_681 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_681 = {maskExt_hi_681, maskExt_lo_681};
  wire [15:0]         maskExt_lo_682 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_682 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_682 = {maskExt_hi_682, maskExt_lo_682};
  wire [15:0]         maskExt_lo_683 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_683 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_683 = {maskExt_hi_683, maskExt_lo_683};
  wire [15:0]         maskExt_lo_684 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_684 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_684 = {maskExt_hi_684, maskExt_lo_684};
  wire [15:0]         maskExt_lo_685 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_685 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_685 = {maskExt_hi_685, maskExt_lo_685};
  wire [15:0]         maskExt_lo_686 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_686 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_686 = {maskExt_hi_686, maskExt_lo_686};
  wire [15:0]         maskExt_lo_687 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_687 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_687 = {maskExt_hi_687, maskExt_lo_687};
  wire [15:0]         maskExt_lo_688 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_688 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_688 = {maskExt_hi_688, maskExt_lo_688};
  wire [15:0]         maskExt_lo_689 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_689 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_689 = {maskExt_hi_689, maskExt_lo_689};
  wire [15:0]         maskExt_lo_690 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_690 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_690 = {maskExt_hi_690, maskExt_lo_690};
  wire [15:0]         maskExt_lo_691 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_691 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_691 = {maskExt_hi_691, maskExt_lo_691};
  wire [15:0]         maskExt_lo_692 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_692 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_692 = {maskExt_hi_692, maskExt_lo_692};
  wire [15:0]         maskExt_lo_693 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_693 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_693 = {maskExt_hi_693, maskExt_lo_693};
  wire [15:0]         maskExt_lo_694 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_694 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_694 = {maskExt_hi_694, maskExt_lo_694};
  wire [15:0]         maskExt_lo_695 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_695 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_695 = {maskExt_hi_695, maskExt_lo_695};
  wire [15:0]         maskExt_lo_696 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_696 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_696 = {maskExt_hi_696, maskExt_lo_696};
  wire [15:0]         maskExt_lo_697 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_697 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_697 = {maskExt_hi_697, maskExt_lo_697};
  wire [15:0]         maskExt_lo_698 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_698 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_698 = {maskExt_hi_698, maskExt_lo_698};
  wire [15:0]         maskExt_lo_699 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_699 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_699 = {maskExt_hi_699, maskExt_lo_699};
  wire [15:0]         maskExt_lo_700 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_700 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_700 = {maskExt_hi_700, maskExt_lo_700};
  wire [15:0]         maskExt_lo_701 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_701 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_701 = {maskExt_hi_701, maskExt_lo_701};
  wire [15:0]         maskExt_lo_702 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_702 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_702 = {maskExt_hi_702, maskExt_lo_702};
  wire [15:0]         maskExt_lo_703 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_703 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_703 = {maskExt_hi_703, maskExt_lo_703};
  wire [15:0]         maskExt_lo_704 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_704 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_704 = {maskExt_hi_704, maskExt_lo_704};
  wire [15:0]         maskExt_lo_705 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_705 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_705 = {maskExt_hi_705, maskExt_lo_705};
  wire [15:0]         maskExt_lo_706 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_706 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_706 = {maskExt_hi_706, maskExt_lo_706};
  wire [15:0]         maskExt_lo_707 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_707 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_707 = {maskExt_hi_707, maskExt_lo_707};
  wire [15:0]         maskExt_lo_708 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_708 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_708 = {maskExt_hi_708, maskExt_lo_708};
  wire [15:0]         maskExt_lo_709 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_709 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_709 = {maskExt_hi_709, maskExt_lo_709};
  wire [15:0]         maskExt_lo_710 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_710 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_710 = {maskExt_hi_710, maskExt_lo_710};
  wire [15:0]         maskExt_lo_711 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_711 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_711 = {maskExt_hi_711, maskExt_lo_711};
  wire [15:0]         maskExt_lo_712 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_712 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_712 = {maskExt_hi_712, maskExt_lo_712};
  wire [15:0]         maskExt_lo_713 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_713 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_713 = {maskExt_hi_713, maskExt_lo_713};
  wire [15:0]         maskExt_lo_714 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_714 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_714 = {maskExt_hi_714, maskExt_lo_714};
  wire [15:0]         maskExt_lo_715 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_715 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_715 = {maskExt_hi_715, maskExt_lo_715};
  wire [15:0]         maskExt_lo_716 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_716 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_716 = {maskExt_hi_716, maskExt_lo_716};
  wire [15:0]         maskExt_lo_717 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_717 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_717 = {maskExt_hi_717, maskExt_lo_717};
  wire [15:0]         maskExt_lo_718 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_718 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_718 = {maskExt_hi_718, maskExt_lo_718};
  wire [15:0]         maskExt_lo_719 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_719 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_719 = {maskExt_hi_719, maskExt_lo_719};
  wire [15:0]         maskExt_lo_720 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_720 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_720 = {maskExt_hi_720, maskExt_lo_720};
  wire [15:0]         maskExt_lo_721 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_721 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_721 = {maskExt_hi_721, maskExt_lo_721};
  wire [15:0]         maskExt_lo_722 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_722 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_722 = {maskExt_hi_722, maskExt_lo_722};
  wire [15:0]         maskExt_lo_723 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_723 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_723 = {maskExt_hi_723, maskExt_lo_723};
  wire [15:0]         maskExt_lo_724 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_724 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_724 = {maskExt_hi_724, maskExt_lo_724};
  wire [15:0]         maskExt_lo_725 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_725 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_725 = {maskExt_hi_725, maskExt_lo_725};
  wire [15:0]         maskExt_lo_726 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_726 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_726 = {maskExt_hi_726, maskExt_lo_726};
  wire [15:0]         maskExt_lo_727 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_727 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_727 = {maskExt_hi_727, maskExt_lo_727};
  wire [15:0]         maskExt_lo_728 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_728 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_728 = {maskExt_hi_728, maskExt_lo_728};
  wire [15:0]         maskExt_lo_729 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_729 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_729 = {maskExt_hi_729, maskExt_lo_729};
  wire [15:0]         maskExt_lo_730 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_730 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_730 = {maskExt_hi_730, maskExt_lo_730};
  wire [15:0]         maskExt_lo_731 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_731 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_731 = {maskExt_hi_731, maskExt_lo_731};
  wire [15:0]         maskExt_lo_732 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_732 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_732 = {maskExt_hi_732, maskExt_lo_732};
  wire [15:0]         maskExt_lo_733 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_733 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_733 = {maskExt_hi_733, maskExt_lo_733};
  wire [15:0]         maskExt_lo_734 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_734 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_734 = {maskExt_hi_734, maskExt_lo_734};
  wire [15:0]         maskExt_lo_735 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_735 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_735 = {maskExt_hi_735, maskExt_lo_735};
  wire [15:0]         maskExt_lo_736 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_736 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_736 = {maskExt_hi_736, maskExt_lo_736};
  wire [15:0]         maskExt_lo_737 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_737 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_737 = {maskExt_hi_737, maskExt_lo_737};
  wire [15:0]         maskExt_lo_738 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_738 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_738 = {maskExt_hi_738, maskExt_lo_738};
  wire [15:0]         maskExt_lo_739 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_739 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_739 = {maskExt_hi_739, maskExt_lo_739};
  wire [15:0]         maskExt_lo_740 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_740 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_740 = {maskExt_hi_740, maskExt_lo_740};
  wire [15:0]         maskExt_lo_741 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_741 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_741 = {maskExt_hi_741, maskExt_lo_741};
  wire [15:0]         maskExt_lo_742 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_742 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_742 = {maskExt_hi_742, maskExt_lo_742};
  wire [15:0]         maskExt_lo_743 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_743 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_743 = {maskExt_hi_743, maskExt_lo_743};
  wire [15:0]         maskExt_lo_744 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_744 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_744 = {maskExt_hi_744, maskExt_lo_744};
  wire [15:0]         maskExt_lo_745 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_745 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_745 = {maskExt_hi_745, maskExt_lo_745};
  wire [15:0]         maskExt_lo_746 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_746 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_746 = {maskExt_hi_746, maskExt_lo_746};
  wire [15:0]         maskExt_lo_747 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_747 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_747 = {maskExt_hi_747, maskExt_lo_747};
  wire [15:0]         maskExt_lo_748 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_748 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_748 = {maskExt_hi_748, maskExt_lo_748};
  wire [15:0]         maskExt_lo_749 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_749 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_749 = {maskExt_hi_749, maskExt_lo_749};
  wire [15:0]         maskExt_lo_750 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_750 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_750 = {maskExt_hi_750, maskExt_lo_750};
  wire [15:0]         maskExt_lo_751 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_751 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_751 = {maskExt_hi_751, maskExt_lo_751};
  wire [15:0]         maskExt_lo_752 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_752 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_752 = {maskExt_hi_752, maskExt_lo_752};
  wire [15:0]         maskExt_lo_753 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_753 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_753 = {maskExt_hi_753, maskExt_lo_753};
  wire [15:0]         maskExt_lo_754 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_754 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_754 = {maskExt_hi_754, maskExt_lo_754};
  wire [15:0]         maskExt_lo_755 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_755 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_755 = {maskExt_hi_755, maskExt_lo_755};
  wire [15:0]         maskExt_lo_756 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_756 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_756 = {maskExt_hi_756, maskExt_lo_756};
  wire [15:0]         maskExt_lo_757 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_757 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_757 = {maskExt_hi_757, maskExt_lo_757};
  wire [15:0]         maskExt_lo_758 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_758 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_758 = {maskExt_hi_758, maskExt_lo_758};
  wire [15:0]         maskExt_lo_759 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_759 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_759 = {maskExt_hi_759, maskExt_lo_759};
  wire [15:0]         maskExt_lo_760 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_760 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_760 = {maskExt_hi_760, maskExt_lo_760};
  wire [15:0]         maskExt_lo_761 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_761 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_761 = {maskExt_hi_761, maskExt_lo_761};
  wire [15:0]         maskExt_lo_762 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_762 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_762 = {maskExt_hi_762, maskExt_lo_762};
  wire [15:0]         maskExt_lo_763 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_763 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_763 = {maskExt_hi_763, maskExt_lo_763};
  wire [15:0]         maskExt_lo_764 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_764 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_764 = {maskExt_hi_764, maskExt_lo_764};
  wire [15:0]         maskExt_lo_765 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_765 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_765 = {maskExt_hi_765, maskExt_lo_765};
  wire [15:0]         maskExt_lo_766 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_766 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_766 = {maskExt_hi_766, maskExt_lo_766};
  wire [15:0]         maskExt_lo_767 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_767 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_767 = {maskExt_hi_767, maskExt_lo_767};
  wire [15:0]         maskExt_lo_768 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_768 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_768 = {maskExt_hi_768, maskExt_lo_768};
  wire [15:0]         maskExt_lo_769 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_769 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_769 = {maskExt_hi_769, maskExt_lo_769};
  wire [15:0]         maskExt_lo_770 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_770 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_770 = {maskExt_hi_770, maskExt_lo_770};
  wire [15:0]         maskExt_lo_771 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_771 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_771 = {maskExt_hi_771, maskExt_lo_771};
  wire [15:0]         maskExt_lo_772 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_772 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_772 = {maskExt_hi_772, maskExt_lo_772};
  wire [15:0]         maskExt_lo_773 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_773 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_773 = {maskExt_hi_773, maskExt_lo_773};
  wire [15:0]         maskExt_lo_774 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_774 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_774 = {maskExt_hi_774, maskExt_lo_774};
  wire [15:0]         maskExt_lo_775 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_775 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_775 = {maskExt_hi_775, maskExt_lo_775};
  wire [15:0]         maskExt_lo_776 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_776 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_776 = {maskExt_hi_776, maskExt_lo_776};
  wire [15:0]         maskExt_lo_777 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_777 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_777 = {maskExt_hi_777, maskExt_lo_777};
  wire [15:0]         maskExt_lo_778 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_778 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_778 = {maskExt_hi_778, maskExt_lo_778};
  wire [15:0]         maskExt_lo_779 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_779 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_779 = {maskExt_hi_779, maskExt_lo_779};
  wire [15:0]         maskExt_lo_780 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_780 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_780 = {maskExt_hi_780, maskExt_lo_780};
  wire [15:0]         maskExt_lo_781 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_781 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_781 = {maskExt_hi_781, maskExt_lo_781};
  wire [15:0]         maskExt_lo_782 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_782 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_782 = {maskExt_hi_782, maskExt_lo_782};
  wire [15:0]         maskExt_lo_783 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_783 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_783 = {maskExt_hi_783, maskExt_lo_783};
  wire [15:0]         maskExt_lo_784 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_784 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_784 = {maskExt_hi_784, maskExt_lo_784};
  wire [15:0]         maskExt_lo_785 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_785 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_785 = {maskExt_hi_785, maskExt_lo_785};
  wire [15:0]         maskExt_lo_786 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_786 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_786 = {maskExt_hi_786, maskExt_lo_786};
  wire [15:0]         maskExt_lo_787 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_787 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_787 = {maskExt_hi_787, maskExt_lo_787};
  wire [15:0]         maskExt_lo_788 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_788 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_788 = {maskExt_hi_788, maskExt_lo_788};
  wire [15:0]         maskExt_lo_789 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_789 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_789 = {maskExt_hi_789, maskExt_lo_789};
  wire [15:0]         maskExt_lo_790 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_790 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_790 = {maskExt_hi_790, maskExt_lo_790};
  wire [15:0]         maskExt_lo_791 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_791 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_791 = {maskExt_hi_791, maskExt_lo_791};
  wire [15:0]         maskExt_lo_792 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_792 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_792 = {maskExt_hi_792, maskExt_lo_792};
  wire [15:0]         maskExt_lo_793 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_793 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_793 = {maskExt_hi_793, maskExt_lo_793};
  wire [15:0]         maskExt_lo_794 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_794 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_794 = {maskExt_hi_794, maskExt_lo_794};
  wire [15:0]         maskExt_lo_795 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_795 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_795 = {maskExt_hi_795, maskExt_lo_795};
  wire [15:0]         maskExt_lo_796 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_796 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_796 = {maskExt_hi_796, maskExt_lo_796};
  wire [15:0]         maskExt_lo_797 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_797 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_797 = {maskExt_hi_797, maskExt_lo_797};
  wire [15:0]         maskExt_lo_798 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_798 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_798 = {maskExt_hi_798, maskExt_lo_798};
  wire [15:0]         maskExt_lo_799 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_799 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_799 = {maskExt_hi_799, maskExt_lo_799};
  wire [15:0]         maskExt_lo_800 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_800 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_800 = {maskExt_hi_800, maskExt_lo_800};
  wire [15:0]         maskExt_lo_801 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_801 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_801 = {maskExt_hi_801, maskExt_lo_801};
  wire [15:0]         maskExt_lo_802 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_802 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_802 = {maskExt_hi_802, maskExt_lo_802};
  wire [15:0]         maskExt_lo_803 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_803 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_803 = {maskExt_hi_803, maskExt_lo_803};
  wire [15:0]         maskExt_lo_804 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_804 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_804 = {maskExt_hi_804, maskExt_lo_804};
  wire [15:0]         maskExt_lo_805 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_805 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_805 = {maskExt_hi_805, maskExt_lo_805};
  wire [15:0]         maskExt_lo_806 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_806 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_806 = {maskExt_hi_806, maskExt_lo_806};
  wire [15:0]         maskExt_lo_807 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_807 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_807 = {maskExt_hi_807, maskExt_lo_807};
  wire [15:0]         maskExt_lo_808 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_808 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_808 = {maskExt_hi_808, maskExt_lo_808};
  wire [15:0]         maskExt_lo_809 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_809 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_809 = {maskExt_hi_809, maskExt_lo_809};
  wire [15:0]         maskExt_lo_810 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_810 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_810 = {maskExt_hi_810, maskExt_lo_810};
  wire [15:0]         maskExt_lo_811 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_811 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_811 = {maskExt_hi_811, maskExt_lo_811};
  wire [15:0]         maskExt_lo_812 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_812 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_812 = {maskExt_hi_812, maskExt_lo_812};
  wire [15:0]         maskExt_lo_813 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_813 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_813 = {maskExt_hi_813, maskExt_lo_813};
  wire [15:0]         maskExt_lo_814 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_814 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_814 = {maskExt_hi_814, maskExt_lo_814};
  wire [15:0]         maskExt_lo_815 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_815 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_815 = {maskExt_hi_815, maskExt_lo_815};
  wire [15:0]         maskExt_lo_816 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_816 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_816 = {maskExt_hi_816, maskExt_lo_816};
  wire [15:0]         maskExt_lo_817 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_817 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_817 = {maskExt_hi_817, maskExt_lo_817};
  wire [15:0]         maskExt_lo_818 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_818 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_818 = {maskExt_hi_818, maskExt_lo_818};
  wire [15:0]         maskExt_lo_819 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_819 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_819 = {maskExt_hi_819, maskExt_lo_819};
  wire [15:0]         maskExt_lo_820 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_820 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_820 = {maskExt_hi_820, maskExt_lo_820};
  wire [15:0]         maskExt_lo_821 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_821 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_821 = {maskExt_hi_821, maskExt_lo_821};
  wire [15:0]         maskExt_lo_822 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_822 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_822 = {maskExt_hi_822, maskExt_lo_822};
  wire [15:0]         maskExt_lo_823 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_823 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_823 = {maskExt_hi_823, maskExt_lo_823};
  wire [15:0]         maskExt_lo_824 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_824 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_824 = {maskExt_hi_824, maskExt_lo_824};
  wire [15:0]         maskExt_lo_825 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_825 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_825 = {maskExt_hi_825, maskExt_lo_825};
  wire [15:0]         maskExt_lo_826 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_826 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_826 = {maskExt_hi_826, maskExt_lo_826};
  wire [15:0]         maskExt_lo_827 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_827 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_827 = {maskExt_hi_827, maskExt_lo_827};
  wire [15:0]         maskExt_lo_828 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_828 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_828 = {maskExt_hi_828, maskExt_lo_828};
  wire [15:0]         maskExt_lo_829 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_829 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_829 = {maskExt_hi_829, maskExt_lo_829};
  wire [15:0]         maskExt_lo_830 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_830 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_830 = {maskExt_hi_830, maskExt_lo_830};
  wire [15:0]         maskExt_lo_831 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_831 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_831 = {maskExt_hi_831, maskExt_lo_831};
  wire [15:0]         maskExt_lo_832 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_832 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_832 = {maskExt_hi_832, maskExt_lo_832};
  wire [15:0]         maskExt_lo_833 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_833 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_833 = {maskExt_hi_833, maskExt_lo_833};
  wire [15:0]         maskExt_lo_834 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_834 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_834 = {maskExt_hi_834, maskExt_lo_834};
  wire [15:0]         maskExt_lo_835 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_835 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_835 = {maskExt_hi_835, maskExt_lo_835};
  wire [15:0]         maskExt_lo_836 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_836 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_836 = {maskExt_hi_836, maskExt_lo_836};
  wire [15:0]         maskExt_lo_837 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_837 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_837 = {maskExt_hi_837, maskExt_lo_837};
  wire [15:0]         maskExt_lo_838 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_838 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_838 = {maskExt_hi_838, maskExt_lo_838};
  wire [15:0]         maskExt_lo_839 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_839 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_839 = {maskExt_hi_839, maskExt_lo_839};
  wire [15:0]         maskExt_lo_840 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_840 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_840 = {maskExt_hi_840, maskExt_lo_840};
  wire [15:0]         maskExt_lo_841 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_841 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_841 = {maskExt_hi_841, maskExt_lo_841};
  wire [15:0]         maskExt_lo_842 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_842 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_842 = {maskExt_hi_842, maskExt_lo_842};
  wire [15:0]         maskExt_lo_843 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_843 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_843 = {maskExt_hi_843, maskExt_lo_843};
  wire [15:0]         maskExt_lo_844 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_844 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_844 = {maskExt_hi_844, maskExt_lo_844};
  wire [15:0]         maskExt_lo_845 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_845 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_845 = {maskExt_hi_845, maskExt_lo_845};
  wire [15:0]         maskExt_lo_846 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_846 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_846 = {maskExt_hi_846, maskExt_lo_846};
  wire [15:0]         maskExt_lo_847 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_847 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_847 = {maskExt_hi_847, maskExt_lo_847};
  wire [15:0]         maskExt_lo_848 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_848 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_848 = {maskExt_hi_848, maskExt_lo_848};
  wire [15:0]         maskExt_lo_849 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_849 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_849 = {maskExt_hi_849, maskExt_lo_849};
  wire [15:0]         maskExt_lo_850 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_850 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_850 = {maskExt_hi_850, maskExt_lo_850};
  wire [15:0]         maskExt_lo_851 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_851 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_851 = {maskExt_hi_851, maskExt_lo_851};
  wire [15:0]         maskExt_lo_852 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_852 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_852 = {maskExt_hi_852, maskExt_lo_852};
  wire [15:0]         maskExt_lo_853 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_853 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_853 = {maskExt_hi_853, maskExt_lo_853};
  wire [15:0]         maskExt_lo_854 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_854 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_854 = {maskExt_hi_854, maskExt_lo_854};
  wire [15:0]         maskExt_lo_855 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_855 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_855 = {maskExt_hi_855, maskExt_lo_855};
  wire [15:0]         maskExt_lo_856 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_856 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_856 = {maskExt_hi_856, maskExt_lo_856};
  wire [15:0]         maskExt_lo_857 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_857 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_857 = {maskExt_hi_857, maskExt_lo_857};
  wire [15:0]         maskExt_lo_858 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_858 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_858 = {maskExt_hi_858, maskExt_lo_858};
  wire [15:0]         maskExt_lo_859 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_859 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_859 = {maskExt_hi_859, maskExt_lo_859};
  wire [15:0]         maskExt_lo_860 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_860 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_860 = {maskExt_hi_860, maskExt_lo_860};
  wire [15:0]         maskExt_lo_861 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_861 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_861 = {maskExt_hi_861, maskExt_lo_861};
  wire [15:0]         maskExt_lo_862 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_862 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_862 = {maskExt_hi_862, maskExt_lo_862};
  wire [15:0]         maskExt_lo_863 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_863 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_863 = {maskExt_hi_863, maskExt_lo_863};
  wire [15:0]         maskExt_lo_864 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_864 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_864 = {maskExt_hi_864, maskExt_lo_864};
  wire [15:0]         maskExt_lo_865 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_865 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_865 = {maskExt_hi_865, maskExt_lo_865};
  wire [15:0]         maskExt_lo_866 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_866 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_866 = {maskExt_hi_866, maskExt_lo_866};
  wire [15:0]         maskExt_lo_867 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_867 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_867 = {maskExt_hi_867, maskExt_lo_867};
  wire [15:0]         maskExt_lo_868 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_868 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_868 = {maskExt_hi_868, maskExt_lo_868};
  wire [15:0]         maskExt_lo_869 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_869 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_869 = {maskExt_hi_869, maskExt_lo_869};
  wire [15:0]         maskExt_lo_870 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_870 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_870 = {maskExt_hi_870, maskExt_lo_870};
  wire [15:0]         maskExt_lo_871 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_871 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_871 = {maskExt_hi_871, maskExt_lo_871};
  wire [15:0]         maskExt_lo_872 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_872 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_872 = {maskExt_hi_872, maskExt_lo_872};
  wire [15:0]         maskExt_lo_873 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_873 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_873 = {maskExt_hi_873, maskExt_lo_873};
  wire [15:0]         maskExt_lo_874 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_874 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_874 = {maskExt_hi_874, maskExt_lo_874};
  wire [15:0]         maskExt_lo_875 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_875 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_875 = {maskExt_hi_875, maskExt_lo_875};
  wire [15:0]         maskExt_lo_876 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_876 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_876 = {maskExt_hi_876, maskExt_lo_876};
  wire [15:0]         maskExt_lo_877 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_877 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_877 = {maskExt_hi_877, maskExt_lo_877};
  wire [15:0]         maskExt_lo_878 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_878 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_878 = {maskExt_hi_878, maskExt_lo_878};
  wire [15:0]         maskExt_lo_879 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_879 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_879 = {maskExt_hi_879, maskExt_lo_879};
  wire [15:0]         maskExt_lo_880 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_880 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_880 = {maskExt_hi_880, maskExt_lo_880};
  wire [15:0]         maskExt_lo_881 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_881 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_881 = {maskExt_hi_881, maskExt_lo_881};
  wire [15:0]         maskExt_lo_882 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_882 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_882 = {maskExt_hi_882, maskExt_lo_882};
  wire [15:0]         maskExt_lo_883 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_883 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_883 = {maskExt_hi_883, maskExt_lo_883};
  wire [15:0]         maskExt_lo_884 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_884 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_884 = {maskExt_hi_884, maskExt_lo_884};
  wire [15:0]         maskExt_lo_885 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_885 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_885 = {maskExt_hi_885, maskExt_lo_885};
  wire [15:0]         maskExt_lo_886 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_886 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_886 = {maskExt_hi_886, maskExt_lo_886};
  wire [15:0]         maskExt_lo_887 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_887 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_887 = {maskExt_hi_887, maskExt_lo_887};
  wire [15:0]         maskExt_lo_888 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_888 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_888 = {maskExt_hi_888, maskExt_lo_888};
  wire [15:0]         maskExt_lo_889 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_889 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_889 = {maskExt_hi_889, maskExt_lo_889};
  wire [15:0]         maskExt_lo_890 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_890 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_890 = {maskExt_hi_890, maskExt_lo_890};
  wire [15:0]         maskExt_lo_891 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_891 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_891 = {maskExt_hi_891, maskExt_lo_891};
  wire [15:0]         maskExt_lo_892 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_892 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_892 = {maskExt_hi_892, maskExt_lo_892};
  wire [15:0]         maskExt_lo_893 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_893 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_893 = {maskExt_hi_893, maskExt_lo_893};
  wire [15:0]         maskExt_lo_894 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_894 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_894 = {maskExt_hi_894, maskExt_lo_894};
  wire [15:0]         maskExt_lo_895 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_895 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_895 = {maskExt_hi_895, maskExt_lo_895};
  wire [15:0]         maskExt_lo_896 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_896 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_896 = {maskExt_hi_896, maskExt_lo_896};
  wire [15:0]         maskExt_lo_897 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_897 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_897 = {maskExt_hi_897, maskExt_lo_897};
  wire [15:0]         maskExt_lo_898 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_898 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_898 = {maskExt_hi_898, maskExt_lo_898};
  wire [15:0]         maskExt_lo_899 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_899 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_899 = {maskExt_hi_899, maskExt_lo_899};
  wire [15:0]         maskExt_lo_900 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_900 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_900 = {maskExt_hi_900, maskExt_lo_900};
  wire [15:0]         maskExt_lo_901 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_901 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_901 = {maskExt_hi_901, maskExt_lo_901};
  wire [15:0]         maskExt_lo_902 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_902 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_902 = {maskExt_hi_902, maskExt_lo_902};
  wire [15:0]         maskExt_lo_903 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_903 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_903 = {maskExt_hi_903, maskExt_lo_903};
  wire [15:0]         maskExt_lo_904 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_904 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_904 = {maskExt_hi_904, maskExt_lo_904};
  wire [15:0]         maskExt_lo_905 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_905 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_905 = {maskExt_hi_905, maskExt_lo_905};
  wire [15:0]         maskExt_lo_906 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_906 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_906 = {maskExt_hi_906, maskExt_lo_906};
  wire [15:0]         maskExt_lo_907 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_907 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_907 = {maskExt_hi_907, maskExt_lo_907};
  wire [15:0]         maskExt_lo_908 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_908 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_908 = {maskExt_hi_908, maskExt_lo_908};
  wire [15:0]         maskExt_lo_909 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_909 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_909 = {maskExt_hi_909, maskExt_lo_909};
  wire [15:0]         maskExt_lo_910 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_910 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_910 = {maskExt_hi_910, maskExt_lo_910};
  wire [15:0]         maskExt_lo_911 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_911 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_911 = {maskExt_hi_911, maskExt_lo_911};
  wire [15:0]         maskExt_lo_912 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_912 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_912 = {maskExt_hi_912, maskExt_lo_912};
  wire [15:0]         maskExt_lo_913 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_913 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_913 = {maskExt_hi_913, maskExt_lo_913};
  wire [15:0]         maskExt_lo_914 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_914 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_914 = {maskExt_hi_914, maskExt_lo_914};
  wire [15:0]         maskExt_lo_915 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_915 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_915 = {maskExt_hi_915, maskExt_lo_915};
  wire [15:0]         maskExt_lo_916 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_916 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_916 = {maskExt_hi_916, maskExt_lo_916};
  wire [15:0]         maskExt_lo_917 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_917 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_917 = {maskExt_hi_917, maskExt_lo_917};
  wire [15:0]         maskExt_lo_918 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_918 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_918 = {maskExt_hi_918, maskExt_lo_918};
  wire [15:0]         maskExt_lo_919 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_919 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_919 = {maskExt_hi_919, maskExt_lo_919};
  wire [15:0]         maskExt_lo_920 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_920 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_920 = {maskExt_hi_920, maskExt_lo_920};
  wire [15:0]         maskExt_lo_921 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_921 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_921 = {maskExt_hi_921, maskExt_lo_921};
  wire [15:0]         maskExt_lo_922 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_922 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_922 = {maskExt_hi_922, maskExt_lo_922};
  wire [15:0]         maskExt_lo_923 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_923 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_923 = {maskExt_hi_923, maskExt_lo_923};
  wire [15:0]         maskExt_lo_924 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_924 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_924 = {maskExt_hi_924, maskExt_lo_924};
  wire [15:0]         maskExt_lo_925 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_925 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_925 = {maskExt_hi_925, maskExt_lo_925};
  wire [15:0]         maskExt_lo_926 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_926 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_926 = {maskExt_hi_926, maskExt_lo_926};
  wire [15:0]         maskExt_lo_927 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_927 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_927 = {maskExt_hi_927, maskExt_lo_927};
  wire [15:0]         maskExt_lo_928 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_928 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_928 = {maskExt_hi_928, maskExt_lo_928};
  wire [15:0]         maskExt_lo_929 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_929 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_929 = {maskExt_hi_929, maskExt_lo_929};
  wire [15:0]         maskExt_lo_930 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_930 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_930 = {maskExt_hi_930, maskExt_lo_930};
  wire [15:0]         maskExt_lo_931 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_931 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_931 = {maskExt_hi_931, maskExt_lo_931};
  wire [15:0]         maskExt_lo_932 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_932 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_932 = {maskExt_hi_932, maskExt_lo_932};
  wire [15:0]         maskExt_lo_933 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_933 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_933 = {maskExt_hi_933, maskExt_lo_933};
  wire [15:0]         maskExt_lo_934 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_934 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_934 = {maskExt_hi_934, maskExt_lo_934};
  wire [15:0]         maskExt_lo_935 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_935 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_935 = {maskExt_hi_935, maskExt_lo_935};
  wire [15:0]         maskExt_lo_936 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_936 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_936 = {maskExt_hi_936, maskExt_lo_936};
  wire [15:0]         maskExt_lo_937 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_937 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_937 = {maskExt_hi_937, maskExt_lo_937};
  wire [15:0]         maskExt_lo_938 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_938 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_938 = {maskExt_hi_938, maskExt_lo_938};
  wire [15:0]         maskExt_lo_939 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_939 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_939 = {maskExt_hi_939, maskExt_lo_939};
  wire [15:0]         maskExt_lo_940 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_940 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_940 = {maskExt_hi_940, maskExt_lo_940};
  wire [15:0]         maskExt_lo_941 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_941 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_941 = {maskExt_hi_941, maskExt_lo_941};
  wire [15:0]         maskExt_lo_942 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_942 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_942 = {maskExt_hi_942, maskExt_lo_942};
  wire [15:0]         maskExt_lo_943 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_943 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_943 = {maskExt_hi_943, maskExt_lo_943};
  wire [15:0]         maskExt_lo_944 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_944 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_944 = {maskExt_hi_944, maskExt_lo_944};
  wire [15:0]         maskExt_lo_945 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_945 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_945 = {maskExt_hi_945, maskExt_lo_945};
  wire [15:0]         maskExt_lo_946 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_946 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_946 = {maskExt_hi_946, maskExt_lo_946};
  wire [15:0]         maskExt_lo_947 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_947 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_947 = {maskExt_hi_947, maskExt_lo_947};
  wire [15:0]         maskExt_lo_948 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_948 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_948 = {maskExt_hi_948, maskExt_lo_948};
  wire [15:0]         maskExt_lo_949 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_949 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_949 = {maskExt_hi_949, maskExt_lo_949};
  wire [15:0]         maskExt_lo_950 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_950 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_950 = {maskExt_hi_950, maskExt_lo_950};
  wire [15:0]         maskExt_lo_951 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_951 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_951 = {maskExt_hi_951, maskExt_lo_951};
  wire [15:0]         maskExt_lo_952 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_952 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_952 = {maskExt_hi_952, maskExt_lo_952};
  wire [15:0]         maskExt_lo_953 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_953 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_953 = {maskExt_hi_953, maskExt_lo_953};
  wire [15:0]         maskExt_lo_954 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_954 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_954 = {maskExt_hi_954, maskExt_lo_954};
  wire [15:0]         maskExt_lo_955 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_955 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_955 = {maskExt_hi_955, maskExt_lo_955};
  wire [15:0]         maskExt_lo_956 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_956 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_956 = {maskExt_hi_956, maskExt_lo_956};
  wire [15:0]         maskExt_lo_957 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_957 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_957 = {maskExt_hi_957, maskExt_lo_957};
  wire [15:0]         maskExt_lo_958 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_958 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_958 = {maskExt_hi_958, maskExt_lo_958};
  wire [15:0]         maskExt_lo_959 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_959 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_959 = {maskExt_hi_959, maskExt_lo_959};
  wire [15:0]         maskExt_lo_960 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_960 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_960 = {maskExt_hi_960, maskExt_lo_960};
  wire [15:0]         maskExt_lo_961 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_961 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_961 = {maskExt_hi_961, maskExt_lo_961};
  wire [15:0]         maskExt_lo_962 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_962 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_962 = {maskExt_hi_962, maskExt_lo_962};
  wire [15:0]         maskExt_lo_963 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_963 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_963 = {maskExt_hi_963, maskExt_lo_963};
  wire [15:0]         maskExt_lo_964 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_964 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_964 = {maskExt_hi_964, maskExt_lo_964};
  wire [15:0]         maskExt_lo_965 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_965 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_965 = {maskExt_hi_965, maskExt_lo_965};
  wire [15:0]         maskExt_lo_966 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_966 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_966 = {maskExt_hi_966, maskExt_lo_966};
  wire [15:0]         maskExt_lo_967 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_967 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_967 = {maskExt_hi_967, maskExt_lo_967};
  wire [15:0]         maskExt_lo_968 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_968 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_968 = {maskExt_hi_968, maskExt_lo_968};
  wire [15:0]         maskExt_lo_969 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_969 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_969 = {maskExt_hi_969, maskExt_lo_969};
  wire [15:0]         maskExt_lo_970 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_970 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_970 = {maskExt_hi_970, maskExt_lo_970};
  wire [15:0]         maskExt_lo_971 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_971 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_971 = {maskExt_hi_971, maskExt_lo_971};
  wire [15:0]         maskExt_lo_972 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_972 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_972 = {maskExt_hi_972, maskExt_lo_972};
  wire [15:0]         maskExt_lo_973 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_973 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_973 = {maskExt_hi_973, maskExt_lo_973};
  wire [15:0]         maskExt_lo_974 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_974 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_974 = {maskExt_hi_974, maskExt_lo_974};
  wire [15:0]         maskExt_lo_975 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_975 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_975 = {maskExt_hi_975, maskExt_lo_975};
  wire [15:0]         maskExt_lo_976 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_976 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_976 = {maskExt_hi_976, maskExt_lo_976};
  wire [15:0]         maskExt_lo_977 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_977 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_977 = {maskExt_hi_977, maskExt_lo_977};
  wire [15:0]         maskExt_lo_978 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_978 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_978 = {maskExt_hi_978, maskExt_lo_978};
  wire [15:0]         maskExt_lo_979 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_979 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_979 = {maskExt_hi_979, maskExt_lo_979};
  wire [15:0]         maskExt_lo_980 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_980 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_980 = {maskExt_hi_980, maskExt_lo_980};
  wire [15:0]         maskExt_lo_981 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_981 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_981 = {maskExt_hi_981, maskExt_lo_981};
  wire [15:0]         maskExt_lo_982 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_982 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_982 = {maskExt_hi_982, maskExt_lo_982};
  wire [15:0]         maskExt_lo_983 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_983 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_983 = {maskExt_hi_983, maskExt_lo_983};
  wire [15:0]         maskExt_lo_984 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_984 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_984 = {maskExt_hi_984, maskExt_lo_984};
  wire [15:0]         maskExt_lo_985 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_985 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_985 = {maskExt_hi_985, maskExt_lo_985};
  wire [15:0]         maskExt_lo_986 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_986 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_986 = {maskExt_hi_986, maskExt_lo_986};
  wire [15:0]         maskExt_lo_987 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_987 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_987 = {maskExt_hi_987, maskExt_lo_987};
  wire [15:0]         maskExt_lo_988 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_988 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_988 = {maskExt_hi_988, maskExt_lo_988};
  wire [15:0]         maskExt_lo_989 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_989 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_989 = {maskExt_hi_989, maskExt_lo_989};
  wire [15:0]         maskExt_lo_990 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_990 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_990 = {maskExt_hi_990, maskExt_lo_990};
  wire [15:0]         maskExt_lo_991 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_991 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_991 = {maskExt_hi_991, maskExt_lo_991};
  wire [15:0]         maskExt_lo_992 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_992 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_992 = {maskExt_hi_992, maskExt_lo_992};
  wire [15:0]         maskExt_lo_993 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_993 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_993 = {maskExt_hi_993, maskExt_lo_993};
  wire [15:0]         maskExt_lo_994 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_994 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_994 = {maskExt_hi_994, maskExt_lo_994};
  wire [15:0]         maskExt_lo_995 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_995 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_995 = {maskExt_hi_995, maskExt_lo_995};
  wire [15:0]         maskExt_lo_996 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_996 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_996 = {maskExt_hi_996, maskExt_lo_996};
  wire [15:0]         maskExt_lo_997 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_997 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_997 = {maskExt_hi_997, maskExt_lo_997};
  wire [15:0]         maskExt_lo_998 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_998 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_998 = {maskExt_hi_998, maskExt_lo_998};
  wire [15:0]         maskExt_lo_999 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_999 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_999 = {maskExt_hi_999, maskExt_lo_999};
  wire [15:0]         maskExt_lo_1000 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1000 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1000 = {maskExt_hi_1000, maskExt_lo_1000};
  wire [15:0]         maskExt_lo_1001 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1001 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1001 = {maskExt_hi_1001, maskExt_lo_1001};
  wire [15:0]         maskExt_lo_1002 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1002 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1002 = {maskExt_hi_1002, maskExt_lo_1002};
  wire [15:0]         maskExt_lo_1003 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1003 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1003 = {maskExt_hi_1003, maskExt_lo_1003};
  wire [15:0]         maskExt_lo_1004 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1004 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1004 = {maskExt_hi_1004, maskExt_lo_1004};
  wire [15:0]         maskExt_lo_1005 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1005 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1005 = {maskExt_hi_1005, maskExt_lo_1005};
  wire [15:0]         maskExt_lo_1006 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1006 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1006 = {maskExt_hi_1006, maskExt_lo_1006};
  wire [15:0]         maskExt_lo_1007 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1007 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1007 = {maskExt_hi_1007, maskExt_lo_1007};
  wire [15:0]         maskExt_lo_1008 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1008 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1008 = {maskExt_hi_1008, maskExt_lo_1008};
  wire [15:0]         maskExt_lo_1009 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1009 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1009 = {maskExt_hi_1009, maskExt_lo_1009};
  wire [15:0]         maskExt_lo_1010 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1010 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1010 = {maskExt_hi_1010, maskExt_lo_1010};
  wire [15:0]         maskExt_lo_1011 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1011 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1011 = {maskExt_hi_1011, maskExt_lo_1011};
  wire [15:0]         maskExt_lo_1012 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1012 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1012 = {maskExt_hi_1012, maskExt_lo_1012};
  wire [15:0]         maskExt_lo_1013 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1013 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1013 = {maskExt_hi_1013, maskExt_lo_1013};
  wire [15:0]         maskExt_lo_1014 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1014 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1014 = {maskExt_hi_1014, maskExt_lo_1014};
  wire [15:0]         maskExt_lo_1015 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1015 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1015 = {maskExt_hi_1015, maskExt_lo_1015};
  wire [15:0]         maskExt_lo_1016 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1016 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1016 = {maskExt_hi_1016, maskExt_lo_1016};
  wire [15:0]         maskExt_lo_1017 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1017 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1017 = {maskExt_hi_1017, maskExt_lo_1017};
  wire [15:0]         maskExt_lo_1018 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1018 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1018 = {maskExt_hi_1018, maskExt_lo_1018};
  wire [15:0]         maskExt_lo_1019 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1019 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1019 = {maskExt_hi_1019, maskExt_lo_1019};
  wire [15:0]         maskExt_lo_1020 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1020 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1020 = {maskExt_hi_1020, maskExt_lo_1020};
  wire [15:0]         maskExt_lo_1021 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1021 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1021 = {maskExt_hi_1021, maskExt_lo_1021};
  wire [15:0]         maskExt_lo_1022 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1022 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1022 = {maskExt_hi_1022, maskExt_lo_1022};
  wire [15:0]         maskExt_lo_1023 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1023 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1023 = {maskExt_hi_1023, maskExt_lo_1023};
  wire [15:0]         maskExt_lo_1024 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1024 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1024 = {maskExt_hi_1024, maskExt_lo_1024};
  wire [15:0]         maskExt_lo_1025 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1025 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1025 = {maskExt_hi_1025, maskExt_lo_1025};
  wire [15:0]         maskExt_lo_1026 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1026 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1026 = {maskExt_hi_1026, maskExt_lo_1026};
  wire [15:0]         maskExt_lo_1027 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1027 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1027 = {maskExt_hi_1027, maskExt_lo_1027};
  wire [15:0]         maskExt_lo_1028 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1028 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1028 = {maskExt_hi_1028, maskExt_lo_1028};
  wire [15:0]         maskExt_lo_1029 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1029 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1029 = {maskExt_hi_1029, maskExt_lo_1029};
  wire [15:0]         maskExt_lo_1030 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1030 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1030 = {maskExt_hi_1030, maskExt_lo_1030};
  wire [15:0]         maskExt_lo_1031 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1031 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1031 = {maskExt_hi_1031, maskExt_lo_1031};
  wire [15:0]         maskExt_lo_1032 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1032 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1032 = {maskExt_hi_1032, maskExt_lo_1032};
  wire [15:0]         maskExt_lo_1033 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1033 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1033 = {maskExt_hi_1033, maskExt_lo_1033};
  wire [15:0]         maskExt_lo_1034 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1034 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1034 = {maskExt_hi_1034, maskExt_lo_1034};
  wire [15:0]         maskExt_lo_1035 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1035 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1035 = {maskExt_hi_1035, maskExt_lo_1035};
  wire [15:0]         maskExt_lo_1036 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1036 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1036 = {maskExt_hi_1036, maskExt_lo_1036};
  wire [15:0]         maskExt_lo_1037 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1037 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1037 = {maskExt_hi_1037, maskExt_lo_1037};
  wire [15:0]         maskExt_lo_1038 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1038 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1038 = {maskExt_hi_1038, maskExt_lo_1038};
  wire [15:0]         maskExt_lo_1039 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1039 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1039 = {maskExt_hi_1039, maskExt_lo_1039};
  wire [15:0]         maskExt_lo_1040 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1040 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1040 = {maskExt_hi_1040, maskExt_lo_1040};
  wire [15:0]         maskExt_lo_1041 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1041 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1041 = {maskExt_hi_1041, maskExt_lo_1041};
  wire [15:0]         maskExt_lo_1042 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1042 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1042 = {maskExt_hi_1042, maskExt_lo_1042};
  wire [15:0]         maskExt_lo_1043 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1043 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1043 = {maskExt_hi_1043, maskExt_lo_1043};
  wire [15:0]         maskExt_lo_1044 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1044 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1044 = {maskExt_hi_1044, maskExt_lo_1044};
  wire [15:0]         maskExt_lo_1045 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1045 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1045 = {maskExt_hi_1045, maskExt_lo_1045};
  wire [15:0]         maskExt_lo_1046 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1046 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1046 = {maskExt_hi_1046, maskExt_lo_1046};
  wire [15:0]         maskExt_lo_1047 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1047 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1047 = {maskExt_hi_1047, maskExt_lo_1047};
  wire [15:0]         maskExt_lo_1048 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1048 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1048 = {maskExt_hi_1048, maskExt_lo_1048};
  wire [15:0]         maskExt_lo_1049 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1049 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1049 = {maskExt_hi_1049, maskExt_lo_1049};
  wire [15:0]         maskExt_lo_1050 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1050 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1050 = {maskExt_hi_1050, maskExt_lo_1050};
  wire [15:0]         maskExt_lo_1051 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1051 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1051 = {maskExt_hi_1051, maskExt_lo_1051};
  wire [15:0]         maskExt_lo_1052 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1052 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1052 = {maskExt_hi_1052, maskExt_lo_1052};
  wire [15:0]         maskExt_lo_1053 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1053 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1053 = {maskExt_hi_1053, maskExt_lo_1053};
  wire [15:0]         maskExt_lo_1054 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1054 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1054 = {maskExt_hi_1054, maskExt_lo_1054};
  wire [15:0]         maskExt_lo_1055 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1055 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1055 = {maskExt_hi_1055, maskExt_lo_1055};
  wire [15:0]         maskExt_lo_1056 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1056 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1056 = {maskExt_hi_1056, maskExt_lo_1056};
  wire [15:0]         maskExt_lo_1057 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1057 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1057 = {maskExt_hi_1057, maskExt_lo_1057};
  wire [15:0]         maskExt_lo_1058 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1058 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1058 = {maskExt_hi_1058, maskExt_lo_1058};
  wire [15:0]         maskExt_lo_1059 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1059 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1059 = {maskExt_hi_1059, maskExt_lo_1059};
  wire [15:0]         maskExt_lo_1060 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1060 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1060 = {maskExt_hi_1060, maskExt_lo_1060};
  wire [15:0]         maskExt_lo_1061 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1061 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1061 = {maskExt_hi_1061, maskExt_lo_1061};
  wire [15:0]         maskExt_lo_1062 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1062 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1062 = {maskExt_hi_1062, maskExt_lo_1062};
  wire [15:0]         maskExt_lo_1063 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1063 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1063 = {maskExt_hi_1063, maskExt_lo_1063};
  wire [15:0]         maskExt_lo_1064 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1064 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1064 = {maskExt_hi_1064, maskExt_lo_1064};
  wire [15:0]         maskExt_lo_1065 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1065 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1065 = {maskExt_hi_1065, maskExt_lo_1065};
  wire [15:0]         maskExt_lo_1066 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1066 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1066 = {maskExt_hi_1066, maskExt_lo_1066};
  wire [15:0]         maskExt_lo_1067 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1067 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1067 = {maskExt_hi_1067, maskExt_lo_1067};
  wire [15:0]         maskExt_lo_1068 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1068 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1068 = {maskExt_hi_1068, maskExt_lo_1068};
  wire [15:0]         maskExt_lo_1069 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1069 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1069 = {maskExt_hi_1069, maskExt_lo_1069};
  wire [15:0]         maskExt_lo_1070 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1070 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1070 = {maskExt_hi_1070, maskExt_lo_1070};
  wire [15:0]         maskExt_lo_1071 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1071 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1071 = {maskExt_hi_1071, maskExt_lo_1071};
  wire [15:0]         maskExt_lo_1072 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1072 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1072 = {maskExt_hi_1072, maskExt_lo_1072};
  wire [15:0]         maskExt_lo_1073 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1073 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1073 = {maskExt_hi_1073, maskExt_lo_1073};
  wire [15:0]         maskExt_lo_1074 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1074 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1074 = {maskExt_hi_1074, maskExt_lo_1074};
  wire [15:0]         maskExt_lo_1075 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1075 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1075 = {maskExt_hi_1075, maskExt_lo_1075};
  wire [15:0]         maskExt_lo_1076 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1076 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1076 = {maskExt_hi_1076, maskExt_lo_1076};
  wire [15:0]         maskExt_lo_1077 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1077 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1077 = {maskExt_hi_1077, maskExt_lo_1077};
  wire [15:0]         maskExt_lo_1078 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1078 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1078 = {maskExt_hi_1078, maskExt_lo_1078};
  wire [15:0]         maskExt_lo_1079 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1079 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1079 = {maskExt_hi_1079, maskExt_lo_1079};
  wire [15:0]         maskExt_lo_1080 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1080 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1080 = {maskExt_hi_1080, maskExt_lo_1080};
  wire [15:0]         maskExt_lo_1081 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1081 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1081 = {maskExt_hi_1081, maskExt_lo_1081};
  wire [15:0]         maskExt_lo_1082 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1082 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1082 = {maskExt_hi_1082, maskExt_lo_1082};
  wire [15:0]         maskExt_lo_1083 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1083 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1083 = {maskExt_hi_1083, maskExt_lo_1083};
  wire [15:0]         maskExt_lo_1084 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1084 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1084 = {maskExt_hi_1084, maskExt_lo_1084};
  wire [15:0]         maskExt_lo_1085 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1085 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1085 = {maskExt_hi_1085, maskExt_lo_1085};
  wire [15:0]         maskExt_lo_1086 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1086 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1086 = {maskExt_hi_1086, maskExt_lo_1086};
  wire [15:0]         maskExt_lo_1087 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1087 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1087 = {maskExt_hi_1087, maskExt_lo_1087};
  wire [15:0]         maskExt_lo_1088 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1088 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1088 = {maskExt_hi_1088, maskExt_lo_1088};
  wire [15:0]         maskExt_lo_1089 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1089 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1089 = {maskExt_hi_1089, maskExt_lo_1089};
  wire [15:0]         maskExt_lo_1090 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1090 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1090 = {maskExt_hi_1090, maskExt_lo_1090};
  wire [15:0]         maskExt_lo_1091 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1091 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1091 = {maskExt_hi_1091, maskExt_lo_1091};
  wire [15:0]         maskExt_lo_1092 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1092 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1092 = {maskExt_hi_1092, maskExt_lo_1092};
  wire [15:0]         maskExt_lo_1093 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1093 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1093 = {maskExt_hi_1093, maskExt_lo_1093};
  wire [15:0]         maskExt_lo_1094 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1094 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1094 = {maskExt_hi_1094, maskExt_lo_1094};
  wire [15:0]         maskExt_lo_1095 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1095 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1095 = {maskExt_hi_1095, maskExt_lo_1095};
  wire [15:0]         maskExt_lo_1096 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1096 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1096 = {maskExt_hi_1096, maskExt_lo_1096};
  wire [15:0]         maskExt_lo_1097 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1097 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1097 = {maskExt_hi_1097, maskExt_lo_1097};
  wire [15:0]         maskExt_lo_1098 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1098 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1098 = {maskExt_hi_1098, maskExt_lo_1098};
  wire [15:0]         maskExt_lo_1099 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1099 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1099 = {maskExt_hi_1099, maskExt_lo_1099};
  wire [15:0]         maskExt_lo_1100 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1100 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1100 = {maskExt_hi_1100, maskExt_lo_1100};
  wire [15:0]         maskExt_lo_1101 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1101 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1101 = {maskExt_hi_1101, maskExt_lo_1101};
  wire [15:0]         maskExt_lo_1102 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1102 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1102 = {maskExt_hi_1102, maskExt_lo_1102};
  wire [15:0]         maskExt_lo_1103 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1103 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1103 = {maskExt_hi_1103, maskExt_lo_1103};
  wire [15:0]         maskExt_lo_1104 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1104 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1104 = {maskExt_hi_1104, maskExt_lo_1104};
  wire [15:0]         maskExt_lo_1105 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1105 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1105 = {maskExt_hi_1105, maskExt_lo_1105};
  wire [15:0]         maskExt_lo_1106 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1106 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1106 = {maskExt_hi_1106, maskExt_lo_1106};
  wire [15:0]         maskExt_lo_1107 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1107 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1107 = {maskExt_hi_1107, maskExt_lo_1107};
  wire [15:0]         maskExt_lo_1108 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1108 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1108 = {maskExt_hi_1108, maskExt_lo_1108};
  wire [15:0]         maskExt_lo_1109 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1109 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1109 = {maskExt_hi_1109, maskExt_lo_1109};
  wire [15:0]         maskExt_lo_1110 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1110 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1110 = {maskExt_hi_1110, maskExt_lo_1110};
  wire [15:0]         maskExt_lo_1111 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1111 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1111 = {maskExt_hi_1111, maskExt_lo_1111};
  wire [15:0]         maskExt_lo_1112 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1112 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1112 = {maskExt_hi_1112, maskExt_lo_1112};
  wire [15:0]         maskExt_lo_1113 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1113 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1113 = {maskExt_hi_1113, maskExt_lo_1113};
  wire [15:0]         maskExt_lo_1114 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1114 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1114 = {maskExt_hi_1114, maskExt_lo_1114};
  wire [15:0]         maskExt_lo_1115 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1115 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1115 = {maskExt_hi_1115, maskExt_lo_1115};
  wire [15:0]         maskExt_lo_1116 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1116 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1116 = {maskExt_hi_1116, maskExt_lo_1116};
  wire [15:0]         maskExt_lo_1117 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1117 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1117 = {maskExt_hi_1117, maskExt_lo_1117};
  wire [15:0]         maskExt_lo_1118 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1118 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1118 = {maskExt_hi_1118, maskExt_lo_1118};
  wire [15:0]         maskExt_lo_1119 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1119 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1119 = {maskExt_hi_1119, maskExt_lo_1119};
  wire [15:0]         maskExt_lo_1120 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1120 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1120 = {maskExt_hi_1120, maskExt_lo_1120};
  wire [15:0]         maskExt_lo_1121 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1121 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1121 = {maskExt_hi_1121, maskExt_lo_1121};
  wire [15:0]         maskExt_lo_1122 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1122 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1122 = {maskExt_hi_1122, maskExt_lo_1122};
  wire [15:0]         maskExt_lo_1123 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1123 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1123 = {maskExt_hi_1123, maskExt_lo_1123};
  wire [15:0]         maskExt_lo_1124 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1124 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1124 = {maskExt_hi_1124, maskExt_lo_1124};
  wire [15:0]         maskExt_lo_1125 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1125 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1125 = {maskExt_hi_1125, maskExt_lo_1125};
  wire [15:0]         maskExt_lo_1126 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1126 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1126 = {maskExt_hi_1126, maskExt_lo_1126};
  wire [15:0]         maskExt_lo_1127 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1127 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1127 = {maskExt_hi_1127, maskExt_lo_1127};
  wire [15:0]         maskExt_lo_1128 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1128 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1128 = {maskExt_hi_1128, maskExt_lo_1128};
  wire [15:0]         maskExt_lo_1129 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1129 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1129 = {maskExt_hi_1129, maskExt_lo_1129};
  wire [15:0]         maskExt_lo_1130 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1130 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1130 = {maskExt_hi_1130, maskExt_lo_1130};
  wire [15:0]         maskExt_lo_1131 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1131 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1131 = {maskExt_hi_1131, maskExt_lo_1131};
  wire [15:0]         maskExt_lo_1132 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1132 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1132 = {maskExt_hi_1132, maskExt_lo_1132};
  wire [15:0]         maskExt_lo_1133 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1133 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1133 = {maskExt_hi_1133, maskExt_lo_1133};
  wire [15:0]         maskExt_lo_1134 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1134 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1134 = {maskExt_hi_1134, maskExt_lo_1134};
  wire [15:0]         maskExt_lo_1135 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1135 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1135 = {maskExt_hi_1135, maskExt_lo_1135};
  wire [15:0]         maskExt_lo_1136 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1136 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1136 = {maskExt_hi_1136, maskExt_lo_1136};
  wire [15:0]         maskExt_lo_1137 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1137 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1137 = {maskExt_hi_1137, maskExt_lo_1137};
  wire [15:0]         maskExt_lo_1138 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1138 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1138 = {maskExt_hi_1138, maskExt_lo_1138};
  wire [15:0]         maskExt_lo_1139 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1139 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1139 = {maskExt_hi_1139, maskExt_lo_1139};
  wire [15:0]         maskExt_lo_1140 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1140 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1140 = {maskExt_hi_1140, maskExt_lo_1140};
  wire [15:0]         maskExt_lo_1141 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1141 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1141 = {maskExt_hi_1141, maskExt_lo_1141};
  wire [15:0]         maskExt_lo_1142 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1142 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1142 = {maskExt_hi_1142, maskExt_lo_1142};
  wire [15:0]         maskExt_lo_1143 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1143 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1143 = {maskExt_hi_1143, maskExt_lo_1143};
  wire [15:0]         maskExt_lo_1144 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1144 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1144 = {maskExt_hi_1144, maskExt_lo_1144};
  wire [15:0]         maskExt_lo_1145 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1145 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1145 = {maskExt_hi_1145, maskExt_lo_1145};
  wire [15:0]         maskExt_lo_1146 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1146 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1146 = {maskExt_hi_1146, maskExt_lo_1146};
  wire [15:0]         maskExt_lo_1147 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1147 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1147 = {maskExt_hi_1147, maskExt_lo_1147};
  wire [15:0]         maskExt_lo_1148 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1148 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1148 = {maskExt_hi_1148, maskExt_lo_1148};
  wire [15:0]         maskExt_lo_1149 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1149 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1149 = {maskExt_hi_1149, maskExt_lo_1149};
  wire [15:0]         maskExt_lo_1150 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1150 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1150 = {maskExt_hi_1150, maskExt_lo_1150};
  wire [15:0]         maskExt_lo_1151 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1151 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1151 = {maskExt_hi_1151, maskExt_lo_1151};
  wire [15:0]         maskExt_lo_1152 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1152 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1152 = {maskExt_hi_1152, maskExt_lo_1152};
  wire [15:0]         maskExt_lo_1153 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1153 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1153 = {maskExt_hi_1153, maskExt_lo_1153};
  wire [15:0]         maskExt_lo_1154 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1154 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1154 = {maskExt_hi_1154, maskExt_lo_1154};
  wire [15:0]         maskExt_lo_1155 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1155 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1155 = {maskExt_hi_1155, maskExt_lo_1155};
  wire [15:0]         maskExt_lo_1156 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1156 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1156 = {maskExt_hi_1156, maskExt_lo_1156};
  wire [15:0]         maskExt_lo_1157 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1157 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1157 = {maskExt_hi_1157, maskExt_lo_1157};
  wire [15:0]         maskExt_lo_1158 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1158 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1158 = {maskExt_hi_1158, maskExt_lo_1158};
  wire [15:0]         maskExt_lo_1159 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1159 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1159 = {maskExt_hi_1159, maskExt_lo_1159};
  wire [15:0]         maskExt_lo_1160 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1160 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1160 = {maskExt_hi_1160, maskExt_lo_1160};
  wire [15:0]         maskExt_lo_1161 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1161 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1161 = {maskExt_hi_1161, maskExt_lo_1161};
  wire [15:0]         maskExt_lo_1162 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1162 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1162 = {maskExt_hi_1162, maskExt_lo_1162};
  wire [15:0]         maskExt_lo_1163 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1163 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1163 = {maskExt_hi_1163, maskExt_lo_1163};
  wire [15:0]         maskExt_lo_1164 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1164 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1164 = {maskExt_hi_1164, maskExt_lo_1164};
  wire [15:0]         maskExt_lo_1165 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1165 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1165 = {maskExt_hi_1165, maskExt_lo_1165};
  wire [15:0]         maskExt_lo_1166 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1166 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1166 = {maskExt_hi_1166, maskExt_lo_1166};
  wire [15:0]         maskExt_lo_1167 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1167 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1167 = {maskExt_hi_1167, maskExt_lo_1167};
  wire [15:0]         maskExt_lo_1168 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1168 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1168 = {maskExt_hi_1168, maskExt_lo_1168};
  wire [15:0]         maskExt_lo_1169 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1169 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1169 = {maskExt_hi_1169, maskExt_lo_1169};
  wire [15:0]         maskExt_lo_1170 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1170 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1170 = {maskExt_hi_1170, maskExt_lo_1170};
  wire [15:0]         maskExt_lo_1171 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1171 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1171 = {maskExt_hi_1171, maskExt_lo_1171};
  wire [15:0]         maskExt_lo_1172 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1172 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1172 = {maskExt_hi_1172, maskExt_lo_1172};
  wire [15:0]         maskExt_lo_1173 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1173 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1173 = {maskExt_hi_1173, maskExt_lo_1173};
  wire [15:0]         maskExt_lo_1174 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1174 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1174 = {maskExt_hi_1174, maskExt_lo_1174};
  wire [15:0]         maskExt_lo_1175 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1175 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1175 = {maskExt_hi_1175, maskExt_lo_1175};
  wire [15:0]         maskExt_lo_1176 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1176 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1176 = {maskExt_hi_1176, maskExt_lo_1176};
  wire [15:0]         maskExt_lo_1177 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1177 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1177 = {maskExt_hi_1177, maskExt_lo_1177};
  wire [15:0]         maskExt_lo_1178 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1178 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1178 = {maskExt_hi_1178, maskExt_lo_1178};
  wire [15:0]         maskExt_lo_1179 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1179 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1179 = {maskExt_hi_1179, maskExt_lo_1179};
  wire [15:0]         maskExt_lo_1180 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1180 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1180 = {maskExt_hi_1180, maskExt_lo_1180};
  wire [15:0]         maskExt_lo_1181 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1181 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1181 = {maskExt_hi_1181, maskExt_lo_1181};
  wire [15:0]         maskExt_lo_1182 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1182 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1182 = {maskExt_hi_1182, maskExt_lo_1182};
  wire [15:0]         maskExt_lo_1183 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1183 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1183 = {maskExt_hi_1183, maskExt_lo_1183};
  wire [15:0]         maskExt_lo_1184 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1184 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1184 = {maskExt_hi_1184, maskExt_lo_1184};
  wire [15:0]         maskExt_lo_1185 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1185 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1185 = {maskExt_hi_1185, maskExt_lo_1185};
  wire [15:0]         maskExt_lo_1186 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1186 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1186 = {maskExt_hi_1186, maskExt_lo_1186};
  wire [15:0]         maskExt_lo_1187 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1187 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1187 = {maskExt_hi_1187, maskExt_lo_1187};
  wire [15:0]         maskExt_lo_1188 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1188 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1188 = {maskExt_hi_1188, maskExt_lo_1188};
  wire [15:0]         maskExt_lo_1189 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1189 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1189 = {maskExt_hi_1189, maskExt_lo_1189};
  wire [15:0]         maskExt_lo_1190 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1190 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1190 = {maskExt_hi_1190, maskExt_lo_1190};
  wire [15:0]         maskExt_lo_1191 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1191 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1191 = {maskExt_hi_1191, maskExt_lo_1191};
  wire [15:0]         maskExt_lo_1192 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1192 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1192 = {maskExt_hi_1192, maskExt_lo_1192};
  wire [15:0]         maskExt_lo_1193 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1193 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1193 = {maskExt_hi_1193, maskExt_lo_1193};
  wire [15:0]         maskExt_lo_1194 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1194 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1194 = {maskExt_hi_1194, maskExt_lo_1194};
  wire [15:0]         maskExt_lo_1195 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1195 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1195 = {maskExt_hi_1195, maskExt_lo_1195};
  wire [15:0]         maskExt_lo_1196 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1196 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1196 = {maskExt_hi_1196, maskExt_lo_1196};
  wire [15:0]         maskExt_lo_1197 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1197 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1197 = {maskExt_hi_1197, maskExt_lo_1197};
  wire [15:0]         maskExt_lo_1198 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1198 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1198 = {maskExt_hi_1198, maskExt_lo_1198};
  wire [15:0]         maskExt_lo_1199 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1199 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1199 = {maskExt_hi_1199, maskExt_lo_1199};
  wire [15:0]         maskExt_lo_1200 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1200 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1200 = {maskExt_hi_1200, maskExt_lo_1200};
  wire [15:0]         maskExt_lo_1201 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1201 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1201 = {maskExt_hi_1201, maskExt_lo_1201};
  wire [15:0]         maskExt_lo_1202 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1202 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1202 = {maskExt_hi_1202, maskExt_lo_1202};
  wire [15:0]         maskExt_lo_1203 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1203 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1203 = {maskExt_hi_1203, maskExt_lo_1203};
  wire [15:0]         maskExt_lo_1204 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1204 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1204 = {maskExt_hi_1204, maskExt_lo_1204};
  wire [15:0]         maskExt_lo_1205 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1205 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1205 = {maskExt_hi_1205, maskExt_lo_1205};
  wire [15:0]         maskExt_lo_1206 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1206 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1206 = {maskExt_hi_1206, maskExt_lo_1206};
  wire [15:0]         maskExt_lo_1207 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1207 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1207 = {maskExt_hi_1207, maskExt_lo_1207};
  wire [15:0]         maskExt_lo_1208 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1208 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1208 = {maskExt_hi_1208, maskExt_lo_1208};
  wire [15:0]         maskExt_lo_1209 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1209 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1209 = {maskExt_hi_1209, maskExt_lo_1209};
  wire [15:0]         maskExt_lo_1210 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1210 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1210 = {maskExt_hi_1210, maskExt_lo_1210};
  wire [15:0]         maskExt_lo_1211 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1211 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1211 = {maskExt_hi_1211, maskExt_lo_1211};
  wire [15:0]         maskExt_lo_1212 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1212 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1212 = {maskExt_hi_1212, maskExt_lo_1212};
  wire [15:0]         maskExt_lo_1213 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1213 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1213 = {maskExt_hi_1213, maskExt_lo_1213};
  wire [15:0]         maskExt_lo_1214 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1214 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1214 = {maskExt_hi_1214, maskExt_lo_1214};
  wire [15:0]         maskExt_lo_1215 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1215 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1215 = {maskExt_hi_1215, maskExt_lo_1215};
  wire [15:0]         maskExt_lo_1216 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1216 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1216 = {maskExt_hi_1216, maskExt_lo_1216};
  wire [15:0]         maskExt_lo_1217 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1217 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1217 = {maskExt_hi_1217, maskExt_lo_1217};
  wire [15:0]         maskExt_lo_1218 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1218 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1218 = {maskExt_hi_1218, maskExt_lo_1218};
  wire [15:0]         maskExt_lo_1219 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1219 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1219 = {maskExt_hi_1219, maskExt_lo_1219};
  wire [15:0]         maskExt_lo_1220 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1220 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1220 = {maskExt_hi_1220, maskExt_lo_1220};
  wire [15:0]         maskExt_lo_1221 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1221 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1221 = {maskExt_hi_1221, maskExt_lo_1221};
  wire [15:0]         maskExt_lo_1222 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1222 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1222 = {maskExt_hi_1222, maskExt_lo_1222};
  wire [15:0]         maskExt_lo_1223 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1223 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1223 = {maskExt_hi_1223, maskExt_lo_1223};
  wire [15:0]         maskExt_lo_1224 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1224 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1224 = {maskExt_hi_1224, maskExt_lo_1224};
  wire [15:0]         maskExt_lo_1225 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1225 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1225 = {maskExt_hi_1225, maskExt_lo_1225};
  wire [15:0]         maskExt_lo_1226 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1226 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1226 = {maskExt_hi_1226, maskExt_lo_1226};
  wire [15:0]         maskExt_lo_1227 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1227 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1227 = {maskExt_hi_1227, maskExt_lo_1227};
  wire [15:0]         maskExt_lo_1228 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1228 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1228 = {maskExt_hi_1228, maskExt_lo_1228};
  wire [15:0]         maskExt_lo_1229 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1229 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1229 = {maskExt_hi_1229, maskExt_lo_1229};
  wire [15:0]         maskExt_lo_1230 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1230 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1230 = {maskExt_hi_1230, maskExt_lo_1230};
  wire [15:0]         maskExt_lo_1231 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1231 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1231 = {maskExt_hi_1231, maskExt_lo_1231};
  wire [15:0]         maskExt_lo_1232 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1232 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1232 = {maskExt_hi_1232, maskExt_lo_1232};
  wire [15:0]         maskExt_lo_1233 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1233 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1233 = {maskExt_hi_1233, maskExt_lo_1233};
  wire [15:0]         maskExt_lo_1234 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1234 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1234 = {maskExt_hi_1234, maskExt_lo_1234};
  wire [15:0]         maskExt_lo_1235 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1235 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1235 = {maskExt_hi_1235, maskExt_lo_1235};
  wire [15:0]         maskExt_lo_1236 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1236 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1236 = {maskExt_hi_1236, maskExt_lo_1236};
  wire [15:0]         maskExt_lo_1237 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1237 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1237 = {maskExt_hi_1237, maskExt_lo_1237};
  wire [15:0]         maskExt_lo_1238 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1238 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1238 = {maskExt_hi_1238, maskExt_lo_1238};
  wire [15:0]         maskExt_lo_1239 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1239 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1239 = {maskExt_hi_1239, maskExt_lo_1239};
  wire [15:0]         maskExt_lo_1240 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1240 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1240 = {maskExt_hi_1240, maskExt_lo_1240};
  wire [15:0]         maskExt_lo_1241 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1241 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1241 = {maskExt_hi_1241, maskExt_lo_1241};
  wire [15:0]         maskExt_lo_1242 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1242 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1242 = {maskExt_hi_1242, maskExt_lo_1242};
  wire [15:0]         maskExt_lo_1243 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1243 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1243 = {maskExt_hi_1243, maskExt_lo_1243};
  wire [15:0]         maskExt_lo_1244 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1244 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1244 = {maskExt_hi_1244, maskExt_lo_1244};
  wire [15:0]         maskExt_lo_1245 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1245 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1245 = {maskExt_hi_1245, maskExt_lo_1245};
  wire [15:0]         maskExt_lo_1246 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1246 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1246 = {maskExt_hi_1246, maskExt_lo_1246};
  wire [15:0]         maskExt_lo_1247 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1247 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1247 = {maskExt_hi_1247, maskExt_lo_1247};
  wire [15:0]         maskExt_lo_1248 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1248 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1248 = {maskExt_hi_1248, maskExt_lo_1248};
  wire [15:0]         maskExt_lo_1249 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1249 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1249 = {maskExt_hi_1249, maskExt_lo_1249};
  wire [15:0]         maskExt_lo_1250 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1250 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1250 = {maskExt_hi_1250, maskExt_lo_1250};
  wire [15:0]         maskExt_lo_1251 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1251 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1251 = {maskExt_hi_1251, maskExt_lo_1251};
  wire [15:0]         maskExt_lo_1252 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1252 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1252 = {maskExt_hi_1252, maskExt_lo_1252};
  wire [15:0]         maskExt_lo_1253 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1253 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1253 = {maskExt_hi_1253, maskExt_lo_1253};
  wire [15:0]         maskExt_lo_1254 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1254 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1254 = {maskExt_hi_1254, maskExt_lo_1254};
  wire [15:0]         maskExt_lo_1255 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1255 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1255 = {maskExt_hi_1255, maskExt_lo_1255};
  wire [15:0]         maskExt_lo_1256 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1256 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1256 = {maskExt_hi_1256, maskExt_lo_1256};
  wire [15:0]         maskExt_lo_1257 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1257 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1257 = {maskExt_hi_1257, maskExt_lo_1257};
  wire [15:0]         maskExt_lo_1258 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1258 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1258 = {maskExt_hi_1258, maskExt_lo_1258};
  wire [15:0]         maskExt_lo_1259 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1259 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1259 = {maskExt_hi_1259, maskExt_lo_1259};
  wire [15:0]         maskExt_lo_1260 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1260 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1260 = {maskExt_hi_1260, maskExt_lo_1260};
  wire [15:0]         maskExt_lo_1261 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1261 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1261 = {maskExt_hi_1261, maskExt_lo_1261};
  wire [15:0]         maskExt_lo_1262 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1262 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1262 = {maskExt_hi_1262, maskExt_lo_1262};
  wire [15:0]         maskExt_lo_1263 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1263 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1263 = {maskExt_hi_1263, maskExt_lo_1263};
  wire [15:0]         maskExt_lo_1264 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1264 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1264 = {maskExt_hi_1264, maskExt_lo_1264};
  wire [15:0]         maskExt_lo_1265 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1265 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1265 = {maskExt_hi_1265, maskExt_lo_1265};
  wire [15:0]         maskExt_lo_1266 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1266 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1266 = {maskExt_hi_1266, maskExt_lo_1266};
  wire [15:0]         maskExt_lo_1267 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1267 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1267 = {maskExt_hi_1267, maskExt_lo_1267};
  wire [15:0]         maskExt_lo_1268 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1268 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1268 = {maskExt_hi_1268, maskExt_lo_1268};
  wire [15:0]         maskExt_lo_1269 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1269 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1269 = {maskExt_hi_1269, maskExt_lo_1269};
  wire [15:0]         maskExt_lo_1270 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1270 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1270 = {maskExt_hi_1270, maskExt_lo_1270};
  wire [15:0]         maskExt_lo_1271 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1271 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1271 = {maskExt_hi_1271, maskExt_lo_1271};
  wire [15:0]         maskExt_lo_1272 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1272 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1272 = {maskExt_hi_1272, maskExt_lo_1272};
  wire [15:0]         maskExt_lo_1273 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1273 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1273 = {maskExt_hi_1273, maskExt_lo_1273};
  wire [15:0]         maskExt_lo_1274 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1274 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1274 = {maskExt_hi_1274, maskExt_lo_1274};
  wire [15:0]         maskExt_lo_1275 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1275 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1275 = {maskExt_hi_1275, maskExt_lo_1275};
  wire [15:0]         maskExt_lo_1276 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1276 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1276 = {maskExt_hi_1276, maskExt_lo_1276};
  wire [15:0]         maskExt_lo_1277 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1277 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1277 = {maskExt_hi_1277, maskExt_lo_1277};
  wire [15:0]         maskExt_lo_1278 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1278 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1278 = {maskExt_hi_1278, maskExt_lo_1278};
  wire [15:0]         maskExt_lo_1279 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1279 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1279 = {maskExt_hi_1279, maskExt_lo_1279};
  wire [15:0]         maskExt_lo_1280 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1280 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1280 = {maskExt_hi_1280, maskExt_lo_1280};
  wire [15:0]         maskExt_lo_1281 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1281 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1281 = {maskExt_hi_1281, maskExt_lo_1281};
  wire [15:0]         maskExt_lo_1282 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1282 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1282 = {maskExt_hi_1282, maskExt_lo_1282};
  wire [15:0]         maskExt_lo_1283 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1283 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1283 = {maskExt_hi_1283, maskExt_lo_1283};
  wire [15:0]         maskExt_lo_1284 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1284 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1284 = {maskExt_hi_1284, maskExt_lo_1284};
  wire [15:0]         maskExt_lo_1285 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1285 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1285 = {maskExt_hi_1285, maskExt_lo_1285};
  wire [15:0]         maskExt_lo_1286 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1286 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1286 = {maskExt_hi_1286, maskExt_lo_1286};
  wire [15:0]         maskExt_lo_1287 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1287 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1287 = {maskExt_hi_1287, maskExt_lo_1287};
  wire [15:0]         maskExt_lo_1288 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1288 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1288 = {maskExt_hi_1288, maskExt_lo_1288};
  wire [15:0]         maskExt_lo_1289 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1289 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1289 = {maskExt_hi_1289, maskExt_lo_1289};
  wire [15:0]         maskExt_lo_1290 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1290 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1290 = {maskExt_hi_1290, maskExt_lo_1290};
  wire [15:0]         maskExt_lo_1291 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1291 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1291 = {maskExt_hi_1291, maskExt_lo_1291};
  wire [15:0]         maskExt_lo_1292 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1292 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1292 = {maskExt_hi_1292, maskExt_lo_1292};
  wire [15:0]         maskExt_lo_1293 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1293 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1293 = {maskExt_hi_1293, maskExt_lo_1293};
  wire [15:0]         maskExt_lo_1294 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1294 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1294 = {maskExt_hi_1294, maskExt_lo_1294};
  wire [15:0]         maskExt_lo_1295 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1295 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1295 = {maskExt_hi_1295, maskExt_lo_1295};
  wire [15:0]         maskExt_lo_1296 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1296 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1296 = {maskExt_hi_1296, maskExt_lo_1296};
  wire [15:0]         maskExt_lo_1297 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1297 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1297 = {maskExt_hi_1297, maskExt_lo_1297};
  wire [15:0]         maskExt_lo_1298 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1298 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1298 = {maskExt_hi_1298, maskExt_lo_1298};
  wire [15:0]         maskExt_lo_1299 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1299 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1299 = {maskExt_hi_1299, maskExt_lo_1299};
  wire [15:0]         maskExt_lo_1300 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1300 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1300 = {maskExt_hi_1300, maskExt_lo_1300};
  wire [15:0]         maskExt_lo_1301 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1301 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1301 = {maskExt_hi_1301, maskExt_lo_1301};
  wire [15:0]         maskExt_lo_1302 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1302 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1302 = {maskExt_hi_1302, maskExt_lo_1302};
  wire [15:0]         maskExt_lo_1303 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1303 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1303 = {maskExt_hi_1303, maskExt_lo_1303};
  wire [15:0]         maskExt_lo_1304 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1304 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1304 = {maskExt_hi_1304, maskExt_lo_1304};
  wire [15:0]         maskExt_lo_1305 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1305 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1305 = {maskExt_hi_1305, maskExt_lo_1305};
  wire [15:0]         maskExt_lo_1306 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1306 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1306 = {maskExt_hi_1306, maskExt_lo_1306};
  wire [15:0]         maskExt_lo_1307 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1307 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1307 = {maskExt_hi_1307, maskExt_lo_1307};
  wire [15:0]         maskExt_lo_1308 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1308 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1308 = {maskExt_hi_1308, maskExt_lo_1308};
  wire [15:0]         maskExt_lo_1309 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1309 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1309 = {maskExt_hi_1309, maskExt_lo_1309};
  wire [15:0]         maskExt_lo_1310 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1310 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1310 = {maskExt_hi_1310, maskExt_lo_1310};
  wire [15:0]         maskExt_lo_1311 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1311 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1311 = {maskExt_hi_1311, maskExt_lo_1311};
  wire [15:0]         maskExt_lo_1312 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1312 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1312 = {maskExt_hi_1312, maskExt_lo_1312};
  wire [15:0]         maskExt_lo_1313 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1313 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1313 = {maskExt_hi_1313, maskExt_lo_1313};
  wire [15:0]         maskExt_lo_1314 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1314 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1314 = {maskExt_hi_1314, maskExt_lo_1314};
  wire [15:0]         maskExt_lo_1315 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1315 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1315 = {maskExt_hi_1315, maskExt_lo_1315};
  wire [15:0]         maskExt_lo_1316 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1316 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1316 = {maskExt_hi_1316, maskExt_lo_1316};
  wire [15:0]         maskExt_lo_1317 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1317 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1317 = {maskExt_hi_1317, maskExt_lo_1317};
  wire [15:0]         maskExt_lo_1318 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1318 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1318 = {maskExt_hi_1318, maskExt_lo_1318};
  wire [15:0]         maskExt_lo_1319 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1319 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1319 = {maskExt_hi_1319, maskExt_lo_1319};
  wire [15:0]         maskExt_lo_1320 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1320 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1320 = {maskExt_hi_1320, maskExt_lo_1320};
  wire [15:0]         maskExt_lo_1321 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1321 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1321 = {maskExt_hi_1321, maskExt_lo_1321};
  wire [15:0]         maskExt_lo_1322 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1322 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1322 = {maskExt_hi_1322, maskExt_lo_1322};
  wire [15:0]         maskExt_lo_1323 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1323 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1323 = {maskExt_hi_1323, maskExt_lo_1323};
  wire [15:0]         maskExt_lo_1324 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1324 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1324 = {maskExt_hi_1324, maskExt_lo_1324};
  wire [15:0]         maskExt_lo_1325 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1325 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1325 = {maskExt_hi_1325, maskExt_lo_1325};
  wire [15:0]         maskExt_lo_1326 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1326 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1326 = {maskExt_hi_1326, maskExt_lo_1326};
  wire [15:0]         maskExt_lo_1327 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1327 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1327 = {maskExt_hi_1327, maskExt_lo_1327};
  wire [15:0]         maskExt_lo_1328 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1328 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1328 = {maskExt_hi_1328, maskExt_lo_1328};
  wire [15:0]         maskExt_lo_1329 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1329 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1329 = {maskExt_hi_1329, maskExt_lo_1329};
  wire [15:0]         maskExt_lo_1330 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1330 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1330 = {maskExt_hi_1330, maskExt_lo_1330};
  wire [15:0]         maskExt_lo_1331 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1331 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1331 = {maskExt_hi_1331, maskExt_lo_1331};
  wire [15:0]         maskExt_lo_1332 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1332 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1332 = {maskExt_hi_1332, maskExt_lo_1332};
  wire [15:0]         maskExt_lo_1333 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1333 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1333 = {maskExt_hi_1333, maskExt_lo_1333};
  wire [15:0]         maskExt_lo_1334 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1334 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1334 = {maskExt_hi_1334, maskExt_lo_1334};
  wire [15:0]         maskExt_lo_1335 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1335 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1335 = {maskExt_hi_1335, maskExt_lo_1335};
  wire [15:0]         maskExt_lo_1336 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1336 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1336 = {maskExt_hi_1336, maskExt_lo_1336};
  wire [15:0]         maskExt_lo_1337 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1337 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1337 = {maskExt_hi_1337, maskExt_lo_1337};
  wire [15:0]         maskExt_lo_1338 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1338 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1338 = {maskExt_hi_1338, maskExt_lo_1338};
  wire [15:0]         maskExt_lo_1339 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1339 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1339 = {maskExt_hi_1339, maskExt_lo_1339};
  wire [15:0]         maskExt_lo_1340 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1340 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1340 = {maskExt_hi_1340, maskExt_lo_1340};
  wire [15:0]         maskExt_lo_1341 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1341 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1341 = {maskExt_hi_1341, maskExt_lo_1341};
  wire [15:0]         maskExt_lo_1342 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1342 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1342 = {maskExt_hi_1342, maskExt_lo_1342};
  wire [15:0]         maskExt_lo_1343 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1343 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1343 = {maskExt_hi_1343, maskExt_lo_1343};
  wire [15:0]         maskExt_lo_1344 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1344 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1344 = {maskExt_hi_1344, maskExt_lo_1344};
  wire [15:0]         maskExt_lo_1345 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1345 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1345 = {maskExt_hi_1345, maskExt_lo_1345};
  wire [15:0]         maskExt_lo_1346 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1346 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1346 = {maskExt_hi_1346, maskExt_lo_1346};
  wire [15:0]         maskExt_lo_1347 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1347 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1347 = {maskExt_hi_1347, maskExt_lo_1347};
  wire [15:0]         maskExt_lo_1348 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1348 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1348 = {maskExt_hi_1348, maskExt_lo_1348};
  wire [15:0]         maskExt_lo_1349 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1349 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1349 = {maskExt_hi_1349, maskExt_lo_1349};
  wire [15:0]         maskExt_lo_1350 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1350 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1350 = {maskExt_hi_1350, maskExt_lo_1350};
  wire [15:0]         maskExt_lo_1351 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1351 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1351 = {maskExt_hi_1351, maskExt_lo_1351};
  wire [15:0]         maskExt_lo_1352 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1352 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1352 = {maskExt_hi_1352, maskExt_lo_1352};
  wire [15:0]         maskExt_lo_1353 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1353 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1353 = {maskExt_hi_1353, maskExt_lo_1353};
  wire [15:0]         maskExt_lo_1354 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1354 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1354 = {maskExt_hi_1354, maskExt_lo_1354};
  wire [15:0]         maskExt_lo_1355 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1355 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1355 = {maskExt_hi_1355, maskExt_lo_1355};
  wire [15:0]         maskExt_lo_1356 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1356 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1356 = {maskExt_hi_1356, maskExt_lo_1356};
  wire [15:0]         maskExt_lo_1357 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1357 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1357 = {maskExt_hi_1357, maskExt_lo_1357};
  wire [15:0]         maskExt_lo_1358 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1358 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1358 = {maskExt_hi_1358, maskExt_lo_1358};
  wire [15:0]         maskExt_lo_1359 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1359 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1359 = {maskExt_hi_1359, maskExt_lo_1359};
  wire [15:0]         maskExt_lo_1360 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1360 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1360 = {maskExt_hi_1360, maskExt_lo_1360};
  wire [15:0]         maskExt_lo_1361 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1361 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1361 = {maskExt_hi_1361, maskExt_lo_1361};
  wire [15:0]         maskExt_lo_1362 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1362 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1362 = {maskExt_hi_1362, maskExt_lo_1362};
  wire [15:0]         maskExt_lo_1363 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1363 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1363 = {maskExt_hi_1363, maskExt_lo_1363};
  wire [15:0]         maskExt_lo_1364 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1364 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1364 = {maskExt_hi_1364, maskExt_lo_1364};
  wire [15:0]         maskExt_lo_1365 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1365 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1365 = {maskExt_hi_1365, maskExt_lo_1365};
  wire [15:0]         maskExt_lo_1366 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1366 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1366 = {maskExt_hi_1366, maskExt_lo_1366};
  wire [15:0]         maskExt_lo_1367 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1367 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1367 = {maskExt_hi_1367, maskExt_lo_1367};
  wire [15:0]         maskExt_lo_1368 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1368 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1368 = {maskExt_hi_1368, maskExt_lo_1368};
  wire [15:0]         maskExt_lo_1369 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1369 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1369 = {maskExt_hi_1369, maskExt_lo_1369};
  wire [15:0]         maskExt_lo_1370 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1370 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1370 = {maskExt_hi_1370, maskExt_lo_1370};
  wire [15:0]         maskExt_lo_1371 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1371 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1371 = {maskExt_hi_1371, maskExt_lo_1371};
  wire [15:0]         maskExt_lo_1372 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1372 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1372 = {maskExt_hi_1372, maskExt_lo_1372};
  wire [15:0]         maskExt_lo_1373 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1373 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1373 = {maskExt_hi_1373, maskExt_lo_1373};
  wire [15:0]         maskExt_lo_1374 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1374 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1374 = {maskExt_hi_1374, maskExt_lo_1374};
  wire [15:0]         maskExt_lo_1375 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1375 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1375 = {maskExt_hi_1375, maskExt_lo_1375};
  wire [15:0]         maskExt_lo_1376 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1376 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1376 = {maskExt_hi_1376, maskExt_lo_1376};
  wire [15:0]         maskExt_lo_1377 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1377 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1377 = {maskExt_hi_1377, maskExt_lo_1377};
  wire [15:0]         maskExt_lo_1378 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1378 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1378 = {maskExt_hi_1378, maskExt_lo_1378};
  wire [15:0]         maskExt_lo_1379 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1379 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1379 = {maskExt_hi_1379, maskExt_lo_1379};
  wire [15:0]         maskExt_lo_1380 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1380 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1380 = {maskExt_hi_1380, maskExt_lo_1380};
  wire [15:0]         maskExt_lo_1381 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1381 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1381 = {maskExt_hi_1381, maskExt_lo_1381};
  wire [15:0]         maskExt_lo_1382 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1382 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1382 = {maskExt_hi_1382, maskExt_lo_1382};
  wire [15:0]         maskExt_lo_1383 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1383 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1383 = {maskExt_hi_1383, maskExt_lo_1383};
  wire [15:0]         maskExt_lo_1384 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1384 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1384 = {maskExt_hi_1384, maskExt_lo_1384};
  wire [15:0]         maskExt_lo_1385 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1385 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1385 = {maskExt_hi_1385, maskExt_lo_1385};
  wire [15:0]         maskExt_lo_1386 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1386 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1386 = {maskExt_hi_1386, maskExt_lo_1386};
  wire [15:0]         maskExt_lo_1387 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1387 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1387 = {maskExt_hi_1387, maskExt_lo_1387};
  wire [15:0]         maskExt_lo_1388 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1388 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1388 = {maskExt_hi_1388, maskExt_lo_1388};
  wire [15:0]         maskExt_lo_1389 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1389 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1389 = {maskExt_hi_1389, maskExt_lo_1389};
  wire [15:0]         maskExt_lo_1390 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1390 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1390 = {maskExt_hi_1390, maskExt_lo_1390};
  wire [15:0]         maskExt_lo_1391 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1391 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1391 = {maskExt_hi_1391, maskExt_lo_1391};
  wire [15:0]         maskExt_lo_1392 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1392 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1392 = {maskExt_hi_1392, maskExt_lo_1392};
  wire [15:0]         maskExt_lo_1393 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1393 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1393 = {maskExt_hi_1393, maskExt_lo_1393};
  wire [15:0]         maskExt_lo_1394 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1394 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1394 = {maskExt_hi_1394, maskExt_lo_1394};
  wire [15:0]         maskExt_lo_1395 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1395 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1395 = {maskExt_hi_1395, maskExt_lo_1395};
  wire [15:0]         maskExt_lo_1396 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1396 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1396 = {maskExt_hi_1396, maskExt_lo_1396};
  wire [15:0]         maskExt_lo_1397 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1397 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1397 = {maskExt_hi_1397, maskExt_lo_1397};
  wire [15:0]         maskExt_lo_1398 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1398 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1398 = {maskExt_hi_1398, maskExt_lo_1398};
  wire [15:0]         maskExt_lo_1399 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1399 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1399 = {maskExt_hi_1399, maskExt_lo_1399};
  wire [15:0]         maskExt_lo_1400 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1400 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1400 = {maskExt_hi_1400, maskExt_lo_1400};
  wire [15:0]         maskExt_lo_1401 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1401 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1401 = {maskExt_hi_1401, maskExt_lo_1401};
  wire [15:0]         maskExt_lo_1402 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1402 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1402 = {maskExt_hi_1402, maskExt_lo_1402};
  wire [15:0]         maskExt_lo_1403 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1403 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1403 = {maskExt_hi_1403, maskExt_lo_1403};
  wire [15:0]         maskExt_lo_1404 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1404 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1404 = {maskExt_hi_1404, maskExt_lo_1404};
  wire [15:0]         maskExt_lo_1405 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1405 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1405 = {maskExt_hi_1405, maskExt_lo_1405};
  wire [15:0]         maskExt_lo_1406 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1406 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1406 = {maskExt_hi_1406, maskExt_lo_1406};
  wire [15:0]         maskExt_lo_1407 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1407 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1407 = {maskExt_hi_1407, maskExt_lo_1407};
  wire [15:0]         maskExt_lo_1408 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1408 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1408 = {maskExt_hi_1408, maskExt_lo_1408};
  wire [15:0]         maskExt_lo_1409 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1409 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1409 = {maskExt_hi_1409, maskExt_lo_1409};
  wire [15:0]         maskExt_lo_1410 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1410 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1410 = {maskExt_hi_1410, maskExt_lo_1410};
  wire [15:0]         maskExt_lo_1411 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1411 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1411 = {maskExt_hi_1411, maskExt_lo_1411};
  wire [15:0]         maskExt_lo_1412 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1412 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1412 = {maskExt_hi_1412, maskExt_lo_1412};
  wire [15:0]         maskExt_lo_1413 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1413 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1413 = {maskExt_hi_1413, maskExt_lo_1413};
  wire [15:0]         maskExt_lo_1414 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1414 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1414 = {maskExt_hi_1414, maskExt_lo_1414};
  wire [15:0]         maskExt_lo_1415 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1415 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1415 = {maskExt_hi_1415, maskExt_lo_1415};
  wire [15:0]         maskExt_lo_1416 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1416 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1416 = {maskExt_hi_1416, maskExt_lo_1416};
  wire [15:0]         maskExt_lo_1417 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1417 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1417 = {maskExt_hi_1417, maskExt_lo_1417};
  wire [15:0]         maskExt_lo_1418 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1418 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1418 = {maskExt_hi_1418, maskExt_lo_1418};
  wire [15:0]         maskExt_lo_1419 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1419 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1419 = {maskExt_hi_1419, maskExt_lo_1419};
  wire [15:0]         maskExt_lo_1420 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1420 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1420 = {maskExt_hi_1420, maskExt_lo_1420};
  wire [15:0]         maskExt_lo_1421 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1421 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1421 = {maskExt_hi_1421, maskExt_lo_1421};
  wire [15:0]         maskExt_lo_1422 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1422 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1422 = {maskExt_hi_1422, maskExt_lo_1422};
  wire [15:0]         maskExt_lo_1423 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1423 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1423 = {maskExt_hi_1423, maskExt_lo_1423};
  wire [15:0]         maskExt_lo_1424 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1424 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1424 = {maskExt_hi_1424, maskExt_lo_1424};
  wire [15:0]         maskExt_lo_1425 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1425 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1425 = {maskExt_hi_1425, maskExt_lo_1425};
  wire [15:0]         maskExt_lo_1426 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1426 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1426 = {maskExt_hi_1426, maskExt_lo_1426};
  wire [15:0]         maskExt_lo_1427 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1427 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1427 = {maskExt_hi_1427, maskExt_lo_1427};
  wire [15:0]         maskExt_lo_1428 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1428 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1428 = {maskExt_hi_1428, maskExt_lo_1428};
  wire [15:0]         maskExt_lo_1429 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1429 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1429 = {maskExt_hi_1429, maskExt_lo_1429};
  wire [15:0]         maskExt_lo_1430 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1430 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1430 = {maskExt_hi_1430, maskExt_lo_1430};
  wire [15:0]         maskExt_lo_1431 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1431 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1431 = {maskExt_hi_1431, maskExt_lo_1431};
  wire [15:0]         maskExt_lo_1432 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1432 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1432 = {maskExt_hi_1432, maskExt_lo_1432};
  wire [15:0]         maskExt_lo_1433 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1433 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1433 = {maskExt_hi_1433, maskExt_lo_1433};
  wire [15:0]         maskExt_lo_1434 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1434 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1434 = {maskExt_hi_1434, maskExt_lo_1434};
  wire [15:0]         maskExt_lo_1435 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1435 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1435 = {maskExt_hi_1435, maskExt_lo_1435};
  wire [15:0]         maskExt_lo_1436 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1436 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1436 = {maskExt_hi_1436, maskExt_lo_1436};
  wire [15:0]         maskExt_lo_1437 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1437 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1437 = {maskExt_hi_1437, maskExt_lo_1437};
  wire [15:0]         maskExt_lo_1438 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1438 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1438 = {maskExt_hi_1438, maskExt_lo_1438};
  wire [15:0]         maskExt_lo_1439 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1439 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1439 = {maskExt_hi_1439, maskExt_lo_1439};
  wire [15:0]         maskExt_lo_1440 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1440 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1440 = {maskExt_hi_1440, maskExt_lo_1440};
  wire [15:0]         maskExt_lo_1441 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1441 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1441 = {maskExt_hi_1441, maskExt_lo_1441};
  wire [15:0]         maskExt_lo_1442 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1442 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1442 = {maskExt_hi_1442, maskExt_lo_1442};
  wire [15:0]         maskExt_lo_1443 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1443 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1443 = {maskExt_hi_1443, maskExt_lo_1443};
  wire [15:0]         maskExt_lo_1444 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1444 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1444 = {maskExt_hi_1444, maskExt_lo_1444};
  wire [15:0]         maskExt_lo_1445 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1445 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1445 = {maskExt_hi_1445, maskExt_lo_1445};
  wire [15:0]         maskExt_lo_1446 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1446 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1446 = {maskExt_hi_1446, maskExt_lo_1446};
  wire [15:0]         maskExt_lo_1447 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1447 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1447 = {maskExt_hi_1447, maskExt_lo_1447};
  wire [15:0]         maskExt_lo_1448 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1448 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1448 = {maskExt_hi_1448, maskExt_lo_1448};
  wire [15:0]         maskExt_lo_1449 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1449 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1449 = {maskExt_hi_1449, maskExt_lo_1449};
  wire [15:0]         maskExt_lo_1450 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1450 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1450 = {maskExt_hi_1450, maskExt_lo_1450};
  wire [15:0]         maskExt_lo_1451 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1451 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1451 = {maskExt_hi_1451, maskExt_lo_1451};
  wire [15:0]         maskExt_lo_1452 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1452 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1452 = {maskExt_hi_1452, maskExt_lo_1452};
  wire [15:0]         maskExt_lo_1453 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1453 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1453 = {maskExt_hi_1453, maskExt_lo_1453};
  wire [15:0]         maskExt_lo_1454 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1454 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1454 = {maskExt_hi_1454, maskExt_lo_1454};
  wire [15:0]         maskExt_lo_1455 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1455 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1455 = {maskExt_hi_1455, maskExt_lo_1455};
  wire [15:0]         maskExt_lo_1456 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1456 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1456 = {maskExt_hi_1456, maskExt_lo_1456};
  wire [15:0]         maskExt_lo_1457 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1457 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1457 = {maskExt_hi_1457, maskExt_lo_1457};
  wire [15:0]         maskExt_lo_1458 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1458 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1458 = {maskExt_hi_1458, maskExt_lo_1458};
  wire [15:0]         maskExt_lo_1459 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1459 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1459 = {maskExt_hi_1459, maskExt_lo_1459};
  wire [15:0]         maskExt_lo_1460 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1460 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1460 = {maskExt_hi_1460, maskExt_lo_1460};
  wire [15:0]         maskExt_lo_1461 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1461 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1461 = {maskExt_hi_1461, maskExt_lo_1461};
  wire [15:0]         maskExt_lo_1462 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1462 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1462 = {maskExt_hi_1462, maskExt_lo_1462};
  wire [15:0]         maskExt_lo_1463 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1463 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1463 = {maskExt_hi_1463, maskExt_lo_1463};
  wire [15:0]         maskExt_lo_1464 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1464 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1464 = {maskExt_hi_1464, maskExt_lo_1464};
  wire [15:0]         maskExt_lo_1465 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1465 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1465 = {maskExt_hi_1465, maskExt_lo_1465};
  wire [15:0]         maskExt_lo_1466 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1466 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1466 = {maskExt_hi_1466, maskExt_lo_1466};
  wire [15:0]         maskExt_lo_1467 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1467 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1467 = {maskExt_hi_1467, maskExt_lo_1467};
  wire [15:0]         maskExt_lo_1468 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1468 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1468 = {maskExt_hi_1468, maskExt_lo_1468};
  wire [15:0]         maskExt_lo_1469 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1469 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1469 = {maskExt_hi_1469, maskExt_lo_1469};
  wire [15:0]         maskExt_lo_1470 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1470 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1470 = {maskExt_hi_1470, maskExt_lo_1470};
  wire [15:0]         maskExt_lo_1471 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1471 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1471 = {maskExt_hi_1471, maskExt_lo_1471};
  wire [15:0]         maskExt_lo_1472 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1472 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1472 = {maskExt_hi_1472, maskExt_lo_1472};
  wire [15:0]         maskExt_lo_1473 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1473 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1473 = {maskExt_hi_1473, maskExt_lo_1473};
  wire [15:0]         maskExt_lo_1474 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1474 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1474 = {maskExt_hi_1474, maskExt_lo_1474};
  wire [15:0]         maskExt_lo_1475 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1475 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1475 = {maskExt_hi_1475, maskExt_lo_1475};
  wire [15:0]         maskExt_lo_1476 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1476 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1476 = {maskExt_hi_1476, maskExt_lo_1476};
  wire [15:0]         maskExt_lo_1477 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1477 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1477 = {maskExt_hi_1477, maskExt_lo_1477};
  wire [15:0]         maskExt_lo_1478 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1478 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1478 = {maskExt_hi_1478, maskExt_lo_1478};
  wire [15:0]         maskExt_lo_1479 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1479 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1479 = {maskExt_hi_1479, maskExt_lo_1479};
  wire [15:0]         maskExt_lo_1480 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1480 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1480 = {maskExt_hi_1480, maskExt_lo_1480};
  wire [15:0]         maskExt_lo_1481 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1481 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1481 = {maskExt_hi_1481, maskExt_lo_1481};
  wire [15:0]         maskExt_lo_1482 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1482 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1482 = {maskExt_hi_1482, maskExt_lo_1482};
  wire [15:0]         maskExt_lo_1483 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1483 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1483 = {maskExt_hi_1483, maskExt_lo_1483};
  wire [15:0]         maskExt_lo_1484 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1484 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1484 = {maskExt_hi_1484, maskExt_lo_1484};
  wire [15:0]         maskExt_lo_1485 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1485 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1485 = {maskExt_hi_1485, maskExt_lo_1485};
  wire [15:0]         maskExt_lo_1486 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1486 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1486 = {maskExt_hi_1486, maskExt_lo_1486};
  wire [15:0]         maskExt_lo_1487 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1487 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1487 = {maskExt_hi_1487, maskExt_lo_1487};
  wire [15:0]         maskExt_lo_1488 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1488 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1488 = {maskExt_hi_1488, maskExt_lo_1488};
  wire [15:0]         maskExt_lo_1489 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1489 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1489 = {maskExt_hi_1489, maskExt_lo_1489};
  wire [15:0]         maskExt_lo_1490 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1490 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1490 = {maskExt_hi_1490, maskExt_lo_1490};
  wire [15:0]         maskExt_lo_1491 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1491 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1491 = {maskExt_hi_1491, maskExt_lo_1491};
  wire [15:0]         maskExt_lo_1492 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1492 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1492 = {maskExt_hi_1492, maskExt_lo_1492};
  wire [15:0]         maskExt_lo_1493 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1493 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1493 = {maskExt_hi_1493, maskExt_lo_1493};
  wire [15:0]         maskExt_lo_1494 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1494 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1494 = {maskExt_hi_1494, maskExt_lo_1494};
  wire [15:0]         maskExt_lo_1495 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1495 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1495 = {maskExt_hi_1495, maskExt_lo_1495};
  wire [15:0]         maskExt_lo_1496 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1496 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1496 = {maskExt_hi_1496, maskExt_lo_1496};
  wire [15:0]         maskExt_lo_1497 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1497 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1497 = {maskExt_hi_1497, maskExt_lo_1497};
  wire [15:0]         maskExt_lo_1498 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1498 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1498 = {maskExt_hi_1498, maskExt_lo_1498};
  wire [15:0]         maskExt_lo_1499 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1499 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1499 = {maskExt_hi_1499, maskExt_lo_1499};
  wire [15:0]         maskExt_lo_1500 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1500 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1500 = {maskExt_hi_1500, maskExt_lo_1500};
  wire [15:0]         maskExt_lo_1501 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1501 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1501 = {maskExt_hi_1501, maskExt_lo_1501};
  wire [15:0]         maskExt_lo_1502 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1502 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1502 = {maskExt_hi_1502, maskExt_lo_1502};
  wire [15:0]         maskExt_lo_1503 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1503 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1503 = {maskExt_hi_1503, maskExt_lo_1503};
  wire [15:0]         maskExt_lo_1504 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1504 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1504 = {maskExt_hi_1504, maskExt_lo_1504};
  wire [15:0]         maskExt_lo_1505 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1505 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1505 = {maskExt_hi_1505, maskExt_lo_1505};
  wire [15:0]         maskExt_lo_1506 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1506 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1506 = {maskExt_hi_1506, maskExt_lo_1506};
  wire [15:0]         maskExt_lo_1507 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1507 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1507 = {maskExt_hi_1507, maskExt_lo_1507};
  wire [15:0]         maskExt_lo_1508 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1508 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1508 = {maskExt_hi_1508, maskExt_lo_1508};
  wire [15:0]         maskExt_lo_1509 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1509 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1509 = {maskExt_hi_1509, maskExt_lo_1509};
  wire [15:0]         maskExt_lo_1510 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1510 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1510 = {maskExt_hi_1510, maskExt_lo_1510};
  wire [15:0]         maskExt_lo_1511 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1511 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1511 = {maskExt_hi_1511, maskExt_lo_1511};
  wire [15:0]         maskExt_lo_1512 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1512 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1512 = {maskExt_hi_1512, maskExt_lo_1512};
  wire [15:0]         maskExt_lo_1513 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1513 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1513 = {maskExt_hi_1513, maskExt_lo_1513};
  wire [15:0]         maskExt_lo_1514 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1514 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1514 = {maskExt_hi_1514, maskExt_lo_1514};
  wire [15:0]         maskExt_lo_1515 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1515 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1515 = {maskExt_hi_1515, maskExt_lo_1515};
  wire [15:0]         maskExt_lo_1516 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1516 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1516 = {maskExt_hi_1516, maskExt_lo_1516};
  wire [15:0]         maskExt_lo_1517 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1517 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1517 = {maskExt_hi_1517, maskExt_lo_1517};
  wire [15:0]         maskExt_lo_1518 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1518 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1518 = {maskExt_hi_1518, maskExt_lo_1518};
  wire [15:0]         maskExt_lo_1519 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1519 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1519 = {maskExt_hi_1519, maskExt_lo_1519};
  wire [15:0]         maskExt_lo_1520 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1520 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1520 = {maskExt_hi_1520, maskExt_lo_1520};
  wire [15:0]         maskExt_lo_1521 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1521 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1521 = {maskExt_hi_1521, maskExt_lo_1521};
  wire [15:0]         maskExt_lo_1522 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1522 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1522 = {maskExt_hi_1522, maskExt_lo_1522};
  wire [15:0]         maskExt_lo_1523 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1523 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1523 = {maskExt_hi_1523, maskExt_lo_1523};
  wire [15:0]         maskExt_lo_1524 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1524 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1524 = {maskExt_hi_1524, maskExt_lo_1524};
  wire [15:0]         maskExt_lo_1525 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1525 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1525 = {maskExt_hi_1525, maskExt_lo_1525};
  wire [15:0]         maskExt_lo_1526 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1526 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1526 = {maskExt_hi_1526, maskExt_lo_1526};
  wire [15:0]         maskExt_lo_1527 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1527 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1527 = {maskExt_hi_1527, maskExt_lo_1527};
  wire [15:0]         maskExt_lo_1528 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1528 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1528 = {maskExt_hi_1528, maskExt_lo_1528};
  wire [15:0]         maskExt_lo_1529 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1529 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1529 = {maskExt_hi_1529, maskExt_lo_1529};
  wire [15:0]         maskExt_lo_1530 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1530 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1530 = {maskExt_hi_1530, maskExt_lo_1530};
  wire [15:0]         maskExt_lo_1531 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1531 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1531 = {maskExt_hi_1531, maskExt_lo_1531};
  wire [15:0]         maskExt_lo_1532 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1532 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1532 = {maskExt_hi_1532, maskExt_lo_1532};
  wire [15:0]         maskExt_lo_1533 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1533 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1533 = {maskExt_hi_1533, maskExt_lo_1533};
  wire [15:0]         maskExt_lo_1534 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1534 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1534 = {maskExt_hi_1534, maskExt_lo_1534};
  wire [15:0]         maskExt_lo_1535 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1535 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1535 = {maskExt_hi_1535, maskExt_lo_1535};
  wire [15:0]         maskExt_lo_1536 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1536 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1536 = {maskExt_hi_1536, maskExt_lo_1536};
  wire [15:0]         maskExt_lo_1537 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1537 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1537 = {maskExt_hi_1537, maskExt_lo_1537};
  wire [15:0]         maskExt_lo_1538 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1538 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1538 = {maskExt_hi_1538, maskExt_lo_1538};
  wire [15:0]         maskExt_lo_1539 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1539 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1539 = {maskExt_hi_1539, maskExt_lo_1539};
  wire [15:0]         maskExt_lo_1540 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1540 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1540 = {maskExt_hi_1540, maskExt_lo_1540};
  wire [15:0]         maskExt_lo_1541 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1541 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1541 = {maskExt_hi_1541, maskExt_lo_1541};
  wire [15:0]         maskExt_lo_1542 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1542 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1542 = {maskExt_hi_1542, maskExt_lo_1542};
  wire [15:0]         maskExt_lo_1543 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1543 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1543 = {maskExt_hi_1543, maskExt_lo_1543};
  wire [15:0]         maskExt_lo_1544 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1544 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1544 = {maskExt_hi_1544, maskExt_lo_1544};
  wire [15:0]         maskExt_lo_1545 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1545 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1545 = {maskExt_hi_1545, maskExt_lo_1545};
  wire [15:0]         maskExt_lo_1546 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1546 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1546 = {maskExt_hi_1546, maskExt_lo_1546};
  wire [15:0]         maskExt_lo_1547 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1547 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1547 = {maskExt_hi_1547, maskExt_lo_1547};
  wire [15:0]         maskExt_lo_1548 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1548 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1548 = {maskExt_hi_1548, maskExt_lo_1548};
  wire [15:0]         maskExt_lo_1549 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1549 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1549 = {maskExt_hi_1549, maskExt_lo_1549};
  wire [15:0]         maskExt_lo_1550 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1550 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1550 = {maskExt_hi_1550, maskExt_lo_1550};
  wire [15:0]         maskExt_lo_1551 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1551 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1551 = {maskExt_hi_1551, maskExt_lo_1551};
  wire [15:0]         maskExt_lo_1552 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1552 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1552 = {maskExt_hi_1552, maskExt_lo_1552};
  wire [15:0]         maskExt_lo_1553 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1553 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1553 = {maskExt_hi_1553, maskExt_lo_1553};
  wire [15:0]         maskExt_lo_1554 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1554 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1554 = {maskExt_hi_1554, maskExt_lo_1554};
  wire [15:0]         maskExt_lo_1555 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1555 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1555 = {maskExt_hi_1555, maskExt_lo_1555};
  wire [15:0]         maskExt_lo_1556 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1556 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1556 = {maskExt_hi_1556, maskExt_lo_1556};
  wire [15:0]         maskExt_lo_1557 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1557 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1557 = {maskExt_hi_1557, maskExt_lo_1557};
  wire [15:0]         maskExt_lo_1558 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1558 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1558 = {maskExt_hi_1558, maskExt_lo_1558};
  wire [15:0]         maskExt_lo_1559 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1559 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1559 = {maskExt_hi_1559, maskExt_lo_1559};
  wire [15:0]         maskExt_lo_1560 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1560 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1560 = {maskExt_hi_1560, maskExt_lo_1560};
  wire [15:0]         maskExt_lo_1561 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1561 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1561 = {maskExt_hi_1561, maskExt_lo_1561};
  wire [15:0]         maskExt_lo_1562 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1562 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1562 = {maskExt_hi_1562, maskExt_lo_1562};
  wire [15:0]         maskExt_lo_1563 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1563 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1563 = {maskExt_hi_1563, maskExt_lo_1563};
  wire [15:0]         maskExt_lo_1564 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1564 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1564 = {maskExt_hi_1564, maskExt_lo_1564};
  wire [15:0]         maskExt_lo_1565 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1565 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1565 = {maskExt_hi_1565, maskExt_lo_1565};
  wire [15:0]         maskExt_lo_1566 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1566 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1566 = {maskExt_hi_1566, maskExt_lo_1566};
  wire [15:0]         maskExt_lo_1567 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1567 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1567 = {maskExt_hi_1567, maskExt_lo_1567};
  wire [15:0]         maskExt_lo_1568 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1568 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1568 = {maskExt_hi_1568, maskExt_lo_1568};
  wire [15:0]         maskExt_lo_1569 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1569 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1569 = {maskExt_hi_1569, maskExt_lo_1569};
  wire [15:0]         maskExt_lo_1570 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1570 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1570 = {maskExt_hi_1570, maskExt_lo_1570};
  wire [15:0]         maskExt_lo_1571 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1571 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1571 = {maskExt_hi_1571, maskExt_lo_1571};
  wire [15:0]         maskExt_lo_1572 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1572 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1572 = {maskExt_hi_1572, maskExt_lo_1572};
  wire [15:0]         maskExt_lo_1573 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1573 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1573 = {maskExt_hi_1573, maskExt_lo_1573};
  wire [15:0]         maskExt_lo_1574 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1574 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1574 = {maskExt_hi_1574, maskExt_lo_1574};
  wire [15:0]         maskExt_lo_1575 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1575 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1575 = {maskExt_hi_1575, maskExt_lo_1575};
  wire [15:0]         maskExt_lo_1576 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1576 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1576 = {maskExt_hi_1576, maskExt_lo_1576};
  wire [15:0]         maskExt_lo_1577 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1577 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1577 = {maskExt_hi_1577, maskExt_lo_1577};
  wire [15:0]         maskExt_lo_1578 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1578 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1578 = {maskExt_hi_1578, maskExt_lo_1578};
  wire [15:0]         maskExt_lo_1579 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1579 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1579 = {maskExt_hi_1579, maskExt_lo_1579};
  wire [15:0]         maskExt_lo_1580 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1580 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1580 = {maskExt_hi_1580, maskExt_lo_1580};
  wire [15:0]         maskExt_lo_1581 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1581 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1581 = {maskExt_hi_1581, maskExt_lo_1581};
  wire [15:0]         maskExt_lo_1582 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1582 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1582 = {maskExt_hi_1582, maskExt_lo_1582};
  wire [15:0]         maskExt_lo_1583 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1583 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1583 = {maskExt_hi_1583, maskExt_lo_1583};
  wire [15:0]         maskExt_lo_1584 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1584 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1584 = {maskExt_hi_1584, maskExt_lo_1584};
  wire [15:0]         maskExt_lo_1585 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1585 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1585 = {maskExt_hi_1585, maskExt_lo_1585};
  wire [15:0]         maskExt_lo_1586 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1586 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1586 = {maskExt_hi_1586, maskExt_lo_1586};
  wire [15:0]         maskExt_lo_1587 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1587 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1587 = {maskExt_hi_1587, maskExt_lo_1587};
  wire [15:0]         maskExt_lo_1588 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1588 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1588 = {maskExt_hi_1588, maskExt_lo_1588};
  wire [15:0]         maskExt_lo_1589 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1589 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1589 = {maskExt_hi_1589, maskExt_lo_1589};
  wire [15:0]         maskExt_lo_1590 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1590 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1590 = {maskExt_hi_1590, maskExt_lo_1590};
  wire [15:0]         maskExt_lo_1591 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1591 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1591 = {maskExt_hi_1591, maskExt_lo_1591};
  wire [15:0]         maskExt_lo_1592 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1592 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1592 = {maskExt_hi_1592, maskExt_lo_1592};
  wire [15:0]         maskExt_lo_1593 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1593 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1593 = {maskExt_hi_1593, maskExt_lo_1593};
  wire [15:0]         maskExt_lo_1594 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1594 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1594 = {maskExt_hi_1594, maskExt_lo_1594};
  wire [15:0]         maskExt_lo_1595 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1595 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1595 = {maskExt_hi_1595, maskExt_lo_1595};
  wire [15:0]         maskExt_lo_1596 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1596 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1596 = {maskExt_hi_1596, maskExt_lo_1596};
  wire [15:0]         maskExt_lo_1597 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1597 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1597 = {maskExt_hi_1597, maskExt_lo_1597};
  wire [15:0]         maskExt_lo_1598 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1598 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1598 = {maskExt_hi_1598, maskExt_lo_1598};
  wire [15:0]         maskExt_lo_1599 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1599 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1599 = {maskExt_hi_1599, maskExt_lo_1599};
  wire [15:0]         maskExt_lo_1600 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1600 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1600 = {maskExt_hi_1600, maskExt_lo_1600};
  wire [15:0]         maskExt_lo_1601 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1601 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1601 = {maskExt_hi_1601, maskExt_lo_1601};
  wire [15:0]         maskExt_lo_1602 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1602 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1602 = {maskExt_hi_1602, maskExt_lo_1602};
  wire [15:0]         maskExt_lo_1603 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1603 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1603 = {maskExt_hi_1603, maskExt_lo_1603};
  wire [15:0]         maskExt_lo_1604 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1604 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1604 = {maskExt_hi_1604, maskExt_lo_1604};
  wire [15:0]         maskExt_lo_1605 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1605 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1605 = {maskExt_hi_1605, maskExt_lo_1605};
  wire [15:0]         maskExt_lo_1606 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1606 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1606 = {maskExt_hi_1606, maskExt_lo_1606};
  wire [15:0]         maskExt_lo_1607 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1607 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1607 = {maskExt_hi_1607, maskExt_lo_1607};
  wire [15:0]         maskExt_lo_1608 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1608 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1608 = {maskExt_hi_1608, maskExt_lo_1608};
  wire [15:0]         maskExt_lo_1609 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1609 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1609 = {maskExt_hi_1609, maskExt_lo_1609};
  wire [15:0]         maskExt_lo_1610 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1610 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1610 = {maskExt_hi_1610, maskExt_lo_1610};
  wire [15:0]         maskExt_lo_1611 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1611 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1611 = {maskExt_hi_1611, maskExt_lo_1611};
  wire [15:0]         maskExt_lo_1612 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1612 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1612 = {maskExt_hi_1612, maskExt_lo_1612};
  wire [15:0]         maskExt_lo_1613 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1613 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1613 = {maskExt_hi_1613, maskExt_lo_1613};
  wire [15:0]         maskExt_lo_1614 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1614 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1614 = {maskExt_hi_1614, maskExt_lo_1614};
  wire [15:0]         maskExt_lo_1615 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1615 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1615 = {maskExt_hi_1615, maskExt_lo_1615};
  wire [15:0]         maskExt_lo_1616 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1616 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1616 = {maskExt_hi_1616, maskExt_lo_1616};
  wire [15:0]         maskExt_lo_1617 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1617 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1617 = {maskExt_hi_1617, maskExt_lo_1617};
  wire [15:0]         maskExt_lo_1618 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1618 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1618 = {maskExt_hi_1618, maskExt_lo_1618};
  wire [15:0]         maskExt_lo_1619 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1619 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1619 = {maskExt_hi_1619, maskExt_lo_1619};
  wire [15:0]         maskExt_lo_1620 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1620 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1620 = {maskExt_hi_1620, maskExt_lo_1620};
  wire [15:0]         maskExt_lo_1621 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1621 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1621 = {maskExt_hi_1621, maskExt_lo_1621};
  wire [15:0]         maskExt_lo_1622 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1622 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1622 = {maskExt_hi_1622, maskExt_lo_1622};
  wire [15:0]         maskExt_lo_1623 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1623 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1623 = {maskExt_hi_1623, maskExt_lo_1623};
  wire [15:0]         maskExt_lo_1624 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1624 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1624 = {maskExt_hi_1624, maskExt_lo_1624};
  wire [15:0]         maskExt_lo_1625 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1625 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1625 = {maskExt_hi_1625, maskExt_lo_1625};
  wire [15:0]         maskExt_lo_1626 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1626 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1626 = {maskExt_hi_1626, maskExt_lo_1626};
  wire [15:0]         maskExt_lo_1627 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1627 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1627 = {maskExt_hi_1627, maskExt_lo_1627};
  wire [15:0]         maskExt_lo_1628 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1628 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1628 = {maskExt_hi_1628, maskExt_lo_1628};
  wire [15:0]         maskExt_lo_1629 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1629 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1629 = {maskExt_hi_1629, maskExt_lo_1629};
  wire [15:0]         maskExt_lo_1630 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1630 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1630 = {maskExt_hi_1630, maskExt_lo_1630};
  wire [15:0]         maskExt_lo_1631 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1631 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1631 = {maskExt_hi_1631, maskExt_lo_1631};
  wire [15:0]         maskExt_lo_1632 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1632 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1632 = {maskExt_hi_1632, maskExt_lo_1632};
  wire [15:0]         maskExt_lo_1633 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1633 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1633 = {maskExt_hi_1633, maskExt_lo_1633};
  wire [15:0]         maskExt_lo_1634 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1634 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1634 = {maskExt_hi_1634, maskExt_lo_1634};
  wire [15:0]         maskExt_lo_1635 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1635 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1635 = {maskExt_hi_1635, maskExt_lo_1635};
  wire [15:0]         maskExt_lo_1636 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1636 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1636 = {maskExt_hi_1636, maskExt_lo_1636};
  wire [15:0]         maskExt_lo_1637 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1637 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1637 = {maskExt_hi_1637, maskExt_lo_1637};
  wire [15:0]         maskExt_lo_1638 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1638 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1638 = {maskExt_hi_1638, maskExt_lo_1638};
  wire [15:0]         maskExt_lo_1639 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1639 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1639 = {maskExt_hi_1639, maskExt_lo_1639};
  wire [15:0]         maskExt_lo_1640 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1640 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1640 = {maskExt_hi_1640, maskExt_lo_1640};
  wire [15:0]         maskExt_lo_1641 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1641 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1641 = {maskExt_hi_1641, maskExt_lo_1641};
  wire [15:0]         maskExt_lo_1642 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1642 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1642 = {maskExt_hi_1642, maskExt_lo_1642};
  wire [15:0]         maskExt_lo_1643 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1643 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1643 = {maskExt_hi_1643, maskExt_lo_1643};
  wire [15:0]         maskExt_lo_1644 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1644 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1644 = {maskExt_hi_1644, maskExt_lo_1644};
  wire [15:0]         maskExt_lo_1645 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1645 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1645 = {maskExt_hi_1645, maskExt_lo_1645};
  wire [15:0]         maskExt_lo_1646 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1646 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1646 = {maskExt_hi_1646, maskExt_lo_1646};
  wire [15:0]         maskExt_lo_1647 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1647 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1647 = {maskExt_hi_1647, maskExt_lo_1647};
  wire [15:0]         maskExt_lo_1648 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1648 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1648 = {maskExt_hi_1648, maskExt_lo_1648};
  wire [15:0]         maskExt_lo_1649 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1649 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1649 = {maskExt_hi_1649, maskExt_lo_1649};
  wire [15:0]         maskExt_lo_1650 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1650 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1650 = {maskExt_hi_1650, maskExt_lo_1650};
  wire [15:0]         maskExt_lo_1651 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1651 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1651 = {maskExt_hi_1651, maskExt_lo_1651};
  wire [15:0]         maskExt_lo_1652 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1652 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1652 = {maskExt_hi_1652, maskExt_lo_1652};
  wire [15:0]         maskExt_lo_1653 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1653 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1653 = {maskExt_hi_1653, maskExt_lo_1653};
  wire [15:0]         maskExt_lo_1654 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1654 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1654 = {maskExt_hi_1654, maskExt_lo_1654};
  wire [15:0]         maskExt_lo_1655 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1655 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1655 = {maskExt_hi_1655, maskExt_lo_1655};
  wire [15:0]         maskExt_lo_1656 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1656 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1656 = {maskExt_hi_1656, maskExt_lo_1656};
  wire [15:0]         maskExt_lo_1657 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1657 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1657 = {maskExt_hi_1657, maskExt_lo_1657};
  wire [15:0]         maskExt_lo_1658 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1658 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1658 = {maskExt_hi_1658, maskExt_lo_1658};
  wire [15:0]         maskExt_lo_1659 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1659 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1659 = {maskExt_hi_1659, maskExt_lo_1659};
  wire [15:0]         maskExt_lo_1660 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1660 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1660 = {maskExt_hi_1660, maskExt_lo_1660};
  wire [15:0]         maskExt_lo_1661 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1661 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1661 = {maskExt_hi_1661, maskExt_lo_1661};
  wire [15:0]         maskExt_lo_1662 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1662 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1662 = {maskExt_hi_1662, maskExt_lo_1662};
  wire [15:0]         maskExt_lo_1663 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1663 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1663 = {maskExt_hi_1663, maskExt_lo_1663};
  wire [15:0]         maskExt_lo_1664 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1664 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1664 = {maskExt_hi_1664, maskExt_lo_1664};
  wire [15:0]         maskExt_lo_1665 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1665 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1665 = {maskExt_hi_1665, maskExt_lo_1665};
  wire [15:0]         maskExt_lo_1666 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1666 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1666 = {maskExt_hi_1666, maskExt_lo_1666};
  wire [15:0]         maskExt_lo_1667 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1667 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1667 = {maskExt_hi_1667, maskExt_lo_1667};
  wire [15:0]         maskExt_lo_1668 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1668 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1668 = {maskExt_hi_1668, maskExt_lo_1668};
  wire [15:0]         maskExt_lo_1669 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1669 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1669 = {maskExt_hi_1669, maskExt_lo_1669};
  wire [15:0]         maskExt_lo_1670 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1670 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1670 = {maskExt_hi_1670, maskExt_lo_1670};
  wire [15:0]         maskExt_lo_1671 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1671 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1671 = {maskExt_hi_1671, maskExt_lo_1671};
  wire [15:0]         maskExt_lo_1672 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1672 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1672 = {maskExt_hi_1672, maskExt_lo_1672};
  wire [15:0]         maskExt_lo_1673 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1673 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1673 = {maskExt_hi_1673, maskExt_lo_1673};
  wire [15:0]         maskExt_lo_1674 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1674 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1674 = {maskExt_hi_1674, maskExt_lo_1674};
  wire [15:0]         maskExt_lo_1675 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1675 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1675 = {maskExt_hi_1675, maskExt_lo_1675};
  wire [15:0]         maskExt_lo_1676 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1676 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1676 = {maskExt_hi_1676, maskExt_lo_1676};
  wire [15:0]         maskExt_lo_1677 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1677 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1677 = {maskExt_hi_1677, maskExt_lo_1677};
  wire [15:0]         maskExt_lo_1678 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1678 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1678 = {maskExt_hi_1678, maskExt_lo_1678};
  wire [15:0]         maskExt_lo_1679 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1679 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1679 = {maskExt_hi_1679, maskExt_lo_1679};
  wire [15:0]         maskExt_lo_1680 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1680 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1680 = {maskExt_hi_1680, maskExt_lo_1680};
  wire [15:0]         maskExt_lo_1681 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1681 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1681 = {maskExt_hi_1681, maskExt_lo_1681};
  wire [15:0]         maskExt_lo_1682 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1682 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1682 = {maskExt_hi_1682, maskExt_lo_1682};
  wire [15:0]         maskExt_lo_1683 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1683 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1683 = {maskExt_hi_1683, maskExt_lo_1683};
  wire [15:0]         maskExt_lo_1684 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1684 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1684 = {maskExt_hi_1684, maskExt_lo_1684};
  wire [15:0]         maskExt_lo_1685 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1685 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1685 = {maskExt_hi_1685, maskExt_lo_1685};
  wire [15:0]         maskExt_lo_1686 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1686 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1686 = {maskExt_hi_1686, maskExt_lo_1686};
  wire [15:0]         maskExt_lo_1687 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1687 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1687 = {maskExt_hi_1687, maskExt_lo_1687};
  wire [15:0]         maskExt_lo_1688 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1688 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1688 = {maskExt_hi_1688, maskExt_lo_1688};
  wire [15:0]         maskExt_lo_1689 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1689 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1689 = {maskExt_hi_1689, maskExt_lo_1689};
  wire [15:0]         maskExt_lo_1690 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1690 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1690 = {maskExt_hi_1690, maskExt_lo_1690};
  wire [15:0]         maskExt_lo_1691 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1691 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1691 = {maskExt_hi_1691, maskExt_lo_1691};
  wire [15:0]         maskExt_lo_1692 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1692 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1692 = {maskExt_hi_1692, maskExt_lo_1692};
  wire [15:0]         maskExt_lo_1693 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1693 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1693 = {maskExt_hi_1693, maskExt_lo_1693};
  wire [15:0]         maskExt_lo_1694 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1694 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1694 = {maskExt_hi_1694, maskExt_lo_1694};
  wire [15:0]         maskExt_lo_1695 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1695 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1695 = {maskExt_hi_1695, maskExt_lo_1695};
  wire [15:0]         maskExt_lo_1696 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1696 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1696 = {maskExt_hi_1696, maskExt_lo_1696};
  wire [15:0]         maskExt_lo_1697 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1697 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1697 = {maskExt_hi_1697, maskExt_lo_1697};
  wire [15:0]         maskExt_lo_1698 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1698 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1698 = {maskExt_hi_1698, maskExt_lo_1698};
  wire [15:0]         maskExt_lo_1699 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1699 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1699 = {maskExt_hi_1699, maskExt_lo_1699};
  wire [15:0]         maskExt_lo_1700 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1700 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1700 = {maskExt_hi_1700, maskExt_lo_1700};
  wire [15:0]         maskExt_lo_1701 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1701 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1701 = {maskExt_hi_1701, maskExt_lo_1701};
  wire [15:0]         maskExt_lo_1702 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1702 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1702 = {maskExt_hi_1702, maskExt_lo_1702};
  wire [15:0]         maskExt_lo_1703 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1703 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1703 = {maskExt_hi_1703, maskExt_lo_1703};
  wire [15:0]         maskExt_lo_1704 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1704 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1704 = {maskExt_hi_1704, maskExt_lo_1704};
  wire [15:0]         maskExt_lo_1705 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1705 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1705 = {maskExt_hi_1705, maskExt_lo_1705};
  wire [15:0]         maskExt_lo_1706 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1706 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1706 = {maskExt_hi_1706, maskExt_lo_1706};
  wire [15:0]         maskExt_lo_1707 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1707 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1707 = {maskExt_hi_1707, maskExt_lo_1707};
  wire [15:0]         maskExt_lo_1708 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1708 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1708 = {maskExt_hi_1708, maskExt_lo_1708};
  wire [15:0]         maskExt_lo_1709 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1709 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1709 = {maskExt_hi_1709, maskExt_lo_1709};
  wire [15:0]         maskExt_lo_1710 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1710 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1710 = {maskExt_hi_1710, maskExt_lo_1710};
  wire [15:0]         maskExt_lo_1711 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1711 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1711 = {maskExt_hi_1711, maskExt_lo_1711};
  wire [15:0]         maskExt_lo_1712 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1712 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1712 = {maskExt_hi_1712, maskExt_lo_1712};
  wire [15:0]         maskExt_lo_1713 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1713 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1713 = {maskExt_hi_1713, maskExt_lo_1713};
  wire [15:0]         maskExt_lo_1714 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1714 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1714 = {maskExt_hi_1714, maskExt_lo_1714};
  wire [15:0]         maskExt_lo_1715 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1715 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1715 = {maskExt_hi_1715, maskExt_lo_1715};
  wire [15:0]         maskExt_lo_1716 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1716 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1716 = {maskExt_hi_1716, maskExt_lo_1716};
  wire [15:0]         maskExt_lo_1717 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1717 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1717 = {maskExt_hi_1717, maskExt_lo_1717};
  wire [15:0]         maskExt_lo_1718 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1718 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1718 = {maskExt_hi_1718, maskExt_lo_1718};
  wire [15:0]         maskExt_lo_1719 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1719 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1719 = {maskExt_hi_1719, maskExt_lo_1719};
  wire [15:0]         maskExt_lo_1720 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1720 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1720 = {maskExt_hi_1720, maskExt_lo_1720};
  wire [15:0]         maskExt_lo_1721 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1721 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1721 = {maskExt_hi_1721, maskExt_lo_1721};
  wire [15:0]         maskExt_lo_1722 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1722 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1722 = {maskExt_hi_1722, maskExt_lo_1722};
  wire [15:0]         maskExt_lo_1723 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1723 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1723 = {maskExt_hi_1723, maskExt_lo_1723};
  wire [15:0]         maskExt_lo_1724 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1724 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1724 = {maskExt_hi_1724, maskExt_lo_1724};
  wire [15:0]         maskExt_lo_1725 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1725 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1725 = {maskExt_hi_1725, maskExt_lo_1725};
  wire [15:0]         maskExt_lo_1726 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1726 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1726 = {maskExt_hi_1726, maskExt_lo_1726};
  wire [15:0]         maskExt_lo_1727 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1727 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1727 = {maskExt_hi_1727, maskExt_lo_1727};
  wire [15:0]         maskExt_lo_1728 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1728 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1728 = {maskExt_hi_1728, maskExt_lo_1728};
  wire [15:0]         maskExt_lo_1729 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1729 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1729 = {maskExt_hi_1729, maskExt_lo_1729};
  wire [15:0]         maskExt_lo_1730 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1730 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1730 = {maskExt_hi_1730, maskExt_lo_1730};
  wire [15:0]         maskExt_lo_1731 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1731 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1731 = {maskExt_hi_1731, maskExt_lo_1731};
  wire [15:0]         maskExt_lo_1732 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1732 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1732 = {maskExt_hi_1732, maskExt_lo_1732};
  wire [15:0]         maskExt_lo_1733 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1733 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1733 = {maskExt_hi_1733, maskExt_lo_1733};
  wire [15:0]         maskExt_lo_1734 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1734 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1734 = {maskExt_hi_1734, maskExt_lo_1734};
  wire [15:0]         maskExt_lo_1735 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1735 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1735 = {maskExt_hi_1735, maskExt_lo_1735};
  wire [15:0]         maskExt_lo_1736 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1736 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1736 = {maskExt_hi_1736, maskExt_lo_1736};
  wire [15:0]         maskExt_lo_1737 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1737 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1737 = {maskExt_hi_1737, maskExt_lo_1737};
  wire [15:0]         maskExt_lo_1738 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1738 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1738 = {maskExt_hi_1738, maskExt_lo_1738};
  wire [15:0]         maskExt_lo_1739 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1739 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1739 = {maskExt_hi_1739, maskExt_lo_1739};
  wire [15:0]         maskExt_lo_1740 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1740 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1740 = {maskExt_hi_1740, maskExt_lo_1740};
  wire [15:0]         maskExt_lo_1741 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1741 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1741 = {maskExt_hi_1741, maskExt_lo_1741};
  wire [15:0]         maskExt_lo_1742 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1742 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1742 = {maskExt_hi_1742, maskExt_lo_1742};
  wire [15:0]         maskExt_lo_1743 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1743 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1743 = {maskExt_hi_1743, maskExt_lo_1743};
  wire [15:0]         maskExt_lo_1744 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1744 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1744 = {maskExt_hi_1744, maskExt_lo_1744};
  wire [15:0]         maskExt_lo_1745 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1745 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1745 = {maskExt_hi_1745, maskExt_lo_1745};
  wire [15:0]         maskExt_lo_1746 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1746 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1746 = {maskExt_hi_1746, maskExt_lo_1746};
  wire [15:0]         maskExt_lo_1747 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1747 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1747 = {maskExt_hi_1747, maskExt_lo_1747};
  wire [15:0]         maskExt_lo_1748 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1748 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1748 = {maskExt_hi_1748, maskExt_lo_1748};
  wire [15:0]         maskExt_lo_1749 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1749 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1749 = {maskExt_hi_1749, maskExt_lo_1749};
  wire [15:0]         maskExt_lo_1750 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1750 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1750 = {maskExt_hi_1750, maskExt_lo_1750};
  wire [15:0]         maskExt_lo_1751 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1751 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1751 = {maskExt_hi_1751, maskExt_lo_1751};
  wire [15:0]         maskExt_lo_1752 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1752 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1752 = {maskExt_hi_1752, maskExt_lo_1752};
  wire [15:0]         maskExt_lo_1753 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1753 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1753 = {maskExt_hi_1753, maskExt_lo_1753};
  wire [15:0]         maskExt_lo_1754 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1754 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1754 = {maskExt_hi_1754, maskExt_lo_1754};
  wire [15:0]         maskExt_lo_1755 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1755 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1755 = {maskExt_hi_1755, maskExt_lo_1755};
  wire [15:0]         maskExt_lo_1756 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1756 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1756 = {maskExt_hi_1756, maskExt_lo_1756};
  wire [15:0]         maskExt_lo_1757 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1757 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1757 = {maskExt_hi_1757, maskExt_lo_1757};
  wire [15:0]         maskExt_lo_1758 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1758 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1758 = {maskExt_hi_1758, maskExt_lo_1758};
  wire [15:0]         maskExt_lo_1759 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1759 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1759 = {maskExt_hi_1759, maskExt_lo_1759};
  wire [15:0]         maskExt_lo_1760 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1760 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1760 = {maskExt_hi_1760, maskExt_lo_1760};
  wire [15:0]         maskExt_lo_1761 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1761 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1761 = {maskExt_hi_1761, maskExt_lo_1761};
  wire [15:0]         maskExt_lo_1762 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1762 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1762 = {maskExt_hi_1762, maskExt_lo_1762};
  wire [15:0]         maskExt_lo_1763 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1763 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1763 = {maskExt_hi_1763, maskExt_lo_1763};
  wire [15:0]         maskExt_lo_1764 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1764 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1764 = {maskExt_hi_1764, maskExt_lo_1764};
  wire [15:0]         maskExt_lo_1765 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1765 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1765 = {maskExt_hi_1765, maskExt_lo_1765};
  wire [15:0]         maskExt_lo_1766 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1766 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1766 = {maskExt_hi_1766, maskExt_lo_1766};
  wire [15:0]         maskExt_lo_1767 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1767 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1767 = {maskExt_hi_1767, maskExt_lo_1767};
  wire [15:0]         maskExt_lo_1768 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1768 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1768 = {maskExt_hi_1768, maskExt_lo_1768};
  wire [15:0]         maskExt_lo_1769 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1769 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1769 = {maskExt_hi_1769, maskExt_lo_1769};
  wire [15:0]         maskExt_lo_1770 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1770 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1770 = {maskExt_hi_1770, maskExt_lo_1770};
  wire [15:0]         maskExt_lo_1771 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1771 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1771 = {maskExt_hi_1771, maskExt_lo_1771};
  wire [15:0]         maskExt_lo_1772 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1772 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1772 = {maskExt_hi_1772, maskExt_lo_1772};
  wire [15:0]         maskExt_lo_1773 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1773 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1773 = {maskExt_hi_1773, maskExt_lo_1773};
  wire [15:0]         maskExt_lo_1774 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1774 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1774 = {maskExt_hi_1774, maskExt_lo_1774};
  wire [15:0]         maskExt_lo_1775 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1775 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1775 = {maskExt_hi_1775, maskExt_lo_1775};
  wire [15:0]         maskExt_lo_1776 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1776 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1776 = {maskExt_hi_1776, maskExt_lo_1776};
  wire [15:0]         maskExt_lo_1777 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1777 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1777 = {maskExt_hi_1777, maskExt_lo_1777};
  wire [15:0]         maskExt_lo_1778 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1778 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1778 = {maskExt_hi_1778, maskExt_lo_1778};
  wire [15:0]         maskExt_lo_1779 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1779 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1779 = {maskExt_hi_1779, maskExt_lo_1779};
  wire [15:0]         maskExt_lo_1780 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1780 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1780 = {maskExt_hi_1780, maskExt_lo_1780};
  wire [15:0]         maskExt_lo_1781 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1781 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1781 = {maskExt_hi_1781, maskExt_lo_1781};
  wire [15:0]         maskExt_lo_1782 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1782 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1782 = {maskExt_hi_1782, maskExt_lo_1782};
  wire [15:0]         maskExt_lo_1783 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1783 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1783 = {maskExt_hi_1783, maskExt_lo_1783};
  wire [15:0]         maskExt_lo_1784 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1784 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1784 = {maskExt_hi_1784, maskExt_lo_1784};
  wire [15:0]         maskExt_lo_1785 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1785 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1785 = {maskExt_hi_1785, maskExt_lo_1785};
  wire [15:0]         maskExt_lo_1786 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1786 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1786 = {maskExt_hi_1786, maskExt_lo_1786};
  wire [15:0]         maskExt_lo_1787 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1787 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1787 = {maskExt_hi_1787, maskExt_lo_1787};
  wire [15:0]         maskExt_lo_1788 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1788 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1788 = {maskExt_hi_1788, maskExt_lo_1788};
  wire [15:0]         maskExt_lo_1789 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1789 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1789 = {maskExt_hi_1789, maskExt_lo_1789};
  wire [15:0]         maskExt_lo_1790 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1790 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1790 = {maskExt_hi_1790, maskExt_lo_1790};
  wire [15:0]         maskExt_lo_1791 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1791 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1791 = {maskExt_hi_1791, maskExt_lo_1791};
  wire [15:0]         maskExt_lo_1792 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1792 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1792 = {maskExt_hi_1792, maskExt_lo_1792};
  wire [15:0]         maskExt_lo_1793 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1793 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1793 = {maskExt_hi_1793, maskExt_lo_1793};
  wire [15:0]         maskExt_lo_1794 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1794 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1794 = {maskExt_hi_1794, maskExt_lo_1794};
  wire [15:0]         maskExt_lo_1795 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1795 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1795 = {maskExt_hi_1795, maskExt_lo_1795};
  wire [15:0]         maskExt_lo_1796 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1796 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1796 = {maskExt_hi_1796, maskExt_lo_1796};
  wire [15:0]         maskExt_lo_1797 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1797 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1797 = {maskExt_hi_1797, maskExt_lo_1797};
  wire [15:0]         maskExt_lo_1798 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1798 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1798 = {maskExt_hi_1798, maskExt_lo_1798};
  wire [15:0]         maskExt_lo_1799 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1799 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1799 = {maskExt_hi_1799, maskExt_lo_1799};
  wire [15:0]         maskExt_lo_1800 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1800 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1800 = {maskExt_hi_1800, maskExt_lo_1800};
  wire [15:0]         maskExt_lo_1801 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1801 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1801 = {maskExt_hi_1801, maskExt_lo_1801};
  wire [15:0]         maskExt_lo_1802 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1802 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1802 = {maskExt_hi_1802, maskExt_lo_1802};
  wire [15:0]         maskExt_lo_1803 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1803 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1803 = {maskExt_hi_1803, maskExt_lo_1803};
  wire [15:0]         maskExt_lo_1804 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1804 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1804 = {maskExt_hi_1804, maskExt_lo_1804};
  wire [15:0]         maskExt_lo_1805 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1805 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1805 = {maskExt_hi_1805, maskExt_lo_1805};
  wire [15:0]         maskExt_lo_1806 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1806 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1806 = {maskExt_hi_1806, maskExt_lo_1806};
  wire [15:0]         maskExt_lo_1807 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1807 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1807 = {maskExt_hi_1807, maskExt_lo_1807};
  wire [15:0]         maskExt_lo_1808 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1808 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1808 = {maskExt_hi_1808, maskExt_lo_1808};
  wire [15:0]         maskExt_lo_1809 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1809 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1809 = {maskExt_hi_1809, maskExt_lo_1809};
  wire [15:0]         maskExt_lo_1810 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1810 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1810 = {maskExt_hi_1810, maskExt_lo_1810};
  wire [15:0]         maskExt_lo_1811 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1811 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1811 = {maskExt_hi_1811, maskExt_lo_1811};
  wire [15:0]         maskExt_lo_1812 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1812 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1812 = {maskExt_hi_1812, maskExt_lo_1812};
  wire [15:0]         maskExt_lo_1813 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1813 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1813 = {maskExt_hi_1813, maskExt_lo_1813};
  wire [15:0]         maskExt_lo_1814 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1814 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1814 = {maskExt_hi_1814, maskExt_lo_1814};
  wire [15:0]         maskExt_lo_1815 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1815 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1815 = {maskExt_hi_1815, maskExt_lo_1815};
  wire [15:0]         maskExt_lo_1816 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1816 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1816 = {maskExt_hi_1816, maskExt_lo_1816};
  wire [15:0]         maskExt_lo_1817 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1817 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1817 = {maskExt_hi_1817, maskExt_lo_1817};
  wire [15:0]         maskExt_lo_1818 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1818 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1818 = {maskExt_hi_1818, maskExt_lo_1818};
  wire [15:0]         maskExt_lo_1819 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1819 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1819 = {maskExt_hi_1819, maskExt_lo_1819};
  wire [15:0]         maskExt_lo_1820 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1820 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1820 = {maskExt_hi_1820, maskExt_lo_1820};
  wire [15:0]         maskExt_lo_1821 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1821 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1821 = {maskExt_hi_1821, maskExt_lo_1821};
  wire [15:0]         maskExt_lo_1822 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1822 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1822 = {maskExt_hi_1822, maskExt_lo_1822};
  wire [15:0]         maskExt_lo_1823 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1823 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1823 = {maskExt_hi_1823, maskExt_lo_1823};
  wire [15:0]         maskExt_lo_1824 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1824 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1824 = {maskExt_hi_1824, maskExt_lo_1824};
  wire [15:0]         maskExt_lo_1825 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1825 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1825 = {maskExt_hi_1825, maskExt_lo_1825};
  wire [15:0]         maskExt_lo_1826 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1826 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1826 = {maskExt_hi_1826, maskExt_lo_1826};
  wire [15:0]         maskExt_lo_1827 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1827 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1827 = {maskExt_hi_1827, maskExt_lo_1827};
  wire [15:0]         maskExt_lo_1828 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1828 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1828 = {maskExt_hi_1828, maskExt_lo_1828};
  wire [15:0]         maskExt_lo_1829 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1829 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1829 = {maskExt_hi_1829, maskExt_lo_1829};
  wire [15:0]         maskExt_lo_1830 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1830 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1830 = {maskExt_hi_1830, maskExt_lo_1830};
  wire [15:0]         maskExt_lo_1831 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1831 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1831 = {maskExt_hi_1831, maskExt_lo_1831};
  wire [15:0]         maskExt_lo_1832 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1832 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1832 = {maskExt_hi_1832, maskExt_lo_1832};
  wire [15:0]         maskExt_lo_1833 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1833 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1833 = {maskExt_hi_1833, maskExt_lo_1833};
  wire [15:0]         maskExt_lo_1834 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1834 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1834 = {maskExt_hi_1834, maskExt_lo_1834};
  wire [15:0]         maskExt_lo_1835 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1835 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1835 = {maskExt_hi_1835, maskExt_lo_1835};
  wire [15:0]         maskExt_lo_1836 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1836 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1836 = {maskExt_hi_1836, maskExt_lo_1836};
  wire [15:0]         maskExt_lo_1837 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1837 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1837 = {maskExt_hi_1837, maskExt_lo_1837};
  wire [15:0]         maskExt_lo_1838 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1838 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1838 = {maskExt_hi_1838, maskExt_lo_1838};
  wire [15:0]         maskExt_lo_1839 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1839 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1839 = {maskExt_hi_1839, maskExt_lo_1839};
  wire [15:0]         maskExt_lo_1840 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1840 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1840 = {maskExt_hi_1840, maskExt_lo_1840};
  wire [15:0]         maskExt_lo_1841 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1841 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1841 = {maskExt_hi_1841, maskExt_lo_1841};
  wire [15:0]         maskExt_lo_1842 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1842 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1842 = {maskExt_hi_1842, maskExt_lo_1842};
  wire [15:0]         maskExt_lo_1843 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1843 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1843 = {maskExt_hi_1843, maskExt_lo_1843};
  wire [15:0]         maskExt_lo_1844 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1844 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1844 = {maskExt_hi_1844, maskExt_lo_1844};
  wire [15:0]         maskExt_lo_1845 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1845 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1845 = {maskExt_hi_1845, maskExt_lo_1845};
  wire [15:0]         maskExt_lo_1846 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1846 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1846 = {maskExt_hi_1846, maskExt_lo_1846};
  wire [15:0]         maskExt_lo_1847 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1847 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1847 = {maskExt_hi_1847, maskExt_lo_1847};
  wire [15:0]         maskExt_lo_1848 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1848 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1848 = {maskExt_hi_1848, maskExt_lo_1848};
  wire [15:0]         maskExt_lo_1849 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1849 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1849 = {maskExt_hi_1849, maskExt_lo_1849};
  wire [15:0]         maskExt_lo_1850 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1850 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1850 = {maskExt_hi_1850, maskExt_lo_1850};
  wire [15:0]         maskExt_lo_1851 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1851 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1851 = {maskExt_hi_1851, maskExt_lo_1851};
  wire [15:0]         maskExt_lo_1852 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1852 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1852 = {maskExt_hi_1852, maskExt_lo_1852};
  wire [15:0]         maskExt_lo_1853 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1853 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1853 = {maskExt_hi_1853, maskExt_lo_1853};
  wire [15:0]         maskExt_lo_1854 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1854 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1854 = {maskExt_hi_1854, maskExt_lo_1854};
  wire [15:0]         maskExt_lo_1855 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1855 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1855 = {maskExt_hi_1855, maskExt_lo_1855};
  wire [15:0]         maskExt_lo_1856 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1856 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1856 = {maskExt_hi_1856, maskExt_lo_1856};
  wire [15:0]         maskExt_lo_1857 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1857 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1857 = {maskExt_hi_1857, maskExt_lo_1857};
  wire [15:0]         maskExt_lo_1858 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1858 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1858 = {maskExt_hi_1858, maskExt_lo_1858};
  wire [15:0]         maskExt_lo_1859 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1859 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1859 = {maskExt_hi_1859, maskExt_lo_1859};
  wire [15:0]         maskExt_lo_1860 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1860 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1860 = {maskExt_hi_1860, maskExt_lo_1860};
  wire [15:0]         maskExt_lo_1861 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1861 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1861 = {maskExt_hi_1861, maskExt_lo_1861};
  wire [15:0]         maskExt_lo_1862 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1862 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1862 = {maskExt_hi_1862, maskExt_lo_1862};
  wire [15:0]         maskExt_lo_1863 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1863 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1863 = {maskExt_hi_1863, maskExt_lo_1863};
  wire [15:0]         maskExt_lo_1864 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1864 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1864 = {maskExt_hi_1864, maskExt_lo_1864};
  wire [15:0]         maskExt_lo_1865 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1865 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1865 = {maskExt_hi_1865, maskExt_lo_1865};
  wire [15:0]         maskExt_lo_1866 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1866 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1866 = {maskExt_hi_1866, maskExt_lo_1866};
  wire [15:0]         maskExt_lo_1867 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1867 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1867 = {maskExt_hi_1867, maskExt_lo_1867};
  wire [15:0]         maskExt_lo_1868 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1868 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1868 = {maskExt_hi_1868, maskExt_lo_1868};
  wire [15:0]         maskExt_lo_1869 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1869 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1869 = {maskExt_hi_1869, maskExt_lo_1869};
  wire [15:0]         maskExt_lo_1870 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1870 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1870 = {maskExt_hi_1870, maskExt_lo_1870};
  wire [15:0]         maskExt_lo_1871 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1871 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1871 = {maskExt_hi_1871, maskExt_lo_1871};
  wire [15:0]         maskExt_lo_1872 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1872 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1872 = {maskExt_hi_1872, maskExt_lo_1872};
  wire [15:0]         maskExt_lo_1873 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1873 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1873 = {maskExt_hi_1873, maskExt_lo_1873};
  wire [15:0]         maskExt_lo_1874 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1874 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1874 = {maskExt_hi_1874, maskExt_lo_1874};
  wire [15:0]         maskExt_lo_1875 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1875 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1875 = {maskExt_hi_1875, maskExt_lo_1875};
  wire [15:0]         maskExt_lo_1876 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1876 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1876 = {maskExt_hi_1876, maskExt_lo_1876};
  wire [15:0]         maskExt_lo_1877 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1877 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1877 = {maskExt_hi_1877, maskExt_lo_1877};
  wire [15:0]         maskExt_lo_1878 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1878 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1878 = {maskExt_hi_1878, maskExt_lo_1878};
  wire [15:0]         maskExt_lo_1879 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1879 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1879 = {maskExt_hi_1879, maskExt_lo_1879};
  wire [15:0]         maskExt_lo_1880 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1880 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1880 = {maskExt_hi_1880, maskExt_lo_1880};
  wire [15:0]         maskExt_lo_1881 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1881 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1881 = {maskExt_hi_1881, maskExt_lo_1881};
  wire [15:0]         maskExt_lo_1882 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1882 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1882 = {maskExt_hi_1882, maskExt_lo_1882};
  wire [15:0]         maskExt_lo_1883 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1883 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1883 = {maskExt_hi_1883, maskExt_lo_1883};
  wire [15:0]         maskExt_lo_1884 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1884 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1884 = {maskExt_hi_1884, maskExt_lo_1884};
  wire [15:0]         maskExt_lo_1885 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1885 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1885 = {maskExt_hi_1885, maskExt_lo_1885};
  wire [15:0]         maskExt_lo_1886 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1886 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1886 = {maskExt_hi_1886, maskExt_lo_1886};
  wire [15:0]         maskExt_lo_1887 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1887 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1887 = {maskExt_hi_1887, maskExt_lo_1887};
  wire [15:0]         maskExt_lo_1888 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1888 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1888 = {maskExt_hi_1888, maskExt_lo_1888};
  wire [15:0]         maskExt_lo_1889 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1889 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1889 = {maskExt_hi_1889, maskExt_lo_1889};
  wire [15:0]         maskExt_lo_1890 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1890 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1890 = {maskExt_hi_1890, maskExt_lo_1890};
  wire [15:0]         maskExt_lo_1891 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1891 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1891 = {maskExt_hi_1891, maskExt_lo_1891};
  wire [15:0]         maskExt_lo_1892 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1892 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1892 = {maskExt_hi_1892, maskExt_lo_1892};
  wire [15:0]         maskExt_lo_1893 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1893 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1893 = {maskExt_hi_1893, maskExt_lo_1893};
  wire [15:0]         maskExt_lo_1894 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1894 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1894 = {maskExt_hi_1894, maskExt_lo_1894};
  wire [15:0]         maskExt_lo_1895 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1895 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1895 = {maskExt_hi_1895, maskExt_lo_1895};
  wire [15:0]         maskExt_lo_1896 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1896 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1896 = {maskExt_hi_1896, maskExt_lo_1896};
  wire [15:0]         maskExt_lo_1897 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1897 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1897 = {maskExt_hi_1897, maskExt_lo_1897};
  wire [15:0]         maskExt_lo_1898 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1898 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1898 = {maskExt_hi_1898, maskExt_lo_1898};
  wire [15:0]         maskExt_lo_1899 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1899 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1899 = {maskExt_hi_1899, maskExt_lo_1899};
  wire [15:0]         maskExt_lo_1900 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1900 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1900 = {maskExt_hi_1900, maskExt_lo_1900};
  wire [15:0]         maskExt_lo_1901 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1901 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1901 = {maskExt_hi_1901, maskExt_lo_1901};
  wire [15:0]         maskExt_lo_1902 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1902 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1902 = {maskExt_hi_1902, maskExt_lo_1902};
  wire [15:0]         maskExt_lo_1903 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1903 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1903 = {maskExt_hi_1903, maskExt_lo_1903};
  wire [15:0]         maskExt_lo_1904 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1904 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1904 = {maskExt_hi_1904, maskExt_lo_1904};
  wire [15:0]         maskExt_lo_1905 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1905 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1905 = {maskExt_hi_1905, maskExt_lo_1905};
  wire [15:0]         maskExt_lo_1906 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1906 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1906 = {maskExt_hi_1906, maskExt_lo_1906};
  wire [15:0]         maskExt_lo_1907 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1907 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1907 = {maskExt_hi_1907, maskExt_lo_1907};
  wire [15:0]         maskExt_lo_1908 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1908 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1908 = {maskExt_hi_1908, maskExt_lo_1908};
  wire [15:0]         maskExt_lo_1909 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1909 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1909 = {maskExt_hi_1909, maskExt_lo_1909};
  wire [15:0]         maskExt_lo_1910 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1910 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1910 = {maskExt_hi_1910, maskExt_lo_1910};
  wire [15:0]         maskExt_lo_1911 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1911 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1911 = {maskExt_hi_1911, maskExt_lo_1911};
  wire [15:0]         maskExt_lo_1912 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1912 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1912 = {maskExt_hi_1912, maskExt_lo_1912};
  wire [15:0]         maskExt_lo_1913 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1913 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1913 = {maskExt_hi_1913, maskExt_lo_1913};
  wire [15:0]         maskExt_lo_1914 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1914 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1914 = {maskExt_hi_1914, maskExt_lo_1914};
  wire [15:0]         maskExt_lo_1915 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1915 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1915 = {maskExt_hi_1915, maskExt_lo_1915};
  wire [15:0]         maskExt_lo_1916 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1916 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1916 = {maskExt_hi_1916, maskExt_lo_1916};
  wire [15:0]         maskExt_lo_1917 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1917 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1917 = {maskExt_hi_1917, maskExt_lo_1917};
  wire [15:0]         maskExt_lo_1918 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1918 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1918 = {maskExt_hi_1918, maskExt_lo_1918};
  wire [15:0]         maskExt_lo_1919 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1919 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1919 = {maskExt_hi_1919, maskExt_lo_1919};
  wire [15:0]         maskExt_lo_1920 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1920 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1920 = {maskExt_hi_1920, maskExt_lo_1920};
  wire [15:0]         maskExt_lo_1921 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1921 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1921 = {maskExt_hi_1921, maskExt_lo_1921};
  wire [15:0]         maskExt_lo_1922 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1922 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1922 = {maskExt_hi_1922, maskExt_lo_1922};
  wire [15:0]         maskExt_lo_1923 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1923 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1923 = {maskExt_hi_1923, maskExt_lo_1923};
  wire [15:0]         maskExt_lo_1924 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1924 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1924 = {maskExt_hi_1924, maskExt_lo_1924};
  wire [15:0]         maskExt_lo_1925 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1925 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1925 = {maskExt_hi_1925, maskExt_lo_1925};
  wire [15:0]         maskExt_lo_1926 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1926 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1926 = {maskExt_hi_1926, maskExt_lo_1926};
  wire [15:0]         maskExt_lo_1927 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1927 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1927 = {maskExt_hi_1927, maskExt_lo_1927};
  wire [15:0]         maskExt_lo_1928 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1928 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1928 = {maskExt_hi_1928, maskExt_lo_1928};
  wire [15:0]         maskExt_lo_1929 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1929 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1929 = {maskExt_hi_1929, maskExt_lo_1929};
  wire [15:0]         maskExt_lo_1930 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1930 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1930 = {maskExt_hi_1930, maskExt_lo_1930};
  wire [15:0]         maskExt_lo_1931 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1931 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1931 = {maskExt_hi_1931, maskExt_lo_1931};
  wire [15:0]         maskExt_lo_1932 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1932 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1932 = {maskExt_hi_1932, maskExt_lo_1932};
  wire [15:0]         maskExt_lo_1933 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1933 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1933 = {maskExt_hi_1933, maskExt_lo_1933};
  wire [15:0]         maskExt_lo_1934 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1934 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1934 = {maskExt_hi_1934, maskExt_lo_1934};
  wire [15:0]         maskExt_lo_1935 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1935 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1935 = {maskExt_hi_1935, maskExt_lo_1935};
  wire [15:0]         maskExt_lo_1936 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1936 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1936 = {maskExt_hi_1936, maskExt_lo_1936};
  wire [15:0]         maskExt_lo_1937 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1937 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1937 = {maskExt_hi_1937, maskExt_lo_1937};
  wire [15:0]         maskExt_lo_1938 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1938 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1938 = {maskExt_hi_1938, maskExt_lo_1938};
  wire [15:0]         maskExt_lo_1939 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1939 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1939 = {maskExt_hi_1939, maskExt_lo_1939};
  wire [15:0]         maskExt_lo_1940 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1940 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1940 = {maskExt_hi_1940, maskExt_lo_1940};
  wire [15:0]         maskExt_lo_1941 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1941 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1941 = {maskExt_hi_1941, maskExt_lo_1941};
  wire [15:0]         maskExt_lo_1942 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1942 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1942 = {maskExt_hi_1942, maskExt_lo_1942};
  wire [15:0]         maskExt_lo_1943 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1943 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1943 = {maskExt_hi_1943, maskExt_lo_1943};
  wire [15:0]         maskExt_lo_1944 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1944 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1944 = {maskExt_hi_1944, maskExt_lo_1944};
  wire [15:0]         maskExt_lo_1945 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1945 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1945 = {maskExt_hi_1945, maskExt_lo_1945};
  wire [15:0]         maskExt_lo_1946 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1946 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1946 = {maskExt_hi_1946, maskExt_lo_1946};
  wire [15:0]         maskExt_lo_1947 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1947 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1947 = {maskExt_hi_1947, maskExt_lo_1947};
  wire [15:0]         maskExt_lo_1948 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1948 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1948 = {maskExt_hi_1948, maskExt_lo_1948};
  wire [15:0]         maskExt_lo_1949 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1949 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1949 = {maskExt_hi_1949, maskExt_lo_1949};
  wire [15:0]         maskExt_lo_1950 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1950 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1950 = {maskExt_hi_1950, maskExt_lo_1950};
  wire [15:0]         maskExt_lo_1951 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1951 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1951 = {maskExt_hi_1951, maskExt_lo_1951};
  wire [15:0]         maskExt_lo_1952 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1952 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1952 = {maskExt_hi_1952, maskExt_lo_1952};
  wire [15:0]         maskExt_lo_1953 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1953 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1953 = {maskExt_hi_1953, maskExt_lo_1953};
  wire [15:0]         maskExt_lo_1954 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1954 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1954 = {maskExt_hi_1954, maskExt_lo_1954};
  wire [15:0]         maskExt_lo_1955 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1955 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1955 = {maskExt_hi_1955, maskExt_lo_1955};
  wire [15:0]         maskExt_lo_1956 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1956 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1956 = {maskExt_hi_1956, maskExt_lo_1956};
  wire [15:0]         maskExt_lo_1957 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1957 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1957 = {maskExt_hi_1957, maskExt_lo_1957};
  wire [15:0]         maskExt_lo_1958 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1958 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1958 = {maskExt_hi_1958, maskExt_lo_1958};
  wire [15:0]         maskExt_lo_1959 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1959 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1959 = {maskExt_hi_1959, maskExt_lo_1959};
  wire [15:0]         maskExt_lo_1960 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1960 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1960 = {maskExt_hi_1960, maskExt_lo_1960};
  wire [15:0]         maskExt_lo_1961 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1961 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1961 = {maskExt_hi_1961, maskExt_lo_1961};
  wire [15:0]         maskExt_lo_1962 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1962 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1962 = {maskExt_hi_1962, maskExt_lo_1962};
  wire [15:0]         maskExt_lo_1963 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1963 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1963 = {maskExt_hi_1963, maskExt_lo_1963};
  wire [15:0]         maskExt_lo_1964 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1964 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1964 = {maskExt_hi_1964, maskExt_lo_1964};
  wire [15:0]         maskExt_lo_1965 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1965 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1965 = {maskExt_hi_1965, maskExt_lo_1965};
  wire [15:0]         maskExt_lo_1966 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1966 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1966 = {maskExt_hi_1966, maskExt_lo_1966};
  wire [15:0]         maskExt_lo_1967 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1967 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1967 = {maskExt_hi_1967, maskExt_lo_1967};
  wire [15:0]         maskExt_lo_1968 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1968 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1968 = {maskExt_hi_1968, maskExt_lo_1968};
  wire [15:0]         maskExt_lo_1969 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1969 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1969 = {maskExt_hi_1969, maskExt_lo_1969};
  wire [15:0]         maskExt_lo_1970 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1970 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1970 = {maskExt_hi_1970, maskExt_lo_1970};
  wire [15:0]         maskExt_lo_1971 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1971 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1971 = {maskExt_hi_1971, maskExt_lo_1971};
  wire [15:0]         maskExt_lo_1972 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1972 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1972 = {maskExt_hi_1972, maskExt_lo_1972};
  wire [15:0]         maskExt_lo_1973 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1973 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1973 = {maskExt_hi_1973, maskExt_lo_1973};
  wire [15:0]         maskExt_lo_1974 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1974 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1974 = {maskExt_hi_1974, maskExt_lo_1974};
  wire [15:0]         maskExt_lo_1975 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1975 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1975 = {maskExt_hi_1975, maskExt_lo_1975};
  wire [15:0]         maskExt_lo_1976 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1976 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1976 = {maskExt_hi_1976, maskExt_lo_1976};
  wire [15:0]         maskExt_lo_1977 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1977 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1977 = {maskExt_hi_1977, maskExt_lo_1977};
  wire [15:0]         maskExt_lo_1978 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1978 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1978 = {maskExt_hi_1978, maskExt_lo_1978};
  wire [15:0]         maskExt_lo_1979 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1979 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1979 = {maskExt_hi_1979, maskExt_lo_1979};
  wire [15:0]         maskExt_lo_1980 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1980 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1980 = {maskExt_hi_1980, maskExt_lo_1980};
  wire [15:0]         maskExt_lo_1981 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1981 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1981 = {maskExt_hi_1981, maskExt_lo_1981};
  wire [15:0]         maskExt_lo_1982 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1982 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1982 = {maskExt_hi_1982, maskExt_lo_1982};
  wire [15:0]         maskExt_lo_1983 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1983 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1983 = {maskExt_hi_1983, maskExt_lo_1983};
  wire [15:0]         maskExt_lo_1984 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1984 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1984 = {maskExt_hi_1984, maskExt_lo_1984};
  wire [15:0]         maskExt_lo_1985 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1985 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1985 = {maskExt_hi_1985, maskExt_lo_1985};
  wire [15:0]         maskExt_lo_1986 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1986 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1986 = {maskExt_hi_1986, maskExt_lo_1986};
  wire [15:0]         maskExt_lo_1987 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1987 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1987 = {maskExt_hi_1987, maskExt_lo_1987};
  wire [15:0]         maskExt_lo_1988 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1988 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1988 = {maskExt_hi_1988, maskExt_lo_1988};
  wire [15:0]         maskExt_lo_1989 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1989 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1989 = {maskExt_hi_1989, maskExt_lo_1989};
  wire [15:0]         maskExt_lo_1990 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1990 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1990 = {maskExt_hi_1990, maskExt_lo_1990};
  wire [15:0]         maskExt_lo_1991 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1991 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1991 = {maskExt_hi_1991, maskExt_lo_1991};
  wire [15:0]         maskExt_lo_1992 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1992 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1992 = {maskExt_hi_1992, maskExt_lo_1992};
  wire [15:0]         maskExt_lo_1993 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1993 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1993 = {maskExt_hi_1993, maskExt_lo_1993};
  wire [15:0]         maskExt_lo_1994 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1994 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1994 = {maskExt_hi_1994, maskExt_lo_1994};
  wire [15:0]         maskExt_lo_1995 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1995 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1995 = {maskExt_hi_1995, maskExt_lo_1995};
  wire [15:0]         maskExt_lo_1996 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1996 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1996 = {maskExt_hi_1996, maskExt_lo_1996};
  wire [15:0]         maskExt_lo_1997 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1997 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1997 = {maskExt_hi_1997, maskExt_lo_1997};
  wire [15:0]         maskExt_lo_1998 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1998 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1998 = {maskExt_hi_1998, maskExt_lo_1998};
  wire [15:0]         maskExt_lo_1999 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1999 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1999 = {maskExt_hi_1999, maskExt_lo_1999};
  wire [15:0]         maskExt_lo_2000 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2000 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_2000 = {maskExt_hi_2000, maskExt_lo_2000};
  wire [15:0]         maskExt_lo_2001 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2001 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_2001 = {maskExt_hi_2001, maskExt_lo_2001};
  wire [15:0]         maskExt_lo_2002 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2002 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_2002 = {maskExt_hi_2002, maskExt_lo_2002};
  wire [15:0]         maskExt_lo_2003 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2003 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_2003 = {maskExt_hi_2003, maskExt_lo_2003};
  wire [15:0]         maskExt_lo_2004 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2004 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_2004 = {maskExt_hi_2004, maskExt_lo_2004};
  wire [15:0]         maskExt_lo_2005 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2005 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_2005 = {maskExt_hi_2005, maskExt_lo_2005};
  wire [15:0]         maskExt_lo_2006 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2006 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_2006 = {maskExt_hi_2006, maskExt_lo_2006};
  wire [15:0]         maskExt_lo_2007 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2007 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_2007 = {maskExt_hi_2007, maskExt_lo_2007};
  wire [15:0]         maskExt_lo_2008 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2008 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_2008 = {maskExt_hi_2008, maskExt_lo_2008};
  wire [15:0]         maskExt_lo_2009 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2009 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_2009 = {maskExt_hi_2009, maskExt_lo_2009};
  wire [15:0]         maskExt_lo_2010 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2010 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_2010 = {maskExt_hi_2010, maskExt_lo_2010};
  wire [15:0]         maskExt_lo_2011 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2011 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_2011 = {maskExt_hi_2011, maskExt_lo_2011};
  wire [15:0]         maskExt_lo_2012 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2012 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_2012 = {maskExt_hi_2012, maskExt_lo_2012};
  wire [15:0]         maskExt_lo_2013 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2013 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_2013 = {maskExt_hi_2013, maskExt_lo_2013};
  wire [15:0]         maskExt_lo_2014 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2014 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_2014 = {maskExt_hi_2014, maskExt_lo_2014};
  wire [15:0]         maskExt_lo_2015 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2015 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_2015 = {maskExt_hi_2015, maskExt_lo_2015};
  wire [15:0]         maskExt_lo_2016 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2016 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_2016 = {maskExt_hi_2016, maskExt_lo_2016};
  wire [15:0]         maskExt_lo_2017 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2017 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_2017 = {maskExt_hi_2017, maskExt_lo_2017};
  wire [15:0]         maskExt_lo_2018 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2018 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_2018 = {maskExt_hi_2018, maskExt_lo_2018};
  wire [15:0]         maskExt_lo_2019 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2019 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_2019 = {maskExt_hi_2019, maskExt_lo_2019};
  wire [15:0]         maskExt_lo_2020 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2020 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_2020 = {maskExt_hi_2020, maskExt_lo_2020};
  wire [15:0]         maskExt_lo_2021 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2021 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_2021 = {maskExt_hi_2021, maskExt_lo_2021};
  wire [15:0]         maskExt_lo_2022 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2022 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_2022 = {maskExt_hi_2022, maskExt_lo_2022};
  wire [15:0]         maskExt_lo_2023 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2023 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_2023 = {maskExt_hi_2023, maskExt_lo_2023};
  wire [15:0]         maskExt_lo_2024 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2024 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_2024 = {maskExt_hi_2024, maskExt_lo_2024};
  wire [15:0]         maskExt_lo_2025 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2025 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_2025 = {maskExt_hi_2025, maskExt_lo_2025};
  wire [15:0]         maskExt_lo_2026 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2026 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_2026 = {maskExt_hi_2026, maskExt_lo_2026};
  wire [15:0]         maskExt_lo_2027 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2027 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_2027 = {maskExt_hi_2027, maskExt_lo_2027};
  wire [15:0]         maskExt_lo_2028 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2028 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_2028 = {maskExt_hi_2028, maskExt_lo_2028};
  wire [15:0]         maskExt_lo_2029 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2029 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_2029 = {maskExt_hi_2029, maskExt_lo_2029};
  wire [15:0]         maskExt_lo_2030 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2030 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_2030 = {maskExt_hi_2030, maskExt_lo_2030};
  wire [15:0]         maskExt_lo_2031 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2031 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_2031 = {maskExt_hi_2031, maskExt_lo_2031};
  wire [15:0]         maskExt_lo_2032 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2032 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_2032 = {maskExt_hi_2032, maskExt_lo_2032};
  wire [15:0]         maskExt_lo_2033 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2033 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_2033 = {maskExt_hi_2033, maskExt_lo_2033};
  wire [15:0]         maskExt_lo_2034 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2034 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_2034 = {maskExt_hi_2034, maskExt_lo_2034};
  wire [15:0]         maskExt_lo_2035 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2035 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_2035 = {maskExt_hi_2035, maskExt_lo_2035};
  wire [15:0]         maskExt_lo_2036 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2036 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_2036 = {maskExt_hi_2036, maskExt_lo_2036};
  wire [15:0]         maskExt_lo_2037 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2037 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_2037 = {maskExt_hi_2037, maskExt_lo_2037};
  wire [15:0]         maskExt_lo_2038 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2038 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_2038 = {maskExt_hi_2038, maskExt_lo_2038};
  wire [15:0]         maskExt_lo_2039 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2039 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_2039 = {maskExt_hi_2039, maskExt_lo_2039};
  wire [15:0]         maskExt_lo_2040 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2040 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_2040 = {maskExt_hi_2040, maskExt_lo_2040};
  wire [15:0]         maskExt_lo_2041 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2041 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_2041 = {maskExt_hi_2041, maskExt_lo_2041};
  wire [15:0]         maskExt_lo_2042 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2042 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_2042 = {maskExt_hi_2042, maskExt_lo_2042};
  wire [15:0]         maskExt_lo_2043 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2043 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_2043 = {maskExt_hi_2043, maskExt_lo_2043};
  wire [15:0]         maskExt_lo_2044 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2044 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_2044 = {maskExt_hi_2044, maskExt_lo_2044};
  wire [15:0]         maskExt_lo_2045 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2045 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_2045 = {maskExt_hi_2045, maskExt_lo_2045};
  wire [15:0]         maskExt_lo_2046 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2046 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_2046 = {maskExt_hi_2046, maskExt_lo_2046};
  wire [15:0]         maskExt_lo_2047 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2047 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_2047 = {maskExt_hi_2047, maskExt_lo_2047};
  wire                alwaysMerge = {request_bits_instructionInformation_mop_0, request_bits_instructionInformation_lumop_0[2:0], request_bits_instructionInformation_lumop_0[4]} == 6'h0;
  wire                useLoadUnit = alwaysMerge & ~request_bits_instructionInformation_isStore_0;
  wire                useStoreUnit = alwaysMerge & request_bits_instructionInformation_isStore_0;
  wire                useOtherUnit = ~alwaysMerge;
  wire                addressCheck = _otherUnit_status_idle & (~useOtherUnit | _loadUnit_status_idle & _storeUnit_status_idle);
  wire                unitReady = useLoadUnit & _loadUnit_status_idle | useStoreUnit & _storeUnit_status_idle | useOtherUnit & _otherUnit_status_idle;
  wire                request_ready_0 = unitReady & addressCheck;
  wire                requestFire = request_ready_0 & request_valid_0;
  wire                reqEnq_0 = useLoadUnit & requestFire;
  wire                reqEnq_1 = useStoreUnit & requestFire;
  wire                reqEnq_2 = useOtherUnit & requestFire;
  wire [11:0]         maskSelect = _loadUnit_maskSelect_valid ? _loadUnit_maskSelect_bits : 12'h0;
  wire [63:0]         _GEN = {v0_1, v0_0};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo_lo = _GEN;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo_lo = _GEN;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo_lo = _GEN;
  wire [63:0]         _GEN_0 = {v0_3, v0_2};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo_hi = _GEN_0;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo_hi = _GEN_0;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo_hi = _GEN_0;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_1 = {v0_5, v0_4};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi_lo = _GEN_1;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi_lo = _GEN_1;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi_lo = _GEN_1;
  wire [63:0]         _GEN_2 = {v0_7, v0_6};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi_hi = _GEN_2;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi_hi = _GEN_2;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi_hi = _GEN_2;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi = {loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_3 = {v0_9, v0_8};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo_lo = _GEN_3;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo_lo = _GEN_3;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo_lo = _GEN_3;
  wire [63:0]         _GEN_4 = {v0_11, v0_10};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo_hi = _GEN_4;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo_hi = _GEN_4;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo_hi = _GEN_4;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo = {loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_5 = {v0_13, v0_12};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi_lo = _GEN_5;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi_lo = _GEN_5;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi_lo = _GEN_5;
  wire [63:0]         _GEN_6 = {v0_15, v0_14};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi_hi = _GEN_6;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi_hi = _GEN_6;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi_hi = _GEN_6;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi = {loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi = {loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_7 = {v0_17, v0_16};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo_lo = _GEN_7;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo_lo = _GEN_7;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo_lo = _GEN_7;
  wire [63:0]         _GEN_8 = {v0_19, v0_18};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo_hi = _GEN_8;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo_hi = _GEN_8;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo_hi = _GEN_8;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo = {loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_9 = {v0_21, v0_20};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi_lo = _GEN_9;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi_lo = _GEN_9;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi_lo = _GEN_9;
  wire [63:0]         _GEN_10 = {v0_23, v0_22};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi_hi = _GEN_10;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi_hi = _GEN_10;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi_hi = _GEN_10;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi = {loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo = {loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_11 = {v0_25, v0_24};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo_lo = _GEN_11;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo_lo = _GEN_11;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo_lo = _GEN_11;
  wire [63:0]         _GEN_12 = {v0_27, v0_26};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo_hi = _GEN_12;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo_hi = _GEN_12;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo_hi = _GEN_12;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo = {loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_13 = {v0_29, v0_28};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi_lo = _GEN_13;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi_lo = _GEN_13;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi_lo = _GEN_13;
  wire [63:0]         _GEN_14 = {v0_31, v0_30};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi_hi = _GEN_14;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi_hi = _GEN_14;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi_hi = _GEN_14;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi = {loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi = {loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi = {loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_lo_lo_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_15 = {v0_33, v0_32};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo_lo = _GEN_15;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo_lo = _GEN_15;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo_lo = _GEN_15;
  wire [63:0]         _GEN_16 = {v0_35, v0_34};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo_hi = _GEN_16;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo_hi = _GEN_16;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo_hi = _GEN_16;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_17 = {v0_37, v0_36};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi_lo = _GEN_17;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi_lo = _GEN_17;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi_lo = _GEN_17;
  wire [63:0]         _GEN_18 = {v0_39, v0_38};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi_hi = _GEN_18;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi_hi = _GEN_18;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi_hi = _GEN_18;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi = {loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo = {loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_19 = {v0_41, v0_40};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo_lo = _GEN_19;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo_lo = _GEN_19;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo_lo = _GEN_19;
  wire [63:0]         _GEN_20 = {v0_43, v0_42};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo_hi = _GEN_20;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo_hi = _GEN_20;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo_hi = _GEN_20;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo = {loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_21 = {v0_45, v0_44};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi_lo = _GEN_21;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi_lo = _GEN_21;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi_lo = _GEN_21;
  wire [63:0]         _GEN_22 = {v0_47, v0_46};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi_hi = _GEN_22;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi_hi = _GEN_22;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi_hi = _GEN_22;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi = {loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi = {loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo = {loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_23 = {v0_49, v0_48};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo_lo = _GEN_23;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo_lo = _GEN_23;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo_lo = _GEN_23;
  wire [63:0]         _GEN_24 = {v0_51, v0_50};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo_hi = _GEN_24;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo_hi = _GEN_24;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo_hi = _GEN_24;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo = {loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_25 = {v0_53, v0_52};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi_lo = _GEN_25;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi_lo = _GEN_25;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi_lo = _GEN_25;
  wire [63:0]         _GEN_26 = {v0_55, v0_54};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi_hi = _GEN_26;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi_hi = _GEN_26;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi_hi = _GEN_26;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi = {loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo = {loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_27 = {v0_57, v0_56};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo_lo = _GEN_27;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo_lo = _GEN_27;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo_lo = _GEN_27;
  wire [63:0]         _GEN_28 = {v0_59, v0_58};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo_hi = _GEN_28;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo_hi = _GEN_28;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo_hi = _GEN_28;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo = {loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_29 = {v0_61, v0_60};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi_lo = _GEN_29;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi_lo = _GEN_29;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi_lo = _GEN_29;
  wire [63:0]         _GEN_30 = {v0_63, v0_62};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi_hi = _GEN_30;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi_hi = _GEN_30;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi_hi = _GEN_30;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi = {loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi = {loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi = {loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_lo_lo_lo_lo_hi = {loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo};
  wire [2047:0]       loadUnit_maskInput_lo_lo_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_31 = {v0_65, v0_64};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo_lo = _GEN_31;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo_lo = _GEN_31;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo_lo = _GEN_31;
  wire [63:0]         _GEN_32 = {v0_67, v0_66};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo_hi = _GEN_32;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo_hi = _GEN_32;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo_hi = _GEN_32;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_33 = {v0_69, v0_68};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi_lo = _GEN_33;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi_lo = _GEN_33;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi_lo = _GEN_33;
  wire [63:0]         _GEN_34 = {v0_71, v0_70};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi_hi = _GEN_34;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi_hi = _GEN_34;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi_hi = _GEN_34;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi = {loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_35 = {v0_73, v0_72};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo_lo = _GEN_35;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo_lo = _GEN_35;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo_lo = _GEN_35;
  wire [63:0]         _GEN_36 = {v0_75, v0_74};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo_hi = _GEN_36;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo_hi = _GEN_36;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo_hi = _GEN_36;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo = {loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_37 = {v0_77, v0_76};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi_lo = _GEN_37;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi_lo = _GEN_37;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi_lo = _GEN_37;
  wire [63:0]         _GEN_38 = {v0_79, v0_78};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi_hi = _GEN_38;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi_hi = _GEN_38;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi_hi = _GEN_38;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi = {loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi = {loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo = {loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_39 = {v0_81, v0_80};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo_lo = _GEN_39;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo_lo = _GEN_39;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo_lo = _GEN_39;
  wire [63:0]         _GEN_40 = {v0_83, v0_82};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo_hi = _GEN_40;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo_hi = _GEN_40;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo_hi = _GEN_40;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo = {loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_41 = {v0_85, v0_84};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi_lo = _GEN_41;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi_lo = _GEN_41;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi_lo = _GEN_41;
  wire [63:0]         _GEN_42 = {v0_87, v0_86};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi_hi = _GEN_42;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi_hi = _GEN_42;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi_hi = _GEN_42;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi = {loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo = {loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_43 = {v0_89, v0_88};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo_lo = _GEN_43;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo_lo = _GEN_43;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo_lo = _GEN_43;
  wire [63:0]         _GEN_44 = {v0_91, v0_90};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo_hi = _GEN_44;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo_hi = _GEN_44;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo_hi = _GEN_44;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo = {loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_45 = {v0_93, v0_92};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi_lo = _GEN_45;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi_lo = _GEN_45;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi_lo = _GEN_45;
  wire [63:0]         _GEN_46 = {v0_95, v0_94};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi_hi = _GEN_46;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi_hi = _GEN_46;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi_hi = _GEN_46;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi = {loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi = {loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi = {loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_lo_lo_lo_hi_lo = {loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_47 = {v0_97, v0_96};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo_lo = _GEN_47;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo_lo = _GEN_47;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo_lo = _GEN_47;
  wire [63:0]         _GEN_48 = {v0_99, v0_98};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo_hi = _GEN_48;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo_hi = _GEN_48;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo_hi = _GEN_48;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_49 = {v0_101, v0_100};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi_lo = _GEN_49;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi_lo = _GEN_49;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi_lo = _GEN_49;
  wire [63:0]         _GEN_50 = {v0_103, v0_102};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi_hi = _GEN_50;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi_hi = _GEN_50;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi_hi = _GEN_50;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi = {loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo = {loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_51 = {v0_105, v0_104};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo_lo = _GEN_51;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo_lo = _GEN_51;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo_lo = _GEN_51;
  wire [63:0]         _GEN_52 = {v0_107, v0_106};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo_hi = _GEN_52;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo_hi = _GEN_52;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo_hi = _GEN_52;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo = {loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_53 = {v0_109, v0_108};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi_lo = _GEN_53;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi_lo = _GEN_53;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi_lo = _GEN_53;
  wire [63:0]         _GEN_54 = {v0_111, v0_110};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi_hi = _GEN_54;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi_hi = _GEN_54;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi_hi = _GEN_54;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi = {loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi = {loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo = {loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_55 = {v0_113, v0_112};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo_lo = _GEN_55;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo_lo = _GEN_55;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo_lo = _GEN_55;
  wire [63:0]         _GEN_56 = {v0_115, v0_114};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo_hi = _GEN_56;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo_hi = _GEN_56;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo_hi = _GEN_56;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo = {loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_57 = {v0_117, v0_116};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi_lo = _GEN_57;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi_lo = _GEN_57;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi_lo = _GEN_57;
  wire [63:0]         _GEN_58 = {v0_119, v0_118};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi_hi = _GEN_58;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi_hi = _GEN_58;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi_hi = _GEN_58;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi = {loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo = {loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_59 = {v0_121, v0_120};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo_lo = _GEN_59;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo_lo = _GEN_59;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo_lo = _GEN_59;
  wire [63:0]         _GEN_60 = {v0_123, v0_122};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo_hi = _GEN_60;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo_hi = _GEN_60;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo_hi = _GEN_60;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo = {loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_61 = {v0_125, v0_124};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi_lo = _GEN_61;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi_lo = _GEN_61;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi_lo = _GEN_61;
  wire [63:0]         _GEN_62 = {v0_127, v0_126};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi_hi = _GEN_62;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi_hi = _GEN_62;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi_hi = _GEN_62;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi = {loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi = {loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi = {loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_lo_lo_lo_hi_hi = {loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo};
  wire [2047:0]       loadUnit_maskInput_lo_lo_lo_lo_hi = {loadUnit_maskInput_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_lo};
  wire [4095:0]       loadUnit_maskInput_lo_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_63 = {v0_129, v0_128};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo_lo = _GEN_63;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo_lo = _GEN_63;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo_lo = _GEN_63;
  wire [63:0]         _GEN_64 = {v0_131, v0_130};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo_hi = _GEN_64;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo_hi = _GEN_64;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo_hi = _GEN_64;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_65 = {v0_133, v0_132};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi_lo = _GEN_65;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi_lo = _GEN_65;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi_lo = _GEN_65;
  wire [63:0]         _GEN_66 = {v0_135, v0_134};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi_hi = _GEN_66;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi_hi = _GEN_66;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi_hi = _GEN_66;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi = {loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_67 = {v0_137, v0_136};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo_lo = _GEN_67;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo_lo = _GEN_67;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo_lo = _GEN_67;
  wire [63:0]         _GEN_68 = {v0_139, v0_138};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo_hi = _GEN_68;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo_hi = _GEN_68;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo_hi = _GEN_68;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo = {loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_69 = {v0_141, v0_140};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi_lo = _GEN_69;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi_lo = _GEN_69;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi_lo = _GEN_69;
  wire [63:0]         _GEN_70 = {v0_143, v0_142};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi_hi = _GEN_70;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi_hi = _GEN_70;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi_hi = _GEN_70;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi = {loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi = {loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_71 = {v0_145, v0_144};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo_lo = _GEN_71;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo_lo = _GEN_71;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo_lo = _GEN_71;
  wire [63:0]         _GEN_72 = {v0_147, v0_146};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo_hi = _GEN_72;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo_hi = _GEN_72;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo_hi = _GEN_72;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo = {loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_73 = {v0_149, v0_148};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi_lo = _GEN_73;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi_lo = _GEN_73;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi_lo = _GEN_73;
  wire [63:0]         _GEN_74 = {v0_151, v0_150};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi_hi = _GEN_74;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi_hi = _GEN_74;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi_hi = _GEN_74;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi = {loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo = {loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_75 = {v0_153, v0_152};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo_lo = _GEN_75;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo_lo = _GEN_75;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo_lo = _GEN_75;
  wire [63:0]         _GEN_76 = {v0_155, v0_154};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo_hi = _GEN_76;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo_hi = _GEN_76;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo_hi = _GEN_76;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo = {loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_77 = {v0_157, v0_156};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi_lo = _GEN_77;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi_lo = _GEN_77;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi_lo = _GEN_77;
  wire [63:0]         _GEN_78 = {v0_159, v0_158};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi_hi = _GEN_78;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi_hi = _GEN_78;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi_hi = _GEN_78;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi = {loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi = {loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi = {loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_lo_lo_hi_lo_lo = {loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_79 = {v0_161, v0_160};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo_lo = _GEN_79;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo_lo = _GEN_79;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo_lo = _GEN_79;
  wire [63:0]         _GEN_80 = {v0_163, v0_162};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo_hi = _GEN_80;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo_hi = _GEN_80;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo_hi = _GEN_80;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_81 = {v0_165, v0_164};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi_lo = _GEN_81;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi_lo = _GEN_81;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi_lo = _GEN_81;
  wire [63:0]         _GEN_82 = {v0_167, v0_166};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi_hi = _GEN_82;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi_hi = _GEN_82;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi_hi = _GEN_82;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi = {loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo = {loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_83 = {v0_169, v0_168};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo_lo = _GEN_83;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo_lo = _GEN_83;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo_lo = _GEN_83;
  wire [63:0]         _GEN_84 = {v0_171, v0_170};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo_hi = _GEN_84;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo_hi = _GEN_84;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo_hi = _GEN_84;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo = {loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_85 = {v0_173, v0_172};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi_lo = _GEN_85;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi_lo = _GEN_85;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi_lo = _GEN_85;
  wire [63:0]         _GEN_86 = {v0_175, v0_174};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi_hi = _GEN_86;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi_hi = _GEN_86;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi_hi = _GEN_86;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi = {loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi = {loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo = {loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_87 = {v0_177, v0_176};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo_lo = _GEN_87;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo_lo = _GEN_87;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo_lo = _GEN_87;
  wire [63:0]         _GEN_88 = {v0_179, v0_178};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo_hi = _GEN_88;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo_hi = _GEN_88;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo_hi = _GEN_88;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo = {loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_89 = {v0_181, v0_180};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi_lo = _GEN_89;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi_lo = _GEN_89;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi_lo = _GEN_89;
  wire [63:0]         _GEN_90 = {v0_183, v0_182};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi_hi = _GEN_90;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi_hi = _GEN_90;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi_hi = _GEN_90;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi = {loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo = {loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_91 = {v0_185, v0_184};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo_lo = _GEN_91;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo_lo = _GEN_91;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo_lo = _GEN_91;
  wire [63:0]         _GEN_92 = {v0_187, v0_186};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo_hi = _GEN_92;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo_hi = _GEN_92;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo_hi = _GEN_92;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo = {loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_93 = {v0_189, v0_188};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi_lo = _GEN_93;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi_lo = _GEN_93;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi_lo = _GEN_93;
  wire [63:0]         _GEN_94 = {v0_191, v0_190};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi_hi = _GEN_94;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi_hi = _GEN_94;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi_hi = _GEN_94;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi = {loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi = {loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi = {loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_lo_lo_hi_lo_hi = {loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo};
  wire [2047:0]       loadUnit_maskInput_lo_lo_lo_hi_lo = {loadUnit_maskInput_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_95 = {v0_193, v0_192};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo_lo = _GEN_95;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo_lo = _GEN_95;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo_lo = _GEN_95;
  wire [63:0]         _GEN_96 = {v0_195, v0_194};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo_hi = _GEN_96;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo_hi = _GEN_96;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo_hi = _GEN_96;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_97 = {v0_197, v0_196};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi_lo = _GEN_97;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi_lo = _GEN_97;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi_lo = _GEN_97;
  wire [63:0]         _GEN_98 = {v0_199, v0_198};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi_hi = _GEN_98;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi_hi = _GEN_98;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi_hi = _GEN_98;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi = {loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_99 = {v0_201, v0_200};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo_lo = _GEN_99;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo_lo = _GEN_99;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo_lo = _GEN_99;
  wire [63:0]         _GEN_100 = {v0_203, v0_202};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo_hi = _GEN_100;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo_hi = _GEN_100;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo_hi = _GEN_100;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo = {loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_101 = {v0_205, v0_204};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi_lo = _GEN_101;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi_lo = _GEN_101;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi_lo = _GEN_101;
  wire [63:0]         _GEN_102 = {v0_207, v0_206};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi_hi = _GEN_102;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi_hi = _GEN_102;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi_hi = _GEN_102;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi = {loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi = {loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo = {loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_103 = {v0_209, v0_208};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo_lo = _GEN_103;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo_lo = _GEN_103;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo_lo = _GEN_103;
  wire [63:0]         _GEN_104 = {v0_211, v0_210};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo_hi = _GEN_104;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo_hi = _GEN_104;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo_hi = _GEN_104;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo = {loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_105 = {v0_213, v0_212};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi_lo = _GEN_105;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi_lo = _GEN_105;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi_lo = _GEN_105;
  wire [63:0]         _GEN_106 = {v0_215, v0_214};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi_hi = _GEN_106;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi_hi = _GEN_106;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi_hi = _GEN_106;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi = {loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo = {loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_107 = {v0_217, v0_216};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo_lo = _GEN_107;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo_lo = _GEN_107;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo_lo = _GEN_107;
  wire [63:0]         _GEN_108 = {v0_219, v0_218};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo_hi = _GEN_108;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo_hi = _GEN_108;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo_hi = _GEN_108;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo = {loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_109 = {v0_221, v0_220};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi_lo = _GEN_109;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi_lo = _GEN_109;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi_lo = _GEN_109;
  wire [63:0]         _GEN_110 = {v0_223, v0_222};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi_hi = _GEN_110;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi_hi = _GEN_110;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi_hi = _GEN_110;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi = {loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi = {loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi = {loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_lo_lo_hi_hi_lo = {loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_111 = {v0_225, v0_224};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo_lo = _GEN_111;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo_lo = _GEN_111;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo_lo = _GEN_111;
  wire [63:0]         _GEN_112 = {v0_227, v0_226};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo_hi = _GEN_112;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo_hi = _GEN_112;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo_hi = _GEN_112;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_113 = {v0_229, v0_228};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi_lo = _GEN_113;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi_lo = _GEN_113;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi_lo = _GEN_113;
  wire [63:0]         _GEN_114 = {v0_231, v0_230};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi_hi = _GEN_114;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi_hi = _GEN_114;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi_hi = _GEN_114;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi = {loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo = {loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_115 = {v0_233, v0_232};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo_lo = _GEN_115;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo_lo = _GEN_115;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo_lo = _GEN_115;
  wire [63:0]         _GEN_116 = {v0_235, v0_234};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo_hi = _GEN_116;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo_hi = _GEN_116;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo_hi = _GEN_116;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo = {loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_117 = {v0_237, v0_236};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi_lo = _GEN_117;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi_lo = _GEN_117;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi_lo = _GEN_117;
  wire [63:0]         _GEN_118 = {v0_239, v0_238};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi_hi = _GEN_118;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi_hi = _GEN_118;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi_hi = _GEN_118;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi = {loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi = {loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo = {loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_119 = {v0_241, v0_240};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo_lo = _GEN_119;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo_lo = _GEN_119;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo_lo = _GEN_119;
  wire [63:0]         _GEN_120 = {v0_243, v0_242};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo_hi = _GEN_120;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo_hi = _GEN_120;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo_hi = _GEN_120;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo = {loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_121 = {v0_245, v0_244};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi_lo = _GEN_121;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi_lo = _GEN_121;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi_lo = _GEN_121;
  wire [63:0]         _GEN_122 = {v0_247, v0_246};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi_hi = _GEN_122;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi_hi = _GEN_122;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi_hi = _GEN_122;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi = {loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo = {loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_123 = {v0_249, v0_248};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo_lo = _GEN_123;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo_lo = _GEN_123;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo_lo = _GEN_123;
  wire [63:0]         _GEN_124 = {v0_251, v0_250};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo_hi = _GEN_124;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo_hi = _GEN_124;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo_hi = _GEN_124;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo = {loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_125 = {v0_253, v0_252};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi_lo = _GEN_125;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi_lo = _GEN_125;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi_lo = _GEN_125;
  wire [63:0]         _GEN_126 = {v0_255, v0_254};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi_hi = _GEN_126;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi_hi = _GEN_126;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi_hi = _GEN_126;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi = {loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi = {loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi = {loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_lo_lo_hi_hi_hi = {loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo};
  wire [2047:0]       loadUnit_maskInput_lo_lo_lo_hi_hi = {loadUnit_maskInput_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_lo};
  wire [4095:0]       loadUnit_maskInput_lo_lo_lo_hi = {loadUnit_maskInput_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_lo};
  wire [8191:0]       loadUnit_maskInput_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo};
  wire [63:0]         _GEN_127 = {v0_257, v0_256};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo_lo = _GEN_127;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo_lo = _GEN_127;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo_lo = _GEN_127;
  wire [63:0]         _GEN_128 = {v0_259, v0_258};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo_hi = _GEN_128;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo_hi = _GEN_128;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo_hi = _GEN_128;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo = {loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_129 = {v0_261, v0_260};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi_lo = _GEN_129;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi_lo = _GEN_129;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi_lo = _GEN_129;
  wire [63:0]         _GEN_130 = {v0_263, v0_262};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi_hi = _GEN_130;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi_hi = _GEN_130;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi_hi = _GEN_130;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi = {loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo = {loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_131 = {v0_265, v0_264};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo_lo = _GEN_131;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo_lo = _GEN_131;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo_lo = _GEN_131;
  wire [63:0]         _GEN_132 = {v0_267, v0_266};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo_hi = _GEN_132;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo_hi = _GEN_132;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo_hi = _GEN_132;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo = {loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_133 = {v0_269, v0_268};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi_lo = _GEN_133;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi_lo = _GEN_133;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi_lo = _GEN_133;
  wire [63:0]         _GEN_134 = {v0_271, v0_270};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi_hi = _GEN_134;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi_hi = _GEN_134;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi_hi = _GEN_134;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi = {loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi = {loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo = {loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_135 = {v0_273, v0_272};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo_lo = _GEN_135;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo_lo = _GEN_135;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo_lo = _GEN_135;
  wire [63:0]         _GEN_136 = {v0_275, v0_274};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo_hi = _GEN_136;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo_hi = _GEN_136;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo_hi = _GEN_136;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo = {loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_137 = {v0_277, v0_276};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi_lo = _GEN_137;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi_lo = _GEN_137;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi_lo = _GEN_137;
  wire [63:0]         _GEN_138 = {v0_279, v0_278};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi_hi = _GEN_138;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi_hi = _GEN_138;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi_hi = _GEN_138;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi = {loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo = {loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_139 = {v0_281, v0_280};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo_lo = _GEN_139;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo_lo = _GEN_139;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo_lo = _GEN_139;
  wire [63:0]         _GEN_140 = {v0_283, v0_282};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo_hi = _GEN_140;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo_hi = _GEN_140;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo_hi = _GEN_140;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo = {loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_141 = {v0_285, v0_284};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi_lo = _GEN_141;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi_lo = _GEN_141;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi_lo = _GEN_141;
  wire [63:0]         _GEN_142 = {v0_287, v0_286};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi_hi = _GEN_142;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi_hi = _GEN_142;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi_hi = _GEN_142;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi = {loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi = {loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi = {loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_lo_hi_lo_lo_lo = {loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_143 = {v0_289, v0_288};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo_lo = _GEN_143;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo_lo = _GEN_143;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo_lo = _GEN_143;
  wire [63:0]         _GEN_144 = {v0_291, v0_290};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo_hi = _GEN_144;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo_hi = _GEN_144;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo_hi = _GEN_144;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo = {loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_145 = {v0_293, v0_292};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi_lo = _GEN_145;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi_lo = _GEN_145;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi_lo = _GEN_145;
  wire [63:0]         _GEN_146 = {v0_295, v0_294};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi_hi = _GEN_146;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi_hi = _GEN_146;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi_hi = _GEN_146;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi = {loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo = {loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_147 = {v0_297, v0_296};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo_lo = _GEN_147;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo_lo = _GEN_147;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo_lo = _GEN_147;
  wire [63:0]         _GEN_148 = {v0_299, v0_298};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo_hi = _GEN_148;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo_hi = _GEN_148;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo_hi = _GEN_148;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo = {loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_149 = {v0_301, v0_300};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi_lo = _GEN_149;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi_lo = _GEN_149;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi_lo = _GEN_149;
  wire [63:0]         _GEN_150 = {v0_303, v0_302};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi_hi = _GEN_150;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi_hi = _GEN_150;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi_hi = _GEN_150;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi = {loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi = {loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo = {loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_151 = {v0_305, v0_304};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo_lo = _GEN_151;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo_lo = _GEN_151;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo_lo = _GEN_151;
  wire [63:0]         _GEN_152 = {v0_307, v0_306};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo_hi = _GEN_152;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo_hi = _GEN_152;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo_hi = _GEN_152;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo = {loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_153 = {v0_309, v0_308};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi_lo = _GEN_153;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi_lo = _GEN_153;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi_lo = _GEN_153;
  wire [63:0]         _GEN_154 = {v0_311, v0_310};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi_hi = _GEN_154;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi_hi = _GEN_154;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi_hi = _GEN_154;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi = {loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo = {loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_155 = {v0_313, v0_312};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo_lo = _GEN_155;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo_lo = _GEN_155;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo_lo = _GEN_155;
  wire [63:0]         _GEN_156 = {v0_315, v0_314};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo_hi = _GEN_156;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo_hi = _GEN_156;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo_hi = _GEN_156;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo = {loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_157 = {v0_317, v0_316};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi_lo = _GEN_157;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi_lo = _GEN_157;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi_lo = _GEN_157;
  wire [63:0]         _GEN_158 = {v0_319, v0_318};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi_hi = _GEN_158;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi_hi = _GEN_158;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi_hi = _GEN_158;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi = {loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi = {loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi = {loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_lo_hi_lo_lo_hi = {loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo};
  wire [2047:0]       loadUnit_maskInput_lo_lo_hi_lo_lo = {loadUnit_maskInput_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_159 = {v0_321, v0_320};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo_lo = _GEN_159;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo_lo = _GEN_159;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo_lo = _GEN_159;
  wire [63:0]         _GEN_160 = {v0_323, v0_322};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo_hi = _GEN_160;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo_hi = _GEN_160;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo_hi = _GEN_160;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo = {loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_161 = {v0_325, v0_324};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi_lo = _GEN_161;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi_lo = _GEN_161;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi_lo = _GEN_161;
  wire [63:0]         _GEN_162 = {v0_327, v0_326};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi_hi = _GEN_162;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi_hi = _GEN_162;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi_hi = _GEN_162;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi = {loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo = {loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_163 = {v0_329, v0_328};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo_lo = _GEN_163;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo_lo = _GEN_163;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo_lo = _GEN_163;
  wire [63:0]         _GEN_164 = {v0_331, v0_330};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo_hi = _GEN_164;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo_hi = _GEN_164;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo_hi = _GEN_164;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo = {loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_165 = {v0_333, v0_332};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi_lo = _GEN_165;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi_lo = _GEN_165;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi_lo = _GEN_165;
  wire [63:0]         _GEN_166 = {v0_335, v0_334};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi_hi = _GEN_166;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi_hi = _GEN_166;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi_hi = _GEN_166;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi = {loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi = {loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo = {loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_167 = {v0_337, v0_336};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo_lo = _GEN_167;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo_lo = _GEN_167;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo_lo = _GEN_167;
  wire [63:0]         _GEN_168 = {v0_339, v0_338};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo_hi = _GEN_168;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo_hi = _GEN_168;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo_hi = _GEN_168;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo = {loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_169 = {v0_341, v0_340};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi_lo = _GEN_169;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi_lo = _GEN_169;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi_lo = _GEN_169;
  wire [63:0]         _GEN_170 = {v0_343, v0_342};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi_hi = _GEN_170;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi_hi = _GEN_170;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi_hi = _GEN_170;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi = {loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo = {loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_171 = {v0_345, v0_344};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo_lo = _GEN_171;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo_lo = _GEN_171;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo_lo = _GEN_171;
  wire [63:0]         _GEN_172 = {v0_347, v0_346};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo_hi = _GEN_172;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo_hi = _GEN_172;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo_hi = _GEN_172;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo = {loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_173 = {v0_349, v0_348};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi_lo = _GEN_173;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi_lo = _GEN_173;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi_lo = _GEN_173;
  wire [63:0]         _GEN_174 = {v0_351, v0_350};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi_hi = _GEN_174;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi_hi = _GEN_174;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi_hi = _GEN_174;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi = {loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi = {loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi = {loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_lo_hi_lo_hi_lo = {loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_175 = {v0_353, v0_352};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo_lo = _GEN_175;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo_lo = _GEN_175;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo_lo = _GEN_175;
  wire [63:0]         _GEN_176 = {v0_355, v0_354};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo_hi = _GEN_176;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo_hi = _GEN_176;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo_hi = _GEN_176;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo = {loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_177 = {v0_357, v0_356};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi_lo = _GEN_177;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi_lo = _GEN_177;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi_lo = _GEN_177;
  wire [63:0]         _GEN_178 = {v0_359, v0_358};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi_hi = _GEN_178;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi_hi = _GEN_178;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi_hi = _GEN_178;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi = {loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo = {loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_179 = {v0_361, v0_360};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo_lo = _GEN_179;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo_lo = _GEN_179;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo_lo = _GEN_179;
  wire [63:0]         _GEN_180 = {v0_363, v0_362};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo_hi = _GEN_180;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo_hi = _GEN_180;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo_hi = _GEN_180;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo = {loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_181 = {v0_365, v0_364};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi_lo = _GEN_181;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi_lo = _GEN_181;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi_lo = _GEN_181;
  wire [63:0]         _GEN_182 = {v0_367, v0_366};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi_hi = _GEN_182;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi_hi = _GEN_182;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi_hi = _GEN_182;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi = {loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi = {loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo = {loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_183 = {v0_369, v0_368};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo_lo = _GEN_183;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo_lo = _GEN_183;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo_lo = _GEN_183;
  wire [63:0]         _GEN_184 = {v0_371, v0_370};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo_hi = _GEN_184;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo_hi = _GEN_184;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo_hi = _GEN_184;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo = {loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_185 = {v0_373, v0_372};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi_lo = _GEN_185;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi_lo = _GEN_185;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi_lo = _GEN_185;
  wire [63:0]         _GEN_186 = {v0_375, v0_374};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi_hi = _GEN_186;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi_hi = _GEN_186;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi_hi = _GEN_186;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi = {loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo = {loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_187 = {v0_377, v0_376};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo_lo = _GEN_187;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo_lo = _GEN_187;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo_lo = _GEN_187;
  wire [63:0]         _GEN_188 = {v0_379, v0_378};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo_hi = _GEN_188;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo_hi = _GEN_188;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo_hi = _GEN_188;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo = {loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_189 = {v0_381, v0_380};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi_lo = _GEN_189;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi_lo = _GEN_189;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi_lo = _GEN_189;
  wire [63:0]         _GEN_190 = {v0_383, v0_382};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi_hi = _GEN_190;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi_hi = _GEN_190;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi_hi = _GEN_190;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi = {loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi = {loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi = {loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_lo_hi_lo_hi_hi = {loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo};
  wire [2047:0]       loadUnit_maskInput_lo_lo_hi_lo_hi = {loadUnit_maskInput_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_lo};
  wire [4095:0]       loadUnit_maskInput_lo_lo_hi_lo = {loadUnit_maskInput_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_191 = {v0_385, v0_384};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo_lo = _GEN_191;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo_lo = _GEN_191;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo_lo = _GEN_191;
  wire [63:0]         _GEN_192 = {v0_387, v0_386};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo_hi = _GEN_192;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo_hi = _GEN_192;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo_hi = _GEN_192;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo = {loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_193 = {v0_389, v0_388};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi_lo = _GEN_193;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi_lo = _GEN_193;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi_lo = _GEN_193;
  wire [63:0]         _GEN_194 = {v0_391, v0_390};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi_hi = _GEN_194;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi_hi = _GEN_194;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi_hi = _GEN_194;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi = {loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo = {loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_195 = {v0_393, v0_392};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo_lo = _GEN_195;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo_lo = _GEN_195;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo_lo = _GEN_195;
  wire [63:0]         _GEN_196 = {v0_395, v0_394};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo_hi = _GEN_196;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo_hi = _GEN_196;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo_hi = _GEN_196;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo = {loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_197 = {v0_397, v0_396};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi_lo = _GEN_197;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi_lo = _GEN_197;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi_lo = _GEN_197;
  wire [63:0]         _GEN_198 = {v0_399, v0_398};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi_hi = _GEN_198;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi_hi = _GEN_198;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi_hi = _GEN_198;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi = {loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi = {loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo = {loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_199 = {v0_401, v0_400};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo_lo = _GEN_199;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo_lo = _GEN_199;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo_lo = _GEN_199;
  wire [63:0]         _GEN_200 = {v0_403, v0_402};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo_hi = _GEN_200;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo_hi = _GEN_200;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo_hi = _GEN_200;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo = {loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_201 = {v0_405, v0_404};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi_lo = _GEN_201;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi_lo = _GEN_201;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi_lo = _GEN_201;
  wire [63:0]         _GEN_202 = {v0_407, v0_406};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi_hi = _GEN_202;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi_hi = _GEN_202;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi_hi = _GEN_202;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi = {loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo = {loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_203 = {v0_409, v0_408};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo_lo = _GEN_203;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo_lo = _GEN_203;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo_lo = _GEN_203;
  wire [63:0]         _GEN_204 = {v0_411, v0_410};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo_hi = _GEN_204;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo_hi = _GEN_204;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo_hi = _GEN_204;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo = {loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_205 = {v0_413, v0_412};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi_lo = _GEN_205;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi_lo = _GEN_205;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi_lo = _GEN_205;
  wire [63:0]         _GEN_206 = {v0_415, v0_414};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi_hi = _GEN_206;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi_hi = _GEN_206;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi_hi = _GEN_206;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi = {loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi = {loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi = {loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_lo_hi_hi_lo_lo = {loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_207 = {v0_417, v0_416};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo_lo = _GEN_207;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo_lo = _GEN_207;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo_lo = _GEN_207;
  wire [63:0]         _GEN_208 = {v0_419, v0_418};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo_hi = _GEN_208;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo_hi = _GEN_208;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo_hi = _GEN_208;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo = {loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_209 = {v0_421, v0_420};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi_lo = _GEN_209;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi_lo = _GEN_209;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi_lo = _GEN_209;
  wire [63:0]         _GEN_210 = {v0_423, v0_422};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi_hi = _GEN_210;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi_hi = _GEN_210;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi_hi = _GEN_210;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi = {loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo = {loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_211 = {v0_425, v0_424};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo_lo = _GEN_211;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo_lo = _GEN_211;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo_lo = _GEN_211;
  wire [63:0]         _GEN_212 = {v0_427, v0_426};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo_hi = _GEN_212;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo_hi = _GEN_212;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo_hi = _GEN_212;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo = {loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_213 = {v0_429, v0_428};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi_lo = _GEN_213;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi_lo = _GEN_213;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi_lo = _GEN_213;
  wire [63:0]         _GEN_214 = {v0_431, v0_430};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi_hi = _GEN_214;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi_hi = _GEN_214;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi_hi = _GEN_214;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi = {loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi = {loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo = {loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_215 = {v0_433, v0_432};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo_lo = _GEN_215;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo_lo = _GEN_215;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo_lo = _GEN_215;
  wire [63:0]         _GEN_216 = {v0_435, v0_434};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo_hi = _GEN_216;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo_hi = _GEN_216;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo_hi = _GEN_216;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo = {loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_217 = {v0_437, v0_436};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi_lo = _GEN_217;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi_lo = _GEN_217;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi_lo = _GEN_217;
  wire [63:0]         _GEN_218 = {v0_439, v0_438};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi_hi = _GEN_218;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi_hi = _GEN_218;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi_hi = _GEN_218;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi = {loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo = {loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_219 = {v0_441, v0_440};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo_lo = _GEN_219;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo_lo = _GEN_219;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo_lo = _GEN_219;
  wire [63:0]         _GEN_220 = {v0_443, v0_442};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo_hi = _GEN_220;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo_hi = _GEN_220;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo_hi = _GEN_220;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo = {loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_221 = {v0_445, v0_444};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi_lo = _GEN_221;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi_lo = _GEN_221;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi_lo = _GEN_221;
  wire [63:0]         _GEN_222 = {v0_447, v0_446};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi_hi = _GEN_222;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi_hi = _GEN_222;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi_hi = _GEN_222;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi = {loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi = {loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi = {loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_lo_hi_hi_lo_hi = {loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo};
  wire [2047:0]       loadUnit_maskInput_lo_lo_hi_hi_lo = {loadUnit_maskInput_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_223 = {v0_449, v0_448};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo_lo = _GEN_223;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo_lo = _GEN_223;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo_lo = _GEN_223;
  wire [63:0]         _GEN_224 = {v0_451, v0_450};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo_hi = _GEN_224;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo_hi = _GEN_224;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo_hi = _GEN_224;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo = {loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_225 = {v0_453, v0_452};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi_lo = _GEN_225;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi_lo = _GEN_225;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi_lo = _GEN_225;
  wire [63:0]         _GEN_226 = {v0_455, v0_454};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi_hi = _GEN_226;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi_hi = _GEN_226;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi_hi = _GEN_226;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi = {loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo = {loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_227 = {v0_457, v0_456};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo_lo = _GEN_227;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo_lo = _GEN_227;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo_lo = _GEN_227;
  wire [63:0]         _GEN_228 = {v0_459, v0_458};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo_hi = _GEN_228;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo_hi = _GEN_228;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo_hi = _GEN_228;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo = {loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_229 = {v0_461, v0_460};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi_lo = _GEN_229;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi_lo = _GEN_229;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi_lo = _GEN_229;
  wire [63:0]         _GEN_230 = {v0_463, v0_462};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi_hi = _GEN_230;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi_hi = _GEN_230;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi_hi = _GEN_230;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi = {loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi = {loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo = {loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_231 = {v0_465, v0_464};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo_lo = _GEN_231;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo_lo = _GEN_231;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo_lo = _GEN_231;
  wire [63:0]         _GEN_232 = {v0_467, v0_466};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo_hi = _GEN_232;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo_hi = _GEN_232;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo_hi = _GEN_232;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo = {loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_233 = {v0_469, v0_468};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi_lo = _GEN_233;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi_lo = _GEN_233;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi_lo = _GEN_233;
  wire [63:0]         _GEN_234 = {v0_471, v0_470};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi_hi = _GEN_234;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi_hi = _GEN_234;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi_hi = _GEN_234;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi = {loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo = {loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_235 = {v0_473, v0_472};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo_lo = _GEN_235;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo_lo = _GEN_235;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo_lo = _GEN_235;
  wire [63:0]         _GEN_236 = {v0_475, v0_474};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo_hi = _GEN_236;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo_hi = _GEN_236;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo_hi = _GEN_236;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo = {loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_237 = {v0_477, v0_476};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi_lo = _GEN_237;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi_lo = _GEN_237;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi_lo = _GEN_237;
  wire [63:0]         _GEN_238 = {v0_479, v0_478};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi_hi = _GEN_238;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi_hi = _GEN_238;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi_hi = _GEN_238;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi = {loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi = {loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi = {loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_lo_hi_hi_hi_lo = {loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_239 = {v0_481, v0_480};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo_lo = _GEN_239;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo_lo = _GEN_239;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo_lo = _GEN_239;
  wire [63:0]         _GEN_240 = {v0_483, v0_482};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo_hi = _GEN_240;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo_hi = _GEN_240;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo_hi = _GEN_240;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo = {loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_241 = {v0_485, v0_484};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi_lo = _GEN_241;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi_lo = _GEN_241;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi_lo = _GEN_241;
  wire [63:0]         _GEN_242 = {v0_487, v0_486};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi_hi = _GEN_242;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi_hi = _GEN_242;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi_hi = _GEN_242;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi = {loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo = {loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_243 = {v0_489, v0_488};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo_lo = _GEN_243;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo_lo = _GEN_243;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo_lo = _GEN_243;
  wire [63:0]         _GEN_244 = {v0_491, v0_490};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo_hi = _GEN_244;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo_hi = _GEN_244;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo_hi = _GEN_244;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo = {loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_245 = {v0_493, v0_492};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi_lo = _GEN_245;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi_lo = _GEN_245;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi_lo = _GEN_245;
  wire [63:0]         _GEN_246 = {v0_495, v0_494};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi_hi = _GEN_246;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi_hi = _GEN_246;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi_hi = _GEN_246;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi = {loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi = {loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo = {loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_247 = {v0_497, v0_496};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo_lo = _GEN_247;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo_lo = _GEN_247;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo_lo = _GEN_247;
  wire [63:0]         _GEN_248 = {v0_499, v0_498};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo_hi = _GEN_248;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo_hi = _GEN_248;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo_hi = _GEN_248;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo = {loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_249 = {v0_501, v0_500};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi_lo = _GEN_249;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi_lo = _GEN_249;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi_lo = _GEN_249;
  wire [63:0]         _GEN_250 = {v0_503, v0_502};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi_hi = _GEN_250;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi_hi = _GEN_250;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi_hi = _GEN_250;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi = {loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo = {loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_251 = {v0_505, v0_504};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo_lo = _GEN_251;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo_lo = _GEN_251;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo_lo = _GEN_251;
  wire [63:0]         _GEN_252 = {v0_507, v0_506};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo_hi = _GEN_252;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo_hi = _GEN_252;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo_hi = _GEN_252;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo = {loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_253 = {v0_509, v0_508};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi_lo = _GEN_253;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi_lo = _GEN_253;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi_lo = _GEN_253;
  wire [63:0]         _GEN_254 = {v0_511, v0_510};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi_hi = _GEN_254;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi_hi = _GEN_254;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi_hi = _GEN_254;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi = {loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi = {loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi = {loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_lo_hi_hi_hi_hi = {loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo};
  wire [2047:0]       loadUnit_maskInput_lo_lo_hi_hi_hi = {loadUnit_maskInput_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_lo};
  wire [4095:0]       loadUnit_maskInput_lo_lo_hi_hi = {loadUnit_maskInput_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_lo};
  wire [8191:0]       loadUnit_maskInput_lo_lo_hi = {loadUnit_maskInput_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo};
  wire [16383:0]      loadUnit_maskInput_lo_lo = {loadUnit_maskInput_lo_lo_hi, loadUnit_maskInput_lo_lo_lo};
  wire [63:0]         _GEN_255 = {v0_513, v0_512};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo_lo = _GEN_255;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo_lo = _GEN_255;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo_lo = _GEN_255;
  wire [63:0]         _GEN_256 = {v0_515, v0_514};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo_hi = _GEN_256;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo_hi = _GEN_256;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo_hi = _GEN_256;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo = {loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_257 = {v0_517, v0_516};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi_lo = _GEN_257;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi_lo = _GEN_257;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi_lo = _GEN_257;
  wire [63:0]         _GEN_258 = {v0_519, v0_518};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi_hi = _GEN_258;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi_hi = _GEN_258;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi_hi = _GEN_258;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi = {loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo = {loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_259 = {v0_521, v0_520};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo_lo = _GEN_259;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo_lo = _GEN_259;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo_lo = _GEN_259;
  wire [63:0]         _GEN_260 = {v0_523, v0_522};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo_hi = _GEN_260;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo_hi = _GEN_260;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo_hi = _GEN_260;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_261 = {v0_525, v0_524};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi_lo = _GEN_261;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi_lo = _GEN_261;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi_lo = _GEN_261;
  wire [63:0]         _GEN_262 = {v0_527, v0_526};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi_hi = _GEN_262;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi_hi = _GEN_262;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi_hi = _GEN_262;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi = {loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi = {loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo = {loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_263 = {v0_529, v0_528};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo_lo = _GEN_263;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo_lo = _GEN_263;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo_lo = _GEN_263;
  wire [63:0]         _GEN_264 = {v0_531, v0_530};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo_hi = _GEN_264;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo_hi = _GEN_264;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo_hi = _GEN_264;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo = {loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_265 = {v0_533, v0_532};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi_lo = _GEN_265;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi_lo = _GEN_265;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi_lo = _GEN_265;
  wire [63:0]         _GEN_266 = {v0_535, v0_534};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi_hi = _GEN_266;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi_hi = _GEN_266;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi_hi = _GEN_266;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi = {loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_267 = {v0_537, v0_536};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo_lo = _GEN_267;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo_lo = _GEN_267;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo_lo = _GEN_267;
  wire [63:0]         _GEN_268 = {v0_539, v0_538};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo_hi = _GEN_268;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo_hi = _GEN_268;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo_hi = _GEN_268;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo = {loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_269 = {v0_541, v0_540};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi_lo = _GEN_269;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi_lo = _GEN_269;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi_lo = _GEN_269;
  wire [63:0]         _GEN_270 = {v0_543, v0_542};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi_hi = _GEN_270;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi_hi = _GEN_270;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi_hi = _GEN_270;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi = {loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi = {loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi = {loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_hi_lo_lo_lo_lo = {loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_271 = {v0_545, v0_544};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo_lo = _GEN_271;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo_lo = _GEN_271;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo_lo = _GEN_271;
  wire [63:0]         _GEN_272 = {v0_547, v0_546};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo_hi = _GEN_272;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo_hi = _GEN_272;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo_hi = _GEN_272;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo = {loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_273 = {v0_549, v0_548};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi_lo = _GEN_273;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi_lo = _GEN_273;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi_lo = _GEN_273;
  wire [63:0]         _GEN_274 = {v0_551, v0_550};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi_hi = _GEN_274;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi_hi = _GEN_274;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi_hi = _GEN_274;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi = {loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo = {loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_275 = {v0_553, v0_552};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo_lo = _GEN_275;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo_lo = _GEN_275;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo_lo = _GEN_275;
  wire [63:0]         _GEN_276 = {v0_555, v0_554};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo_hi = _GEN_276;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo_hi = _GEN_276;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo_hi = _GEN_276;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_277 = {v0_557, v0_556};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi_lo = _GEN_277;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi_lo = _GEN_277;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi_lo = _GEN_277;
  wire [63:0]         _GEN_278 = {v0_559, v0_558};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi_hi = _GEN_278;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi_hi = _GEN_278;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi_hi = _GEN_278;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi = {loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi = {loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_279 = {v0_561, v0_560};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo_lo = _GEN_279;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo_lo = _GEN_279;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo_lo = _GEN_279;
  wire [63:0]         _GEN_280 = {v0_563, v0_562};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo_hi = _GEN_280;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo_hi = _GEN_280;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo_hi = _GEN_280;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo = {loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_281 = {v0_565, v0_564};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi_lo = _GEN_281;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi_lo = _GEN_281;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi_lo = _GEN_281;
  wire [63:0]         _GEN_282 = {v0_567, v0_566};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi_hi = _GEN_282;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi_hi = _GEN_282;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi_hi = _GEN_282;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi = {loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo = {loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_283 = {v0_569, v0_568};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo_lo = _GEN_283;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo_lo = _GEN_283;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo_lo = _GEN_283;
  wire [63:0]         _GEN_284 = {v0_571, v0_570};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo_hi = _GEN_284;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo_hi = _GEN_284;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo_hi = _GEN_284;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo = {loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_285 = {v0_573, v0_572};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi_lo = _GEN_285;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi_lo = _GEN_285;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi_lo = _GEN_285;
  wire [63:0]         _GEN_286 = {v0_575, v0_574};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi_hi = _GEN_286;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi_hi = _GEN_286;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi_hi = _GEN_286;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi = {loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi = {loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi = {loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_hi_lo_lo_lo_hi = {loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo};
  wire [2047:0]       loadUnit_maskInput_lo_hi_lo_lo_lo = {loadUnit_maskInput_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_287 = {v0_577, v0_576};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo_lo = _GEN_287;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo_lo = _GEN_287;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo_lo = _GEN_287;
  wire [63:0]         _GEN_288 = {v0_579, v0_578};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo_hi = _GEN_288;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo_hi = _GEN_288;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo_hi = _GEN_288;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo = {loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_289 = {v0_581, v0_580};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi_lo = _GEN_289;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi_lo = _GEN_289;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi_lo = _GEN_289;
  wire [63:0]         _GEN_290 = {v0_583, v0_582};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi_hi = _GEN_290;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi_hi = _GEN_290;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi_hi = _GEN_290;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi = {loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo = {loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_291 = {v0_585, v0_584};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo_lo = _GEN_291;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo_lo = _GEN_291;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo_lo = _GEN_291;
  wire [63:0]         _GEN_292 = {v0_587, v0_586};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo_hi = _GEN_292;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo_hi = _GEN_292;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo_hi = _GEN_292;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_293 = {v0_589, v0_588};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi_lo = _GEN_293;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi_lo = _GEN_293;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi_lo = _GEN_293;
  wire [63:0]         _GEN_294 = {v0_591, v0_590};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi_hi = _GEN_294;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi_hi = _GEN_294;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi_hi = _GEN_294;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi = {loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi = {loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo = {loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_295 = {v0_593, v0_592};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo_lo = _GEN_295;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo_lo = _GEN_295;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo_lo = _GEN_295;
  wire [63:0]         _GEN_296 = {v0_595, v0_594};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo_hi = _GEN_296;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo_hi = _GEN_296;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo_hi = _GEN_296;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo = {loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_297 = {v0_597, v0_596};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi_lo = _GEN_297;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi_lo = _GEN_297;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi_lo = _GEN_297;
  wire [63:0]         _GEN_298 = {v0_599, v0_598};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi_hi = _GEN_298;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi_hi = _GEN_298;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi_hi = _GEN_298;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi = {loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_299 = {v0_601, v0_600};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo_lo = _GEN_299;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo_lo = _GEN_299;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo_lo = _GEN_299;
  wire [63:0]         _GEN_300 = {v0_603, v0_602};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo_hi = _GEN_300;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo_hi = _GEN_300;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo_hi = _GEN_300;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo = {loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_301 = {v0_605, v0_604};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi_lo = _GEN_301;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi_lo = _GEN_301;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi_lo = _GEN_301;
  wire [63:0]         _GEN_302 = {v0_607, v0_606};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi_hi = _GEN_302;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi_hi = _GEN_302;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi_hi = _GEN_302;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi = {loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi = {loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi = {loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_hi_lo_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_303 = {v0_609, v0_608};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo_lo = _GEN_303;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo_lo = _GEN_303;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo_lo = _GEN_303;
  wire [63:0]         _GEN_304 = {v0_611, v0_610};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo_hi = _GEN_304;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo_hi = _GEN_304;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo_hi = _GEN_304;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo = {loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_305 = {v0_613, v0_612};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi_lo = _GEN_305;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi_lo = _GEN_305;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi_lo = _GEN_305;
  wire [63:0]         _GEN_306 = {v0_615, v0_614};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi_hi = _GEN_306;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi_hi = _GEN_306;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi_hi = _GEN_306;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi = {loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo = {loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_307 = {v0_617, v0_616};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo_lo = _GEN_307;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo_lo = _GEN_307;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo_lo = _GEN_307;
  wire [63:0]         _GEN_308 = {v0_619, v0_618};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo_hi = _GEN_308;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo_hi = _GEN_308;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo_hi = _GEN_308;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_309 = {v0_621, v0_620};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi_lo = _GEN_309;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi_lo = _GEN_309;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi_lo = _GEN_309;
  wire [63:0]         _GEN_310 = {v0_623, v0_622};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi_hi = _GEN_310;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi_hi = _GEN_310;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi_hi = _GEN_310;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi = {loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi = {loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo = {loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_311 = {v0_625, v0_624};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo_lo = _GEN_311;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo_lo = _GEN_311;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo_lo = _GEN_311;
  wire [63:0]         _GEN_312 = {v0_627, v0_626};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo_hi = _GEN_312;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo_hi = _GEN_312;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo_hi = _GEN_312;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo = {loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_313 = {v0_629, v0_628};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi_lo = _GEN_313;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi_lo = _GEN_313;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi_lo = _GEN_313;
  wire [63:0]         _GEN_314 = {v0_631, v0_630};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi_hi = _GEN_314;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi_hi = _GEN_314;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi_hi = _GEN_314;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi = {loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo = {loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_315 = {v0_633, v0_632};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo_lo = _GEN_315;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo_lo = _GEN_315;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo_lo = _GEN_315;
  wire [63:0]         _GEN_316 = {v0_635, v0_634};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo_hi = _GEN_316;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo_hi = _GEN_316;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo_hi = _GEN_316;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo = {loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_317 = {v0_637, v0_636};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi_lo = _GEN_317;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi_lo = _GEN_317;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi_lo = _GEN_317;
  wire [63:0]         _GEN_318 = {v0_639, v0_638};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi_hi = _GEN_318;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi_hi = _GEN_318;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi_hi = _GEN_318;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi = {loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi = {loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi = {loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_hi_lo_lo_hi_hi = {loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo};
  wire [2047:0]       loadUnit_maskInput_lo_hi_lo_lo_hi = {loadUnit_maskInput_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_lo};
  wire [4095:0]       loadUnit_maskInput_lo_hi_lo_lo = {loadUnit_maskInput_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_319 = {v0_641, v0_640};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo_lo = _GEN_319;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo_lo = _GEN_319;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo_lo = _GEN_319;
  wire [63:0]         _GEN_320 = {v0_643, v0_642};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo_hi = _GEN_320;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo_hi = _GEN_320;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo_hi = _GEN_320;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo = {loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_321 = {v0_645, v0_644};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi_lo = _GEN_321;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi_lo = _GEN_321;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi_lo = _GEN_321;
  wire [63:0]         _GEN_322 = {v0_647, v0_646};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi_hi = _GEN_322;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi_hi = _GEN_322;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi_hi = _GEN_322;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi = {loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo = {loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_323 = {v0_649, v0_648};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo_lo = _GEN_323;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo_lo = _GEN_323;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo_lo = _GEN_323;
  wire [63:0]         _GEN_324 = {v0_651, v0_650};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo_hi = _GEN_324;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo_hi = _GEN_324;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo_hi = _GEN_324;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_325 = {v0_653, v0_652};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi_lo = _GEN_325;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi_lo = _GEN_325;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi_lo = _GEN_325;
  wire [63:0]         _GEN_326 = {v0_655, v0_654};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi_hi = _GEN_326;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi_hi = _GEN_326;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi_hi = _GEN_326;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi = {loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi = {loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo = {loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_327 = {v0_657, v0_656};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo_lo = _GEN_327;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo_lo = _GEN_327;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo_lo = _GEN_327;
  wire [63:0]         _GEN_328 = {v0_659, v0_658};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo_hi = _GEN_328;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo_hi = _GEN_328;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo_hi = _GEN_328;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo = {loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_329 = {v0_661, v0_660};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi_lo = _GEN_329;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi_lo = _GEN_329;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi_lo = _GEN_329;
  wire [63:0]         _GEN_330 = {v0_663, v0_662};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi_hi = _GEN_330;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi_hi = _GEN_330;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi_hi = _GEN_330;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi = {loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_331 = {v0_665, v0_664};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo_lo = _GEN_331;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo_lo = _GEN_331;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo_lo = _GEN_331;
  wire [63:0]         _GEN_332 = {v0_667, v0_666};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo_hi = _GEN_332;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo_hi = _GEN_332;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo_hi = _GEN_332;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_333 = {v0_669, v0_668};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi_lo = _GEN_333;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi_lo = _GEN_333;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi_lo = _GEN_333;
  wire [63:0]         _GEN_334 = {v0_671, v0_670};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi_hi = _GEN_334;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi_hi = _GEN_334;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi_hi = _GEN_334;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi = {loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi = {loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi = {loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_hi_lo_hi_lo_lo = {loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_335 = {v0_673, v0_672};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo_lo = _GEN_335;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo_lo = _GEN_335;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo_lo = _GEN_335;
  wire [63:0]         _GEN_336 = {v0_675, v0_674};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo_hi = _GEN_336;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo_hi = _GEN_336;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo_hi = _GEN_336;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo = {loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_337 = {v0_677, v0_676};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi_lo = _GEN_337;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi_lo = _GEN_337;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi_lo = _GEN_337;
  wire [63:0]         _GEN_338 = {v0_679, v0_678};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi_hi = _GEN_338;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi_hi = _GEN_338;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi_hi = _GEN_338;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi = {loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo = {loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_339 = {v0_681, v0_680};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo_lo = _GEN_339;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo_lo = _GEN_339;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo_lo = _GEN_339;
  wire [63:0]         _GEN_340 = {v0_683, v0_682};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo_hi = _GEN_340;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo_hi = _GEN_340;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo_hi = _GEN_340;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_341 = {v0_685, v0_684};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi_lo = _GEN_341;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi_lo = _GEN_341;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi_lo = _GEN_341;
  wire [63:0]         _GEN_342 = {v0_687, v0_686};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi_hi = _GEN_342;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi_hi = _GEN_342;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi_hi = _GEN_342;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi = {loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi = {loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_343 = {v0_689, v0_688};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo_lo = _GEN_343;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo_lo = _GEN_343;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo_lo = _GEN_343;
  wire [63:0]         _GEN_344 = {v0_691, v0_690};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo_hi = _GEN_344;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo_hi = _GEN_344;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo_hi = _GEN_344;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo = {loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_345 = {v0_693, v0_692};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi_lo = _GEN_345;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi_lo = _GEN_345;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi_lo = _GEN_345;
  wire [63:0]         _GEN_346 = {v0_695, v0_694};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi_hi = _GEN_346;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi_hi = _GEN_346;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi_hi = _GEN_346;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi = {loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_347 = {v0_697, v0_696};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo_lo = _GEN_347;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo_lo = _GEN_347;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo_lo = _GEN_347;
  wire [63:0]         _GEN_348 = {v0_699, v0_698};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo_hi = _GEN_348;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo_hi = _GEN_348;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo_hi = _GEN_348;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_349 = {v0_701, v0_700};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi_lo = _GEN_349;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi_lo = _GEN_349;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi_lo = _GEN_349;
  wire [63:0]         _GEN_350 = {v0_703, v0_702};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi_hi = _GEN_350;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi_hi = _GEN_350;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi_hi = _GEN_350;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi = {loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi = {loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi = {loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_hi_lo_hi_lo_hi = {loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo};
  wire [2047:0]       loadUnit_maskInput_lo_hi_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_351 = {v0_705, v0_704};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo_lo = _GEN_351;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo_lo = _GEN_351;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo_lo = _GEN_351;
  wire [63:0]         _GEN_352 = {v0_707, v0_706};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo_hi = _GEN_352;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo_hi = _GEN_352;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo_hi = _GEN_352;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo = {loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_353 = {v0_709, v0_708};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi_lo = _GEN_353;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi_lo = _GEN_353;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi_lo = _GEN_353;
  wire [63:0]         _GEN_354 = {v0_711, v0_710};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi_hi = _GEN_354;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi_hi = _GEN_354;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi_hi = _GEN_354;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi = {loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo = {loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_355 = {v0_713, v0_712};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo_lo = _GEN_355;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo_lo = _GEN_355;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo_lo = _GEN_355;
  wire [63:0]         _GEN_356 = {v0_715, v0_714};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo_hi = _GEN_356;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo_hi = _GEN_356;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo_hi = _GEN_356;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_357 = {v0_717, v0_716};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi_lo = _GEN_357;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi_lo = _GEN_357;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi_lo = _GEN_357;
  wire [63:0]         _GEN_358 = {v0_719, v0_718};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi_hi = _GEN_358;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi_hi = _GEN_358;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi_hi = _GEN_358;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi = {loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi = {loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo = {loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_359 = {v0_721, v0_720};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo_lo = _GEN_359;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo_lo = _GEN_359;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo_lo = _GEN_359;
  wire [63:0]         _GEN_360 = {v0_723, v0_722};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo_hi = _GEN_360;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo_hi = _GEN_360;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo_hi = _GEN_360;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo = {loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_361 = {v0_725, v0_724};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi_lo = _GEN_361;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi_lo = _GEN_361;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi_lo = _GEN_361;
  wire [63:0]         _GEN_362 = {v0_727, v0_726};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi_hi = _GEN_362;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi_hi = _GEN_362;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi_hi = _GEN_362;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi = {loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_363 = {v0_729, v0_728};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo_lo = _GEN_363;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo_lo = _GEN_363;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo_lo = _GEN_363;
  wire [63:0]         _GEN_364 = {v0_731, v0_730};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo_hi = _GEN_364;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo_hi = _GEN_364;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo_hi = _GEN_364;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_365 = {v0_733, v0_732};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi_lo = _GEN_365;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi_lo = _GEN_365;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi_lo = _GEN_365;
  wire [63:0]         _GEN_366 = {v0_735, v0_734};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi_hi = _GEN_366;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi_hi = _GEN_366;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi_hi = _GEN_366;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi = {loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi = {loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi = {loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_hi_lo_hi_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_367 = {v0_737, v0_736};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo_lo = _GEN_367;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo_lo = _GEN_367;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo_lo = _GEN_367;
  wire [63:0]         _GEN_368 = {v0_739, v0_738};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo_hi = _GEN_368;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo_hi = _GEN_368;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo_hi = _GEN_368;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo = {loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_369 = {v0_741, v0_740};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi_lo = _GEN_369;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi_lo = _GEN_369;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi_lo = _GEN_369;
  wire [63:0]         _GEN_370 = {v0_743, v0_742};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi_hi = _GEN_370;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi_hi = _GEN_370;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi_hi = _GEN_370;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi = {loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo = {loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_371 = {v0_745, v0_744};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo_lo = _GEN_371;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo_lo = _GEN_371;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo_lo = _GEN_371;
  wire [63:0]         _GEN_372 = {v0_747, v0_746};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo_hi = _GEN_372;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo_hi = _GEN_372;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo_hi = _GEN_372;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_373 = {v0_749, v0_748};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi_lo = _GEN_373;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi_lo = _GEN_373;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi_lo = _GEN_373;
  wire [63:0]         _GEN_374 = {v0_751, v0_750};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi_hi = _GEN_374;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi_hi = _GEN_374;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi_hi = _GEN_374;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi = {loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi = {loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_375 = {v0_753, v0_752};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo_lo = _GEN_375;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo_lo = _GEN_375;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo_lo = _GEN_375;
  wire [63:0]         _GEN_376 = {v0_755, v0_754};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo_hi = _GEN_376;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo_hi = _GEN_376;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo_hi = _GEN_376;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo = {loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_377 = {v0_757, v0_756};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi_lo = _GEN_377;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi_lo = _GEN_377;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi_lo = _GEN_377;
  wire [63:0]         _GEN_378 = {v0_759, v0_758};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi_hi = _GEN_378;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi_hi = _GEN_378;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi_hi = _GEN_378;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi = {loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_379 = {v0_761, v0_760};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo_lo = _GEN_379;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo_lo = _GEN_379;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo_lo = _GEN_379;
  wire [63:0]         _GEN_380 = {v0_763, v0_762};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo_hi = _GEN_380;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo_hi = _GEN_380;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo_hi = _GEN_380;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_381 = {v0_765, v0_764};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi_lo = _GEN_381;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi_lo = _GEN_381;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi_lo = _GEN_381;
  wire [63:0]         _GEN_382 = {v0_767, v0_766};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi_hi = _GEN_382;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi_hi = _GEN_382;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi_hi = _GEN_382;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi = {loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi = {loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi = {loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_hi_lo_hi_hi_hi = {loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo};
  wire [2047:0]       loadUnit_maskInput_lo_hi_lo_hi_hi = {loadUnit_maskInput_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_lo};
  wire [4095:0]       loadUnit_maskInput_lo_hi_lo_hi = {loadUnit_maskInput_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_lo};
  wire [8191:0]       loadUnit_maskInput_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_lo};
  wire [63:0]         _GEN_383 = {v0_769, v0_768};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo_lo = _GEN_383;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo_lo = _GEN_383;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo_lo = _GEN_383;
  wire [63:0]         _GEN_384 = {v0_771, v0_770};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo_hi = _GEN_384;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo_hi = _GEN_384;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo_hi = _GEN_384;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo = {loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_385 = {v0_773, v0_772};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi_lo = _GEN_385;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi_lo = _GEN_385;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi_lo = _GEN_385;
  wire [63:0]         _GEN_386 = {v0_775, v0_774};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi_hi = _GEN_386;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi_hi = _GEN_386;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi_hi = _GEN_386;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi = {loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo = {loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_387 = {v0_777, v0_776};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo_lo = _GEN_387;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo_lo = _GEN_387;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo_lo = _GEN_387;
  wire [63:0]         _GEN_388 = {v0_779, v0_778};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo_hi = _GEN_388;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo_hi = _GEN_388;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo_hi = _GEN_388;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo = {loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_389 = {v0_781, v0_780};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi_lo = _GEN_389;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi_lo = _GEN_389;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi_lo = _GEN_389;
  wire [63:0]         _GEN_390 = {v0_783, v0_782};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi_hi = _GEN_390;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi_hi = _GEN_390;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi_hi = _GEN_390;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi = {loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi = {loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo = {loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_391 = {v0_785, v0_784};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo_lo = _GEN_391;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo_lo = _GEN_391;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo_lo = _GEN_391;
  wire [63:0]         _GEN_392 = {v0_787, v0_786};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo_hi = _GEN_392;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo_hi = _GEN_392;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo_hi = _GEN_392;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo = {loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_393 = {v0_789, v0_788};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi_lo = _GEN_393;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi_lo = _GEN_393;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi_lo = _GEN_393;
  wire [63:0]         _GEN_394 = {v0_791, v0_790};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi_hi = _GEN_394;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi_hi = _GEN_394;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi_hi = _GEN_394;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi = {loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo = {loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_395 = {v0_793, v0_792};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo_lo = _GEN_395;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo_lo = _GEN_395;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo_lo = _GEN_395;
  wire [63:0]         _GEN_396 = {v0_795, v0_794};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo_hi = _GEN_396;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo_hi = _GEN_396;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo_hi = _GEN_396;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo = {loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_397 = {v0_797, v0_796};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi_lo = _GEN_397;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi_lo = _GEN_397;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi_lo = _GEN_397;
  wire [63:0]         _GEN_398 = {v0_799, v0_798};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi_hi = _GEN_398;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi_hi = _GEN_398;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi_hi = _GEN_398;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi = {loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi = {loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi = {loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_hi_hi_lo_lo_lo = {loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_399 = {v0_801, v0_800};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo_lo = _GEN_399;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo_lo = _GEN_399;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo_lo = _GEN_399;
  wire [63:0]         _GEN_400 = {v0_803, v0_802};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo_hi = _GEN_400;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo_hi = _GEN_400;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo_hi = _GEN_400;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo = {loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_401 = {v0_805, v0_804};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi_lo = _GEN_401;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi_lo = _GEN_401;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi_lo = _GEN_401;
  wire [63:0]         _GEN_402 = {v0_807, v0_806};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi_hi = _GEN_402;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi_hi = _GEN_402;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi_hi = _GEN_402;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi = {loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo = {loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_403 = {v0_809, v0_808};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo_lo = _GEN_403;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo_lo = _GEN_403;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo_lo = _GEN_403;
  wire [63:0]         _GEN_404 = {v0_811, v0_810};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo_hi = _GEN_404;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo_hi = _GEN_404;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo_hi = _GEN_404;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo = {loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_405 = {v0_813, v0_812};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi_lo = _GEN_405;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi_lo = _GEN_405;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi_lo = _GEN_405;
  wire [63:0]         _GEN_406 = {v0_815, v0_814};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi_hi = _GEN_406;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi_hi = _GEN_406;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi_hi = _GEN_406;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi = {loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi = {loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo = {loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_407 = {v0_817, v0_816};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo_lo = _GEN_407;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo_lo = _GEN_407;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo_lo = _GEN_407;
  wire [63:0]         _GEN_408 = {v0_819, v0_818};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo_hi = _GEN_408;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo_hi = _GEN_408;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo_hi = _GEN_408;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo = {loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_409 = {v0_821, v0_820};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi_lo = _GEN_409;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi_lo = _GEN_409;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi_lo = _GEN_409;
  wire [63:0]         _GEN_410 = {v0_823, v0_822};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi_hi = _GEN_410;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi_hi = _GEN_410;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi_hi = _GEN_410;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi = {loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo = {loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_411 = {v0_825, v0_824};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo_lo = _GEN_411;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo_lo = _GEN_411;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo_lo = _GEN_411;
  wire [63:0]         _GEN_412 = {v0_827, v0_826};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo_hi = _GEN_412;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo_hi = _GEN_412;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo_hi = _GEN_412;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo = {loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_413 = {v0_829, v0_828};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi_lo = _GEN_413;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi_lo = _GEN_413;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi_lo = _GEN_413;
  wire [63:0]         _GEN_414 = {v0_831, v0_830};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi_hi = _GEN_414;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi_hi = _GEN_414;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi_hi = _GEN_414;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi = {loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi = {loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi = {loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_hi_hi_lo_lo_hi = {loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo};
  wire [2047:0]       loadUnit_maskInput_lo_hi_hi_lo_lo = {loadUnit_maskInput_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_415 = {v0_833, v0_832};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo_lo = _GEN_415;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo_lo = _GEN_415;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo_lo = _GEN_415;
  wire [63:0]         _GEN_416 = {v0_835, v0_834};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo_hi = _GEN_416;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo_hi = _GEN_416;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo_hi = _GEN_416;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo = {loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_417 = {v0_837, v0_836};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi_lo = _GEN_417;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi_lo = _GEN_417;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi_lo = _GEN_417;
  wire [63:0]         _GEN_418 = {v0_839, v0_838};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi_hi = _GEN_418;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi_hi = _GEN_418;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi_hi = _GEN_418;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi = {loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo = {loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_419 = {v0_841, v0_840};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo_lo = _GEN_419;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo_lo = _GEN_419;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo_lo = _GEN_419;
  wire [63:0]         _GEN_420 = {v0_843, v0_842};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo_hi = _GEN_420;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo_hi = _GEN_420;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo_hi = _GEN_420;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo = {loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_421 = {v0_845, v0_844};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi_lo = _GEN_421;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi_lo = _GEN_421;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi_lo = _GEN_421;
  wire [63:0]         _GEN_422 = {v0_847, v0_846};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi_hi = _GEN_422;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi_hi = _GEN_422;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi_hi = _GEN_422;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi = {loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi = {loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo = {loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_423 = {v0_849, v0_848};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo_lo = _GEN_423;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo_lo = _GEN_423;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo_lo = _GEN_423;
  wire [63:0]         _GEN_424 = {v0_851, v0_850};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo_hi = _GEN_424;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo_hi = _GEN_424;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo_hi = _GEN_424;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo = {loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_425 = {v0_853, v0_852};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi_lo = _GEN_425;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi_lo = _GEN_425;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi_lo = _GEN_425;
  wire [63:0]         _GEN_426 = {v0_855, v0_854};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi_hi = _GEN_426;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi_hi = _GEN_426;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi_hi = _GEN_426;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi = {loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo = {loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_427 = {v0_857, v0_856};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo_lo = _GEN_427;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo_lo = _GEN_427;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo_lo = _GEN_427;
  wire [63:0]         _GEN_428 = {v0_859, v0_858};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo_hi = _GEN_428;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo_hi = _GEN_428;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo_hi = _GEN_428;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo = {loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_429 = {v0_861, v0_860};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi_lo = _GEN_429;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi_lo = _GEN_429;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi_lo = _GEN_429;
  wire [63:0]         _GEN_430 = {v0_863, v0_862};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi_hi = _GEN_430;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi_hi = _GEN_430;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi_hi = _GEN_430;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi = {loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi = {loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi = {loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_hi_hi_lo_hi_lo = {loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_431 = {v0_865, v0_864};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo_lo = _GEN_431;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo_lo = _GEN_431;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo_lo = _GEN_431;
  wire [63:0]         _GEN_432 = {v0_867, v0_866};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo_hi = _GEN_432;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo_hi = _GEN_432;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo_hi = _GEN_432;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo = {loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_433 = {v0_869, v0_868};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi_lo = _GEN_433;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi_lo = _GEN_433;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi_lo = _GEN_433;
  wire [63:0]         _GEN_434 = {v0_871, v0_870};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi_hi = _GEN_434;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi_hi = _GEN_434;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi_hi = _GEN_434;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi = {loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo = {loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_435 = {v0_873, v0_872};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo_lo = _GEN_435;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo_lo = _GEN_435;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo_lo = _GEN_435;
  wire [63:0]         _GEN_436 = {v0_875, v0_874};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo_hi = _GEN_436;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo_hi = _GEN_436;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo_hi = _GEN_436;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo = {loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_437 = {v0_877, v0_876};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi_lo = _GEN_437;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi_lo = _GEN_437;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi_lo = _GEN_437;
  wire [63:0]         _GEN_438 = {v0_879, v0_878};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi_hi = _GEN_438;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi_hi = _GEN_438;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi_hi = _GEN_438;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi = {loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi = {loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo = {loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_439 = {v0_881, v0_880};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo_lo = _GEN_439;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo_lo = _GEN_439;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo_lo = _GEN_439;
  wire [63:0]         _GEN_440 = {v0_883, v0_882};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo_hi = _GEN_440;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo_hi = _GEN_440;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo_hi = _GEN_440;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo = {loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_441 = {v0_885, v0_884};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi_lo = _GEN_441;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi_lo = _GEN_441;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi_lo = _GEN_441;
  wire [63:0]         _GEN_442 = {v0_887, v0_886};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi_hi = _GEN_442;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi_hi = _GEN_442;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi_hi = _GEN_442;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi = {loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo = {loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_443 = {v0_889, v0_888};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo_lo = _GEN_443;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo_lo = _GEN_443;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo_lo = _GEN_443;
  wire [63:0]         _GEN_444 = {v0_891, v0_890};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo_hi = _GEN_444;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo_hi = _GEN_444;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo_hi = _GEN_444;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo = {loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_445 = {v0_893, v0_892};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi_lo = _GEN_445;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi_lo = _GEN_445;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi_lo = _GEN_445;
  wire [63:0]         _GEN_446 = {v0_895, v0_894};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi_hi = _GEN_446;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi_hi = _GEN_446;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi_hi = _GEN_446;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi = {loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi = {loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi = {loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_hi_hi_lo_hi_hi = {loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo};
  wire [2047:0]       loadUnit_maskInput_lo_hi_hi_lo_hi = {loadUnit_maskInput_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_lo};
  wire [4095:0]       loadUnit_maskInput_lo_hi_hi_lo = {loadUnit_maskInput_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_447 = {v0_897, v0_896};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo_lo = _GEN_447;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo_lo = _GEN_447;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo_lo = _GEN_447;
  wire [63:0]         _GEN_448 = {v0_899, v0_898};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo_hi = _GEN_448;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo_hi = _GEN_448;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo_hi = _GEN_448;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo = {loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_449 = {v0_901, v0_900};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi_lo = _GEN_449;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi_lo = _GEN_449;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi_lo = _GEN_449;
  wire [63:0]         _GEN_450 = {v0_903, v0_902};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi_hi = _GEN_450;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi_hi = _GEN_450;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi_hi = _GEN_450;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi = {loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo = {loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_451 = {v0_905, v0_904};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo_lo = _GEN_451;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo_lo = _GEN_451;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo_lo = _GEN_451;
  wire [63:0]         _GEN_452 = {v0_907, v0_906};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo_hi = _GEN_452;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo_hi = _GEN_452;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo_hi = _GEN_452;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo = {loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_453 = {v0_909, v0_908};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi_lo = _GEN_453;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi_lo = _GEN_453;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi_lo = _GEN_453;
  wire [63:0]         _GEN_454 = {v0_911, v0_910};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi_hi = _GEN_454;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi_hi = _GEN_454;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi_hi = _GEN_454;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi = {loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo = {loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_455 = {v0_913, v0_912};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo_lo = _GEN_455;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo_lo = _GEN_455;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo_lo = _GEN_455;
  wire [63:0]         _GEN_456 = {v0_915, v0_914};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo_hi = _GEN_456;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo_hi = _GEN_456;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo_hi = _GEN_456;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo = {loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_457 = {v0_917, v0_916};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi_lo = _GEN_457;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi_lo = _GEN_457;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi_lo = _GEN_457;
  wire [63:0]         _GEN_458 = {v0_919, v0_918};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi_hi = _GEN_458;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi_hi = _GEN_458;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi_hi = _GEN_458;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi = {loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo = {loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_459 = {v0_921, v0_920};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo_lo = _GEN_459;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo_lo = _GEN_459;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo_lo = _GEN_459;
  wire [63:0]         _GEN_460 = {v0_923, v0_922};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo_hi = _GEN_460;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo_hi = _GEN_460;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo_hi = _GEN_460;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo = {loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_461 = {v0_925, v0_924};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi_lo = _GEN_461;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi_lo = _GEN_461;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi_lo = _GEN_461;
  wire [63:0]         _GEN_462 = {v0_927, v0_926};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi_hi = _GEN_462;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi_hi = _GEN_462;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi_hi = _GEN_462;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi = {loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_hi_hi_hi_lo_lo = {loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_463 = {v0_929, v0_928};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo_lo = _GEN_463;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo_lo = _GEN_463;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo_lo = _GEN_463;
  wire [63:0]         _GEN_464 = {v0_931, v0_930};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo_hi = _GEN_464;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo_hi = _GEN_464;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo_hi = _GEN_464;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo = {loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_465 = {v0_933, v0_932};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi_lo = _GEN_465;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi_lo = _GEN_465;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi_lo = _GEN_465;
  wire [63:0]         _GEN_466 = {v0_935, v0_934};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi_hi = _GEN_466;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi_hi = _GEN_466;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi_hi = _GEN_466;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi = {loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo = {loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_467 = {v0_937, v0_936};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo_lo = _GEN_467;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo_lo = _GEN_467;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo_lo = _GEN_467;
  wire [63:0]         _GEN_468 = {v0_939, v0_938};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo_hi = _GEN_468;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo_hi = _GEN_468;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo_hi = _GEN_468;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo = {loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_469 = {v0_941, v0_940};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi_lo = _GEN_469;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi_lo = _GEN_469;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi_lo = _GEN_469;
  wire [63:0]         _GEN_470 = {v0_943, v0_942};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi_hi = _GEN_470;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi_hi = _GEN_470;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi_hi = _GEN_470;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi = {loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo = {loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_471 = {v0_945, v0_944};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo_lo = _GEN_471;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo_lo = _GEN_471;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo_lo = _GEN_471;
  wire [63:0]         _GEN_472 = {v0_947, v0_946};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo_hi = _GEN_472;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo_hi = _GEN_472;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo_hi = _GEN_472;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo = {loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_473 = {v0_949, v0_948};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi_lo = _GEN_473;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi_lo = _GEN_473;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi_lo = _GEN_473;
  wire [63:0]         _GEN_474 = {v0_951, v0_950};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi_hi = _GEN_474;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi_hi = _GEN_474;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi_hi = _GEN_474;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi = {loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo = {loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_475 = {v0_953, v0_952};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo_lo = _GEN_475;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo_lo = _GEN_475;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo_lo = _GEN_475;
  wire [63:0]         _GEN_476 = {v0_955, v0_954};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo_hi = _GEN_476;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo_hi = _GEN_476;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo_hi = _GEN_476;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo = {loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_477 = {v0_957, v0_956};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi_lo = _GEN_477;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi_lo = _GEN_477;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi_lo = _GEN_477;
  wire [63:0]         _GEN_478 = {v0_959, v0_958};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi_hi = _GEN_478;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi_hi = _GEN_478;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi_hi = _GEN_478;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_hi_hi_hi_lo_hi = {loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo};
  wire [2047:0]       loadUnit_maskInput_lo_hi_hi_hi_lo = {loadUnit_maskInput_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_479 = {v0_961, v0_960};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo_lo = _GEN_479;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo_lo = _GEN_479;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo_lo = _GEN_479;
  wire [63:0]         _GEN_480 = {v0_963, v0_962};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo_hi = _GEN_480;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo_hi = _GEN_480;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo_hi = _GEN_480;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo = {loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_481 = {v0_965, v0_964};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi_lo = _GEN_481;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi_lo = _GEN_481;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi_lo = _GEN_481;
  wire [63:0]         _GEN_482 = {v0_967, v0_966};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi_hi = _GEN_482;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi_hi = _GEN_482;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi_hi = _GEN_482;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi = {loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo = {loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_483 = {v0_969, v0_968};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo_lo = _GEN_483;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo_lo = _GEN_483;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo_lo = _GEN_483;
  wire [63:0]         _GEN_484 = {v0_971, v0_970};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo_hi = _GEN_484;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo_hi = _GEN_484;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo_hi = _GEN_484;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo = {loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_485 = {v0_973, v0_972};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi_lo = _GEN_485;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi_lo = _GEN_485;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi_lo = _GEN_485;
  wire [63:0]         _GEN_486 = {v0_975, v0_974};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi_hi = _GEN_486;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi_hi = _GEN_486;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi_hi = _GEN_486;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi = {loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo = {loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_487 = {v0_977, v0_976};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo_lo = _GEN_487;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo_lo = _GEN_487;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo_lo = _GEN_487;
  wire [63:0]         _GEN_488 = {v0_979, v0_978};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo_hi = _GEN_488;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo_hi = _GEN_488;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo_hi = _GEN_488;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo = {loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_489 = {v0_981, v0_980};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi_lo = _GEN_489;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi_lo = _GEN_489;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi_lo = _GEN_489;
  wire [63:0]         _GEN_490 = {v0_983, v0_982};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi_hi = _GEN_490;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi_hi = _GEN_490;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi_hi = _GEN_490;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi = {loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo = {loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_491 = {v0_985, v0_984};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo_lo = _GEN_491;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo_lo = _GEN_491;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo_lo = _GEN_491;
  wire [63:0]         _GEN_492 = {v0_987, v0_986};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo_hi = _GEN_492;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo_hi = _GEN_492;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo_hi = _GEN_492;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo = {loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_493 = {v0_989, v0_988};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi_lo = _GEN_493;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi_lo = _GEN_493;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi_lo = _GEN_493;
  wire [63:0]         _GEN_494 = {v0_991, v0_990};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi_hi = _GEN_494;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi_hi = _GEN_494;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi_hi = _GEN_494;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi = {loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_hi_hi_hi_hi_lo = {loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_495 = {v0_993, v0_992};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo_lo = _GEN_495;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo_lo = _GEN_495;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo_lo = _GEN_495;
  wire [63:0]         _GEN_496 = {v0_995, v0_994};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo_hi = _GEN_496;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo_hi = _GEN_496;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo_hi = _GEN_496;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo = {loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_497 = {v0_997, v0_996};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi_lo = _GEN_497;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi_lo = _GEN_497;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi_lo = _GEN_497;
  wire [63:0]         _GEN_498 = {v0_999, v0_998};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi_hi = _GEN_498;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi_hi = _GEN_498;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi_hi = _GEN_498;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi = {loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo = {loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_499 = {v0_1001, v0_1000};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo_lo = _GEN_499;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo_lo = _GEN_499;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo_lo = _GEN_499;
  wire [63:0]         _GEN_500 = {v0_1003, v0_1002};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo_hi = _GEN_500;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo_hi = _GEN_500;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo_hi = _GEN_500;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo = {loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_501 = {v0_1005, v0_1004};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi_lo = _GEN_501;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi_lo = _GEN_501;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi_lo = _GEN_501;
  wire [63:0]         _GEN_502 = {v0_1007, v0_1006};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi_hi = _GEN_502;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi_hi = _GEN_502;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi_hi = _GEN_502;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi = {loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo = {loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_503 = {v0_1009, v0_1008};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo_lo = _GEN_503;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo_lo = _GEN_503;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo_lo = _GEN_503;
  wire [63:0]         _GEN_504 = {v0_1011, v0_1010};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo_hi = _GEN_504;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo_hi = _GEN_504;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo_hi = _GEN_504;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo = {loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_505 = {v0_1013, v0_1012};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi_lo = _GEN_505;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi_lo = _GEN_505;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi_lo = _GEN_505;
  wire [63:0]         _GEN_506 = {v0_1015, v0_1014};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi_hi = _GEN_506;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi_hi = _GEN_506;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi_hi = _GEN_506;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi = {loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo = {loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_507 = {v0_1017, v0_1016};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo_lo = _GEN_507;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo_lo = _GEN_507;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo_lo = _GEN_507;
  wire [63:0]         _GEN_508 = {v0_1019, v0_1018};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo_hi = _GEN_508;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo_hi = _GEN_508;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo_hi = _GEN_508;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo = {loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_509 = {v0_1021, v0_1020};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi_lo = _GEN_509;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi_lo = _GEN_509;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi_lo = _GEN_509;
  wire [63:0]         _GEN_510 = {v0_1023, v0_1022};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi_hi = _GEN_510;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi_hi = _GEN_510;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi_hi = _GEN_510;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_hi_hi_hi_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo};
  wire [2047:0]       loadUnit_maskInput_lo_hi_hi_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_lo};
  wire [4095:0]       loadUnit_maskInput_lo_hi_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_lo};
  wire [8191:0]       loadUnit_maskInput_lo_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_lo};
  wire [16383:0]      loadUnit_maskInput_lo_hi = {loadUnit_maskInput_lo_hi_hi, loadUnit_maskInput_lo_hi_lo};
  wire [32767:0]      loadUnit_maskInput_lo = {loadUnit_maskInput_lo_hi, loadUnit_maskInput_lo_lo};
  wire [63:0]         _GEN_511 = {v0_1025, v0_1024};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo_lo = _GEN_511;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo_lo = _GEN_511;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo_lo = _GEN_511;
  wire [63:0]         _GEN_512 = {v0_1027, v0_1026};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo_hi = _GEN_512;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo_hi = _GEN_512;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo_hi = _GEN_512;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo = {loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_513 = {v0_1029, v0_1028};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi_lo = _GEN_513;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi_lo = _GEN_513;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi_lo = _GEN_513;
  wire [63:0]         _GEN_514 = {v0_1031, v0_1030};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi_hi = _GEN_514;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi_hi = _GEN_514;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi_hi = _GEN_514;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi = {loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo = {loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_515 = {v0_1033, v0_1032};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo_lo = _GEN_515;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo_lo = _GEN_515;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo_lo = _GEN_515;
  wire [63:0]         _GEN_516 = {v0_1035, v0_1034};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo_hi = _GEN_516;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo_hi = _GEN_516;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo_hi = _GEN_516;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo = {loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_517 = {v0_1037, v0_1036};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi_lo = _GEN_517;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi_lo = _GEN_517;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi_lo = _GEN_517;
  wire [63:0]         _GEN_518 = {v0_1039, v0_1038};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi_hi = _GEN_518;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi_hi = _GEN_518;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi_hi = _GEN_518;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi = {loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi = {loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo = {loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_519 = {v0_1041, v0_1040};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo_lo = _GEN_519;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo_lo = _GEN_519;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo_lo = _GEN_519;
  wire [63:0]         _GEN_520 = {v0_1043, v0_1042};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo_hi = _GEN_520;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo_hi = _GEN_520;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo_hi = _GEN_520;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo = {loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_521 = {v0_1045, v0_1044};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi_lo = _GEN_521;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi_lo = _GEN_521;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi_lo = _GEN_521;
  wire [63:0]         _GEN_522 = {v0_1047, v0_1046};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi_hi = _GEN_522;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi_hi = _GEN_522;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi_hi = _GEN_522;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi = {loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo = {loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_523 = {v0_1049, v0_1048};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo_lo = _GEN_523;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo_lo = _GEN_523;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo_lo = _GEN_523;
  wire [63:0]         _GEN_524 = {v0_1051, v0_1050};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo_hi = _GEN_524;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo_hi = _GEN_524;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo_hi = _GEN_524;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo = {loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_525 = {v0_1053, v0_1052};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi_lo = _GEN_525;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi_lo = _GEN_525;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi_lo = _GEN_525;
  wire [63:0]         _GEN_526 = {v0_1055, v0_1054};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi_hi = _GEN_526;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi_hi = _GEN_526;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi_hi = _GEN_526;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi = {loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi = {loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi = {loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_lo_lo_lo_lo_lo = {loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_527 = {v0_1057, v0_1056};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo_lo = _GEN_527;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo_lo = _GEN_527;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo_lo = _GEN_527;
  wire [63:0]         _GEN_528 = {v0_1059, v0_1058};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo_hi = _GEN_528;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo_hi = _GEN_528;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo_hi = _GEN_528;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo = {loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_529 = {v0_1061, v0_1060};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi_lo = _GEN_529;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi_lo = _GEN_529;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi_lo = _GEN_529;
  wire [63:0]         _GEN_530 = {v0_1063, v0_1062};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi_hi = _GEN_530;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi_hi = _GEN_530;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi_hi = _GEN_530;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi = {loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo = {loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_531 = {v0_1065, v0_1064};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo_lo = _GEN_531;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo_lo = _GEN_531;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo_lo = _GEN_531;
  wire [63:0]         _GEN_532 = {v0_1067, v0_1066};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo_hi = _GEN_532;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo_hi = _GEN_532;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo_hi = _GEN_532;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo = {loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_533 = {v0_1069, v0_1068};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi_lo = _GEN_533;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi_lo = _GEN_533;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi_lo = _GEN_533;
  wire [63:0]         _GEN_534 = {v0_1071, v0_1070};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi_hi = _GEN_534;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi_hi = _GEN_534;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi_hi = _GEN_534;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi = {loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi = {loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo = {loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_535 = {v0_1073, v0_1072};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo_lo = _GEN_535;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo_lo = _GEN_535;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo_lo = _GEN_535;
  wire [63:0]         _GEN_536 = {v0_1075, v0_1074};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo_hi = _GEN_536;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo_hi = _GEN_536;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo_hi = _GEN_536;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo = {loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_537 = {v0_1077, v0_1076};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi_lo = _GEN_537;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi_lo = _GEN_537;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi_lo = _GEN_537;
  wire [63:0]         _GEN_538 = {v0_1079, v0_1078};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi_hi = _GEN_538;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi_hi = _GEN_538;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi_hi = _GEN_538;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi = {loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo = {loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_539 = {v0_1081, v0_1080};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo_lo = _GEN_539;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo_lo = _GEN_539;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo_lo = _GEN_539;
  wire [63:0]         _GEN_540 = {v0_1083, v0_1082};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo_hi = _GEN_540;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo_hi = _GEN_540;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo_hi = _GEN_540;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo = {loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_541 = {v0_1085, v0_1084};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi_lo = _GEN_541;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi_lo = _GEN_541;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi_lo = _GEN_541;
  wire [63:0]         _GEN_542 = {v0_1087, v0_1086};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi_hi = _GEN_542;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi_hi = _GEN_542;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi_hi = _GEN_542;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi = {loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi = {loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi = {loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_lo_lo_lo_lo_hi = {loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo};
  wire [2047:0]       loadUnit_maskInput_hi_lo_lo_lo_lo = {loadUnit_maskInput_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_543 = {v0_1089, v0_1088};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo_lo = _GEN_543;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo_lo = _GEN_543;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo_lo = _GEN_543;
  wire [63:0]         _GEN_544 = {v0_1091, v0_1090};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo_hi = _GEN_544;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo_hi = _GEN_544;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo_hi = _GEN_544;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo = {loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_545 = {v0_1093, v0_1092};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi_lo = _GEN_545;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi_lo = _GEN_545;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi_lo = _GEN_545;
  wire [63:0]         _GEN_546 = {v0_1095, v0_1094};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi_hi = _GEN_546;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi_hi = _GEN_546;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi_hi = _GEN_546;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi = {loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo = {loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_547 = {v0_1097, v0_1096};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo_lo = _GEN_547;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo_lo = _GEN_547;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo_lo = _GEN_547;
  wire [63:0]         _GEN_548 = {v0_1099, v0_1098};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo_hi = _GEN_548;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo_hi = _GEN_548;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo_hi = _GEN_548;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo = {loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_549 = {v0_1101, v0_1100};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi_lo = _GEN_549;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi_lo = _GEN_549;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi_lo = _GEN_549;
  wire [63:0]         _GEN_550 = {v0_1103, v0_1102};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi_hi = _GEN_550;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi_hi = _GEN_550;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi_hi = _GEN_550;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi = {loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi = {loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo = {loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_551 = {v0_1105, v0_1104};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo_lo = _GEN_551;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo_lo = _GEN_551;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo_lo = _GEN_551;
  wire [63:0]         _GEN_552 = {v0_1107, v0_1106};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo_hi = _GEN_552;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo_hi = _GEN_552;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo_hi = _GEN_552;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo = {loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_553 = {v0_1109, v0_1108};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi_lo = _GEN_553;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi_lo = _GEN_553;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi_lo = _GEN_553;
  wire [63:0]         _GEN_554 = {v0_1111, v0_1110};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi_hi = _GEN_554;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi_hi = _GEN_554;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi_hi = _GEN_554;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi = {loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo = {loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_555 = {v0_1113, v0_1112};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo_lo = _GEN_555;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo_lo = _GEN_555;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo_lo = _GEN_555;
  wire [63:0]         _GEN_556 = {v0_1115, v0_1114};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo_hi = _GEN_556;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo_hi = _GEN_556;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo_hi = _GEN_556;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo = {loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_557 = {v0_1117, v0_1116};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi_lo = _GEN_557;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi_lo = _GEN_557;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi_lo = _GEN_557;
  wire [63:0]         _GEN_558 = {v0_1119, v0_1118};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi_hi = _GEN_558;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi_hi = _GEN_558;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi_hi = _GEN_558;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi = {loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi = {loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi = {loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_lo_lo_lo_hi_lo = {loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_559 = {v0_1121, v0_1120};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo_lo = _GEN_559;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo_lo = _GEN_559;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo_lo = _GEN_559;
  wire [63:0]         _GEN_560 = {v0_1123, v0_1122};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo_hi = _GEN_560;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo_hi = _GEN_560;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo_hi = _GEN_560;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo = {loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_561 = {v0_1125, v0_1124};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi_lo = _GEN_561;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi_lo = _GEN_561;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi_lo = _GEN_561;
  wire [63:0]         _GEN_562 = {v0_1127, v0_1126};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi_hi = _GEN_562;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi_hi = _GEN_562;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi_hi = _GEN_562;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi = {loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo = {loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_563 = {v0_1129, v0_1128};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo_lo = _GEN_563;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo_lo = _GEN_563;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo_lo = _GEN_563;
  wire [63:0]         _GEN_564 = {v0_1131, v0_1130};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo_hi = _GEN_564;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo_hi = _GEN_564;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo_hi = _GEN_564;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo = {loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_565 = {v0_1133, v0_1132};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi_lo = _GEN_565;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi_lo = _GEN_565;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi_lo = _GEN_565;
  wire [63:0]         _GEN_566 = {v0_1135, v0_1134};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi_hi = _GEN_566;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi_hi = _GEN_566;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi_hi = _GEN_566;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi = {loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi = {loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo = {loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_567 = {v0_1137, v0_1136};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo_lo = _GEN_567;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo_lo = _GEN_567;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo_lo = _GEN_567;
  wire [63:0]         _GEN_568 = {v0_1139, v0_1138};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo_hi = _GEN_568;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo_hi = _GEN_568;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo_hi = _GEN_568;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo = {loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_569 = {v0_1141, v0_1140};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi_lo = _GEN_569;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi_lo = _GEN_569;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi_lo = _GEN_569;
  wire [63:0]         _GEN_570 = {v0_1143, v0_1142};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi_hi = _GEN_570;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi_hi = _GEN_570;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi_hi = _GEN_570;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi = {loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo = {loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_571 = {v0_1145, v0_1144};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo_lo = _GEN_571;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo_lo = _GEN_571;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo_lo = _GEN_571;
  wire [63:0]         _GEN_572 = {v0_1147, v0_1146};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo_hi = _GEN_572;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo_hi = _GEN_572;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo_hi = _GEN_572;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo = {loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_573 = {v0_1149, v0_1148};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi_lo = _GEN_573;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi_lo = _GEN_573;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi_lo = _GEN_573;
  wire [63:0]         _GEN_574 = {v0_1151, v0_1150};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi_hi = _GEN_574;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi_hi = _GEN_574;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi_hi = _GEN_574;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi = {loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi = {loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi = {loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_lo_lo_lo_hi_hi = {loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo};
  wire [2047:0]       loadUnit_maskInput_hi_lo_lo_lo_hi = {loadUnit_maskInput_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_lo};
  wire [4095:0]       loadUnit_maskInput_hi_lo_lo_lo = {loadUnit_maskInput_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_575 = {v0_1153, v0_1152};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo_lo = _GEN_575;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo_lo = _GEN_575;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo_lo = _GEN_575;
  wire [63:0]         _GEN_576 = {v0_1155, v0_1154};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo_hi = _GEN_576;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo_hi = _GEN_576;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo_hi = _GEN_576;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo = {loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_577 = {v0_1157, v0_1156};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi_lo = _GEN_577;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi_lo = _GEN_577;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi_lo = _GEN_577;
  wire [63:0]         _GEN_578 = {v0_1159, v0_1158};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi_hi = _GEN_578;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi_hi = _GEN_578;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi_hi = _GEN_578;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi = {loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo = {loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_579 = {v0_1161, v0_1160};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo_lo = _GEN_579;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo_lo = _GEN_579;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo_lo = _GEN_579;
  wire [63:0]         _GEN_580 = {v0_1163, v0_1162};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo_hi = _GEN_580;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo_hi = _GEN_580;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo_hi = _GEN_580;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo = {loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_581 = {v0_1165, v0_1164};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi_lo = _GEN_581;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi_lo = _GEN_581;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi_lo = _GEN_581;
  wire [63:0]         _GEN_582 = {v0_1167, v0_1166};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi_hi = _GEN_582;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi_hi = _GEN_582;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi_hi = _GEN_582;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi = {loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi = {loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo = {loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_583 = {v0_1169, v0_1168};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo_lo = _GEN_583;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo_lo = _GEN_583;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo_lo = _GEN_583;
  wire [63:0]         _GEN_584 = {v0_1171, v0_1170};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo_hi = _GEN_584;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo_hi = _GEN_584;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo_hi = _GEN_584;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo = {loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_585 = {v0_1173, v0_1172};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi_lo = _GEN_585;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi_lo = _GEN_585;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi_lo = _GEN_585;
  wire [63:0]         _GEN_586 = {v0_1175, v0_1174};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi_hi = _GEN_586;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi_hi = _GEN_586;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi_hi = _GEN_586;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi = {loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo = {loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_587 = {v0_1177, v0_1176};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo_lo = _GEN_587;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo_lo = _GEN_587;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo_lo = _GEN_587;
  wire [63:0]         _GEN_588 = {v0_1179, v0_1178};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo_hi = _GEN_588;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo_hi = _GEN_588;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo_hi = _GEN_588;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo = {loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_589 = {v0_1181, v0_1180};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi_lo = _GEN_589;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi_lo = _GEN_589;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi_lo = _GEN_589;
  wire [63:0]         _GEN_590 = {v0_1183, v0_1182};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi_hi = _GEN_590;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi_hi = _GEN_590;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi_hi = _GEN_590;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi = {loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi = {loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi = {loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_lo_lo_hi_lo_lo = {loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_591 = {v0_1185, v0_1184};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo_lo = _GEN_591;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo_lo = _GEN_591;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo_lo = _GEN_591;
  wire [63:0]         _GEN_592 = {v0_1187, v0_1186};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo_hi = _GEN_592;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo_hi = _GEN_592;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo_hi = _GEN_592;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo = {loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_593 = {v0_1189, v0_1188};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi_lo = _GEN_593;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi_lo = _GEN_593;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi_lo = _GEN_593;
  wire [63:0]         _GEN_594 = {v0_1191, v0_1190};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi_hi = _GEN_594;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi_hi = _GEN_594;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi_hi = _GEN_594;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi = {loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo = {loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_595 = {v0_1193, v0_1192};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo_lo = _GEN_595;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo_lo = _GEN_595;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo_lo = _GEN_595;
  wire [63:0]         _GEN_596 = {v0_1195, v0_1194};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo_hi = _GEN_596;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo_hi = _GEN_596;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo_hi = _GEN_596;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo = {loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_597 = {v0_1197, v0_1196};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi_lo = _GEN_597;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi_lo = _GEN_597;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi_lo = _GEN_597;
  wire [63:0]         _GEN_598 = {v0_1199, v0_1198};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi_hi = _GEN_598;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi_hi = _GEN_598;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi_hi = _GEN_598;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi = {loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi = {loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo = {loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_599 = {v0_1201, v0_1200};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo_lo = _GEN_599;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo_lo = _GEN_599;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo_lo = _GEN_599;
  wire [63:0]         _GEN_600 = {v0_1203, v0_1202};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo_hi = _GEN_600;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo_hi = _GEN_600;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo_hi = _GEN_600;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo = {loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_601 = {v0_1205, v0_1204};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi_lo = _GEN_601;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi_lo = _GEN_601;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi_lo = _GEN_601;
  wire [63:0]         _GEN_602 = {v0_1207, v0_1206};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi_hi = _GEN_602;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi_hi = _GEN_602;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi_hi = _GEN_602;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi = {loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo = {loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_603 = {v0_1209, v0_1208};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo_lo = _GEN_603;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo_lo = _GEN_603;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo_lo = _GEN_603;
  wire [63:0]         _GEN_604 = {v0_1211, v0_1210};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo_hi = _GEN_604;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo_hi = _GEN_604;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo_hi = _GEN_604;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo = {loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_605 = {v0_1213, v0_1212};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi_lo = _GEN_605;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi_lo = _GEN_605;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi_lo = _GEN_605;
  wire [63:0]         _GEN_606 = {v0_1215, v0_1214};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi_hi = _GEN_606;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi_hi = _GEN_606;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi_hi = _GEN_606;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi = {loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi = {loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi = {loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_lo_lo_hi_lo_hi = {loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo};
  wire [2047:0]       loadUnit_maskInput_hi_lo_lo_hi_lo = {loadUnit_maskInput_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_607 = {v0_1217, v0_1216};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo_lo = _GEN_607;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo_lo = _GEN_607;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo_lo = _GEN_607;
  wire [63:0]         _GEN_608 = {v0_1219, v0_1218};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo_hi = _GEN_608;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo_hi = _GEN_608;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo_hi = _GEN_608;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo = {loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_609 = {v0_1221, v0_1220};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi_lo = _GEN_609;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi_lo = _GEN_609;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi_lo = _GEN_609;
  wire [63:0]         _GEN_610 = {v0_1223, v0_1222};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi_hi = _GEN_610;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi_hi = _GEN_610;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi_hi = _GEN_610;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi = {loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo = {loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_611 = {v0_1225, v0_1224};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo_lo = _GEN_611;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo_lo = _GEN_611;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo_lo = _GEN_611;
  wire [63:0]         _GEN_612 = {v0_1227, v0_1226};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo_hi = _GEN_612;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo_hi = _GEN_612;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo_hi = _GEN_612;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo = {loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_613 = {v0_1229, v0_1228};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi_lo = _GEN_613;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi_lo = _GEN_613;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi_lo = _GEN_613;
  wire [63:0]         _GEN_614 = {v0_1231, v0_1230};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi_hi = _GEN_614;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi_hi = _GEN_614;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi_hi = _GEN_614;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi = {loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi = {loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo = {loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_615 = {v0_1233, v0_1232};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo_lo = _GEN_615;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo_lo = _GEN_615;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo_lo = _GEN_615;
  wire [63:0]         _GEN_616 = {v0_1235, v0_1234};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo_hi = _GEN_616;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo_hi = _GEN_616;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo_hi = _GEN_616;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo = {loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_617 = {v0_1237, v0_1236};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi_lo = _GEN_617;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi_lo = _GEN_617;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi_lo = _GEN_617;
  wire [63:0]         _GEN_618 = {v0_1239, v0_1238};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi_hi = _GEN_618;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi_hi = _GEN_618;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi_hi = _GEN_618;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi = {loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo = {loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_619 = {v0_1241, v0_1240};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo_lo = _GEN_619;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo_lo = _GEN_619;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo_lo = _GEN_619;
  wire [63:0]         _GEN_620 = {v0_1243, v0_1242};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo_hi = _GEN_620;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo_hi = _GEN_620;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo_hi = _GEN_620;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo = {loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_621 = {v0_1245, v0_1244};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi_lo = _GEN_621;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi_lo = _GEN_621;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi_lo = _GEN_621;
  wire [63:0]         _GEN_622 = {v0_1247, v0_1246};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi_hi = _GEN_622;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi_hi = _GEN_622;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi_hi = _GEN_622;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi = {loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi = {loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi = {loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_lo_lo_hi_hi_lo = {loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_623 = {v0_1249, v0_1248};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo_lo = _GEN_623;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo_lo = _GEN_623;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo_lo = _GEN_623;
  wire [63:0]         _GEN_624 = {v0_1251, v0_1250};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo_hi = _GEN_624;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo_hi = _GEN_624;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo_hi = _GEN_624;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo = {loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_625 = {v0_1253, v0_1252};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi_lo = _GEN_625;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi_lo = _GEN_625;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi_lo = _GEN_625;
  wire [63:0]         _GEN_626 = {v0_1255, v0_1254};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi_hi = _GEN_626;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi_hi = _GEN_626;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi_hi = _GEN_626;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi = {loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo = {loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_627 = {v0_1257, v0_1256};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo_lo = _GEN_627;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo_lo = _GEN_627;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo_lo = _GEN_627;
  wire [63:0]         _GEN_628 = {v0_1259, v0_1258};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo_hi = _GEN_628;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo_hi = _GEN_628;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo_hi = _GEN_628;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo = {loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_629 = {v0_1261, v0_1260};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi_lo = _GEN_629;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi_lo = _GEN_629;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi_lo = _GEN_629;
  wire [63:0]         _GEN_630 = {v0_1263, v0_1262};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi_hi = _GEN_630;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi_hi = _GEN_630;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi_hi = _GEN_630;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi = {loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi = {loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo = {loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_631 = {v0_1265, v0_1264};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo_lo = _GEN_631;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo_lo = _GEN_631;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo_lo = _GEN_631;
  wire [63:0]         _GEN_632 = {v0_1267, v0_1266};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo_hi = _GEN_632;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo_hi = _GEN_632;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo_hi = _GEN_632;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo = {loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_633 = {v0_1269, v0_1268};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi_lo = _GEN_633;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi_lo = _GEN_633;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi_lo = _GEN_633;
  wire [63:0]         _GEN_634 = {v0_1271, v0_1270};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi_hi = _GEN_634;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi_hi = _GEN_634;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi_hi = _GEN_634;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi = {loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo = {loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_635 = {v0_1273, v0_1272};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo_lo = _GEN_635;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo_lo = _GEN_635;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo_lo = _GEN_635;
  wire [63:0]         _GEN_636 = {v0_1275, v0_1274};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo_hi = _GEN_636;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo_hi = _GEN_636;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo_hi = _GEN_636;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo = {loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_637 = {v0_1277, v0_1276};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi_lo = _GEN_637;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi_lo = _GEN_637;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi_lo = _GEN_637;
  wire [63:0]         _GEN_638 = {v0_1279, v0_1278};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi_hi = _GEN_638;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi_hi = _GEN_638;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi_hi = _GEN_638;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi = {loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi = {loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi = {loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_lo_lo_hi_hi_hi = {loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo};
  wire [2047:0]       loadUnit_maskInput_hi_lo_lo_hi_hi = {loadUnit_maskInput_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_lo};
  wire [4095:0]       loadUnit_maskInput_hi_lo_lo_hi = {loadUnit_maskInput_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_lo};
  wire [8191:0]       loadUnit_maskInput_hi_lo_lo = {loadUnit_maskInput_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo};
  wire [63:0]         _GEN_639 = {v0_1281, v0_1280};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo_lo = _GEN_639;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo_lo = _GEN_639;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo_lo = _GEN_639;
  wire [63:0]         _GEN_640 = {v0_1283, v0_1282};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo_hi = _GEN_640;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo_hi = _GEN_640;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo_hi = _GEN_640;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo = {loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_641 = {v0_1285, v0_1284};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi_lo = _GEN_641;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi_lo = _GEN_641;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi_lo = _GEN_641;
  wire [63:0]         _GEN_642 = {v0_1287, v0_1286};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi_hi = _GEN_642;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi_hi = _GEN_642;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi_hi = _GEN_642;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi = {loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo = {loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_643 = {v0_1289, v0_1288};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo_lo = _GEN_643;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo_lo = _GEN_643;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo_lo = _GEN_643;
  wire [63:0]         _GEN_644 = {v0_1291, v0_1290};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo_hi = _GEN_644;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo_hi = _GEN_644;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo_hi = _GEN_644;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo = {loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_645 = {v0_1293, v0_1292};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi_lo = _GEN_645;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi_lo = _GEN_645;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi_lo = _GEN_645;
  wire [63:0]         _GEN_646 = {v0_1295, v0_1294};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi_hi = _GEN_646;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi_hi = _GEN_646;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi_hi = _GEN_646;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi = {loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi = {loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo = {loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_647 = {v0_1297, v0_1296};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo_lo = _GEN_647;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo_lo = _GEN_647;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo_lo = _GEN_647;
  wire [63:0]         _GEN_648 = {v0_1299, v0_1298};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo_hi = _GEN_648;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo_hi = _GEN_648;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo_hi = _GEN_648;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo = {loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_649 = {v0_1301, v0_1300};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi_lo = _GEN_649;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi_lo = _GEN_649;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi_lo = _GEN_649;
  wire [63:0]         _GEN_650 = {v0_1303, v0_1302};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi_hi = _GEN_650;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi_hi = _GEN_650;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi_hi = _GEN_650;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo = {loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_651 = {v0_1305, v0_1304};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo_lo = _GEN_651;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo_lo = _GEN_651;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo_lo = _GEN_651;
  wire [63:0]         _GEN_652 = {v0_1307, v0_1306};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo_hi = _GEN_652;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo_hi = _GEN_652;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo_hi = _GEN_652;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo = {loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_653 = {v0_1309, v0_1308};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi_lo = _GEN_653;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi_lo = _GEN_653;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi_lo = _GEN_653;
  wire [63:0]         _GEN_654 = {v0_1311, v0_1310};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi_hi = _GEN_654;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi_hi = _GEN_654;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi_hi = _GEN_654;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi = {loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi = {loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi = {loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_lo_hi_lo_lo_lo = {loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_655 = {v0_1313, v0_1312};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo_lo = _GEN_655;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo_lo = _GEN_655;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo_lo = _GEN_655;
  wire [63:0]         _GEN_656 = {v0_1315, v0_1314};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo_hi = _GEN_656;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo_hi = _GEN_656;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo_hi = _GEN_656;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo = {loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_657 = {v0_1317, v0_1316};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi_lo = _GEN_657;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi_lo = _GEN_657;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi_lo = _GEN_657;
  wire [63:0]         _GEN_658 = {v0_1319, v0_1318};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi_hi = _GEN_658;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi_hi = _GEN_658;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi_hi = _GEN_658;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi = {loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo = {loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_659 = {v0_1321, v0_1320};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo_lo = _GEN_659;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo_lo = _GEN_659;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo_lo = _GEN_659;
  wire [63:0]         _GEN_660 = {v0_1323, v0_1322};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo_hi = _GEN_660;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo_hi = _GEN_660;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo_hi = _GEN_660;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo = {loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_661 = {v0_1325, v0_1324};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi_lo = _GEN_661;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi_lo = _GEN_661;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi_lo = _GEN_661;
  wire [63:0]         _GEN_662 = {v0_1327, v0_1326};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi_hi = _GEN_662;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi_hi = _GEN_662;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi_hi = _GEN_662;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi = {loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo = {loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_663 = {v0_1329, v0_1328};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo_lo = _GEN_663;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo_lo = _GEN_663;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo_lo = _GEN_663;
  wire [63:0]         _GEN_664 = {v0_1331, v0_1330};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo_hi = _GEN_664;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo_hi = _GEN_664;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo_hi = _GEN_664;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo = {loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_665 = {v0_1333, v0_1332};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi_lo = _GEN_665;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi_lo = _GEN_665;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi_lo = _GEN_665;
  wire [63:0]         _GEN_666 = {v0_1335, v0_1334};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi_hi = _GEN_666;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi_hi = _GEN_666;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi_hi = _GEN_666;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo = {loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_667 = {v0_1337, v0_1336};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo_lo = _GEN_667;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo_lo = _GEN_667;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo_lo = _GEN_667;
  wire [63:0]         _GEN_668 = {v0_1339, v0_1338};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo_hi = _GEN_668;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo_hi = _GEN_668;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo_hi = _GEN_668;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo = {loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_669 = {v0_1341, v0_1340};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi_lo = _GEN_669;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi_lo = _GEN_669;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi_lo = _GEN_669;
  wire [63:0]         _GEN_670 = {v0_1343, v0_1342};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi_hi = _GEN_670;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi_hi = _GEN_670;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi_hi = _GEN_670;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi = {loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi = {loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi = {loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_lo_hi_lo_lo_hi = {loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo};
  wire [2047:0]       loadUnit_maskInput_hi_lo_hi_lo_lo = {loadUnit_maskInput_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_671 = {v0_1345, v0_1344};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo_lo = _GEN_671;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo_lo = _GEN_671;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo_lo = _GEN_671;
  wire [63:0]         _GEN_672 = {v0_1347, v0_1346};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo_hi = _GEN_672;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo_hi = _GEN_672;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo_hi = _GEN_672;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo = {loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_673 = {v0_1349, v0_1348};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi_lo = _GEN_673;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi_lo = _GEN_673;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi_lo = _GEN_673;
  wire [63:0]         _GEN_674 = {v0_1351, v0_1350};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi_hi = _GEN_674;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi_hi = _GEN_674;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi_hi = _GEN_674;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi = {loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo = {loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_675 = {v0_1353, v0_1352};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo_lo = _GEN_675;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo_lo = _GEN_675;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo_lo = _GEN_675;
  wire [63:0]         _GEN_676 = {v0_1355, v0_1354};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo_hi = _GEN_676;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo_hi = _GEN_676;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo_hi = _GEN_676;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo = {loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_677 = {v0_1357, v0_1356};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi_lo = _GEN_677;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi_lo = _GEN_677;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi_lo = _GEN_677;
  wire [63:0]         _GEN_678 = {v0_1359, v0_1358};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi_hi = _GEN_678;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi_hi = _GEN_678;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi_hi = _GEN_678;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi = {loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi = {loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo = {loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_679 = {v0_1361, v0_1360};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo_lo = _GEN_679;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo_lo = _GEN_679;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo_lo = _GEN_679;
  wire [63:0]         _GEN_680 = {v0_1363, v0_1362};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo_hi = _GEN_680;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo_hi = _GEN_680;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo_hi = _GEN_680;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo = {loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_681 = {v0_1365, v0_1364};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi_lo = _GEN_681;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi_lo = _GEN_681;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi_lo = _GEN_681;
  wire [63:0]         _GEN_682 = {v0_1367, v0_1366};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi_hi = _GEN_682;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi_hi = _GEN_682;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi_hi = _GEN_682;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo = {loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_683 = {v0_1369, v0_1368};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo_lo = _GEN_683;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo_lo = _GEN_683;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo_lo = _GEN_683;
  wire [63:0]         _GEN_684 = {v0_1371, v0_1370};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo_hi = _GEN_684;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo_hi = _GEN_684;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo_hi = _GEN_684;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo = {loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_685 = {v0_1373, v0_1372};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi_lo = _GEN_685;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi_lo = _GEN_685;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi_lo = _GEN_685;
  wire [63:0]         _GEN_686 = {v0_1375, v0_1374};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi_hi = _GEN_686;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi_hi = _GEN_686;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi_hi = _GEN_686;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi = {loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi = {loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_lo_hi_lo_hi_lo = {loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_687 = {v0_1377, v0_1376};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo_lo = _GEN_687;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo_lo = _GEN_687;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo_lo = _GEN_687;
  wire [63:0]         _GEN_688 = {v0_1379, v0_1378};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo_hi = _GEN_688;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo_hi = _GEN_688;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo_hi = _GEN_688;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo = {loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_689 = {v0_1381, v0_1380};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi_lo = _GEN_689;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi_lo = _GEN_689;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi_lo = _GEN_689;
  wire [63:0]         _GEN_690 = {v0_1383, v0_1382};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi_hi = _GEN_690;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi_hi = _GEN_690;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi_hi = _GEN_690;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi = {loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo = {loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_691 = {v0_1385, v0_1384};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo_lo = _GEN_691;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo_lo = _GEN_691;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo_lo = _GEN_691;
  wire [63:0]         _GEN_692 = {v0_1387, v0_1386};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo_hi = _GEN_692;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo_hi = _GEN_692;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo_hi = _GEN_692;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo = {loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_693 = {v0_1389, v0_1388};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi_lo = _GEN_693;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi_lo = _GEN_693;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi_lo = _GEN_693;
  wire [63:0]         _GEN_694 = {v0_1391, v0_1390};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi_hi = _GEN_694;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi_hi = _GEN_694;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi_hi = _GEN_694;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi = {loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo = {loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_695 = {v0_1393, v0_1392};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo_lo = _GEN_695;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo_lo = _GEN_695;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo_lo = _GEN_695;
  wire [63:0]         _GEN_696 = {v0_1395, v0_1394};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo_hi = _GEN_696;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo_hi = _GEN_696;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo_hi = _GEN_696;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo = {loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_697 = {v0_1397, v0_1396};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi_lo = _GEN_697;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi_lo = _GEN_697;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi_lo = _GEN_697;
  wire [63:0]         _GEN_698 = {v0_1399, v0_1398};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi_hi = _GEN_698;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi_hi = _GEN_698;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi_hi = _GEN_698;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo = {loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_699 = {v0_1401, v0_1400};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo_lo = _GEN_699;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo_lo = _GEN_699;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo_lo = _GEN_699;
  wire [63:0]         _GEN_700 = {v0_1403, v0_1402};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo_hi = _GEN_700;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo_hi = _GEN_700;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo_hi = _GEN_700;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo = {loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_701 = {v0_1405, v0_1404};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi_lo = _GEN_701;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi_lo = _GEN_701;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi_lo = _GEN_701;
  wire [63:0]         _GEN_702 = {v0_1407, v0_1406};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi_hi = _GEN_702;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi_hi = _GEN_702;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi_hi = _GEN_702;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi = {loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi = {loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi = {loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_lo_hi_lo_hi_hi = {loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo};
  wire [2047:0]       loadUnit_maskInput_hi_lo_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_lo};
  wire [4095:0]       loadUnit_maskInput_hi_lo_hi_lo = {loadUnit_maskInput_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_703 = {v0_1409, v0_1408};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo_lo = _GEN_703;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo_lo = _GEN_703;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo_lo = _GEN_703;
  wire [63:0]         _GEN_704 = {v0_1411, v0_1410};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo_hi = _GEN_704;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo_hi = _GEN_704;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo_hi = _GEN_704;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo = {loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_705 = {v0_1413, v0_1412};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi_lo = _GEN_705;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi_lo = _GEN_705;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi_lo = _GEN_705;
  wire [63:0]         _GEN_706 = {v0_1415, v0_1414};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi_hi = _GEN_706;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi_hi = _GEN_706;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi_hi = _GEN_706;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi = {loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo = {loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_707 = {v0_1417, v0_1416};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo_lo = _GEN_707;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo_lo = _GEN_707;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo_lo = _GEN_707;
  wire [63:0]         _GEN_708 = {v0_1419, v0_1418};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo_hi = _GEN_708;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo_hi = _GEN_708;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo_hi = _GEN_708;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo = {loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_709 = {v0_1421, v0_1420};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi_lo = _GEN_709;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi_lo = _GEN_709;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi_lo = _GEN_709;
  wire [63:0]         _GEN_710 = {v0_1423, v0_1422};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi_hi = _GEN_710;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi_hi = _GEN_710;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi_hi = _GEN_710;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi = {loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi = {loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo = {loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_711 = {v0_1425, v0_1424};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo_lo = _GEN_711;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo_lo = _GEN_711;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo_lo = _GEN_711;
  wire [63:0]         _GEN_712 = {v0_1427, v0_1426};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo_hi = _GEN_712;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo_hi = _GEN_712;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo_hi = _GEN_712;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo = {loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_713 = {v0_1429, v0_1428};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi_lo = _GEN_713;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi_lo = _GEN_713;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi_lo = _GEN_713;
  wire [63:0]         _GEN_714 = {v0_1431, v0_1430};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi_hi = _GEN_714;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi_hi = _GEN_714;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi_hi = _GEN_714;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo = {loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_715 = {v0_1433, v0_1432};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo_lo = _GEN_715;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo_lo = _GEN_715;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo_lo = _GEN_715;
  wire [63:0]         _GEN_716 = {v0_1435, v0_1434};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo_hi = _GEN_716;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo_hi = _GEN_716;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo_hi = _GEN_716;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo = {loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_717 = {v0_1437, v0_1436};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi_lo = _GEN_717;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi_lo = _GEN_717;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi_lo = _GEN_717;
  wire [63:0]         _GEN_718 = {v0_1439, v0_1438};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi_hi = _GEN_718;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi_hi = _GEN_718;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi_hi = _GEN_718;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi = {loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi = {loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi = {loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_lo_hi_hi_lo_lo = {loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_719 = {v0_1441, v0_1440};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo_lo = _GEN_719;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo_lo = _GEN_719;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo_lo = _GEN_719;
  wire [63:0]         _GEN_720 = {v0_1443, v0_1442};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo_hi = _GEN_720;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo_hi = _GEN_720;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo_hi = _GEN_720;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo = {loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_721 = {v0_1445, v0_1444};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi_lo = _GEN_721;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi_lo = _GEN_721;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi_lo = _GEN_721;
  wire [63:0]         _GEN_722 = {v0_1447, v0_1446};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi_hi = _GEN_722;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi_hi = _GEN_722;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi_hi = _GEN_722;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi = {loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo = {loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_723 = {v0_1449, v0_1448};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo_lo = _GEN_723;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo_lo = _GEN_723;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo_lo = _GEN_723;
  wire [63:0]         _GEN_724 = {v0_1451, v0_1450};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo_hi = _GEN_724;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo_hi = _GEN_724;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo_hi = _GEN_724;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo = {loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_725 = {v0_1453, v0_1452};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi_lo = _GEN_725;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi_lo = _GEN_725;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi_lo = _GEN_725;
  wire [63:0]         _GEN_726 = {v0_1455, v0_1454};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi_hi = _GEN_726;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi_hi = _GEN_726;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi_hi = _GEN_726;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi = {loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo = {loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_727 = {v0_1457, v0_1456};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo_lo = _GEN_727;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo_lo = _GEN_727;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo_lo = _GEN_727;
  wire [63:0]         _GEN_728 = {v0_1459, v0_1458};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo_hi = _GEN_728;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo_hi = _GEN_728;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo_hi = _GEN_728;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo = {loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_729 = {v0_1461, v0_1460};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi_lo = _GEN_729;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi_lo = _GEN_729;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi_lo = _GEN_729;
  wire [63:0]         _GEN_730 = {v0_1463, v0_1462};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi_hi = _GEN_730;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi_hi = _GEN_730;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi_hi = _GEN_730;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo = {loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_731 = {v0_1465, v0_1464};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo_lo = _GEN_731;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo_lo = _GEN_731;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo_lo = _GEN_731;
  wire [63:0]         _GEN_732 = {v0_1467, v0_1466};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo_hi = _GEN_732;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo_hi = _GEN_732;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo_hi = _GEN_732;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo = {loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_733 = {v0_1469, v0_1468};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi_lo = _GEN_733;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi_lo = _GEN_733;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi_lo = _GEN_733;
  wire [63:0]         _GEN_734 = {v0_1471, v0_1470};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi_hi = _GEN_734;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi_hi = _GEN_734;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi_hi = _GEN_734;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi = {loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi = {loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi = {loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_lo_hi_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo};
  wire [2047:0]       loadUnit_maskInput_hi_lo_hi_hi_lo = {loadUnit_maskInput_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_735 = {v0_1473, v0_1472};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo_lo = _GEN_735;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo_lo = _GEN_735;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo_lo = _GEN_735;
  wire [63:0]         _GEN_736 = {v0_1475, v0_1474};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo_hi = _GEN_736;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo_hi = _GEN_736;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo_hi = _GEN_736;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo = {loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_737 = {v0_1477, v0_1476};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi_lo = _GEN_737;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi_lo = _GEN_737;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi_lo = _GEN_737;
  wire [63:0]         _GEN_738 = {v0_1479, v0_1478};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi_hi = _GEN_738;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi_hi = _GEN_738;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi_hi = _GEN_738;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi = {loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo = {loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_739 = {v0_1481, v0_1480};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo_lo = _GEN_739;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo_lo = _GEN_739;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo_lo = _GEN_739;
  wire [63:0]         _GEN_740 = {v0_1483, v0_1482};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo_hi = _GEN_740;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo_hi = _GEN_740;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo_hi = _GEN_740;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo = {loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_741 = {v0_1485, v0_1484};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi_lo = _GEN_741;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi_lo = _GEN_741;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi_lo = _GEN_741;
  wire [63:0]         _GEN_742 = {v0_1487, v0_1486};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi_hi = _GEN_742;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi_hi = _GEN_742;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi_hi = _GEN_742;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi = {loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi = {loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo = {loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_743 = {v0_1489, v0_1488};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo_lo = _GEN_743;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo_lo = _GEN_743;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo_lo = _GEN_743;
  wire [63:0]         _GEN_744 = {v0_1491, v0_1490};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo_hi = _GEN_744;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo_hi = _GEN_744;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo_hi = _GEN_744;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo = {loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_745 = {v0_1493, v0_1492};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi_lo = _GEN_745;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi_lo = _GEN_745;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi_lo = _GEN_745;
  wire [63:0]         _GEN_746 = {v0_1495, v0_1494};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi_hi = _GEN_746;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi_hi = _GEN_746;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi_hi = _GEN_746;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo = {loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_747 = {v0_1497, v0_1496};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo_lo = _GEN_747;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo_lo = _GEN_747;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo_lo = _GEN_747;
  wire [63:0]         _GEN_748 = {v0_1499, v0_1498};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo_hi = _GEN_748;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo_hi = _GEN_748;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo_hi = _GEN_748;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo = {loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_749 = {v0_1501, v0_1500};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi_lo = _GEN_749;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi_lo = _GEN_749;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi_lo = _GEN_749;
  wire [63:0]         _GEN_750 = {v0_1503, v0_1502};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi_hi = _GEN_750;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi_hi = _GEN_750;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi_hi = _GEN_750;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi = {loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi = {loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_lo_hi_hi_hi_lo = {loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_751 = {v0_1505, v0_1504};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo_lo = _GEN_751;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo_lo = _GEN_751;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo_lo = _GEN_751;
  wire [63:0]         _GEN_752 = {v0_1507, v0_1506};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo_hi = _GEN_752;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo_hi = _GEN_752;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo_hi = _GEN_752;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo = {loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_753 = {v0_1509, v0_1508};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi_lo = _GEN_753;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi_lo = _GEN_753;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi_lo = _GEN_753;
  wire [63:0]         _GEN_754 = {v0_1511, v0_1510};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi_hi = _GEN_754;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi_hi = _GEN_754;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi_hi = _GEN_754;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi = {loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo = {loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_755 = {v0_1513, v0_1512};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo_lo = _GEN_755;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo_lo = _GEN_755;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo_lo = _GEN_755;
  wire [63:0]         _GEN_756 = {v0_1515, v0_1514};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo_hi = _GEN_756;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo_hi = _GEN_756;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo_hi = _GEN_756;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo = {loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_757 = {v0_1517, v0_1516};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi_lo = _GEN_757;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi_lo = _GEN_757;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi_lo = _GEN_757;
  wire [63:0]         _GEN_758 = {v0_1519, v0_1518};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi_hi = _GEN_758;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi_hi = _GEN_758;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi_hi = _GEN_758;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi = {loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo = {loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_759 = {v0_1521, v0_1520};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo_lo = _GEN_759;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo_lo = _GEN_759;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo_lo = _GEN_759;
  wire [63:0]         _GEN_760 = {v0_1523, v0_1522};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo_hi = _GEN_760;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo_hi = _GEN_760;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo_hi = _GEN_760;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo = {loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_761 = {v0_1525, v0_1524};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi_lo = _GEN_761;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi_lo = _GEN_761;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi_lo = _GEN_761;
  wire [63:0]         _GEN_762 = {v0_1527, v0_1526};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi_hi = _GEN_762;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi_hi = _GEN_762;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi_hi = _GEN_762;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo = {loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_763 = {v0_1529, v0_1528};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo_lo = _GEN_763;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo_lo = _GEN_763;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo_lo = _GEN_763;
  wire [63:0]         _GEN_764 = {v0_1531, v0_1530};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo_hi = _GEN_764;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo_hi = _GEN_764;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo_hi = _GEN_764;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo = {loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_765 = {v0_1533, v0_1532};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi_lo = _GEN_765;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi_lo = _GEN_765;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi_lo = _GEN_765;
  wire [63:0]         _GEN_766 = {v0_1535, v0_1534};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi_hi = _GEN_766;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi_hi = _GEN_766;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi_hi = _GEN_766;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi = {loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi = {loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi = {loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_lo_hi_hi_hi_hi = {loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo};
  wire [2047:0]       loadUnit_maskInput_hi_lo_hi_hi_hi = {loadUnit_maskInput_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_lo};
  wire [4095:0]       loadUnit_maskInput_hi_lo_hi_hi = {loadUnit_maskInput_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_lo};
  wire [8191:0]       loadUnit_maskInput_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo};
  wire [16383:0]      loadUnit_maskInput_hi_lo = {loadUnit_maskInput_hi_lo_hi, loadUnit_maskInput_hi_lo_lo};
  wire [63:0]         _GEN_767 = {v0_1537, v0_1536};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo_lo = _GEN_767;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo_lo = _GEN_767;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo_lo = _GEN_767;
  wire [63:0]         _GEN_768 = {v0_1539, v0_1538};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo_hi = _GEN_768;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo_hi = _GEN_768;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo_hi = _GEN_768;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo = {loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_769 = {v0_1541, v0_1540};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi_lo = _GEN_769;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi_lo = _GEN_769;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi_lo = _GEN_769;
  wire [63:0]         _GEN_770 = {v0_1543, v0_1542};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi_hi = _GEN_770;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi_hi = _GEN_770;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi_hi = _GEN_770;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi = {loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo = {loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_771 = {v0_1545, v0_1544};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo_lo = _GEN_771;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo_lo = _GEN_771;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo_lo = _GEN_771;
  wire [63:0]         _GEN_772 = {v0_1547, v0_1546};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo_hi = _GEN_772;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo_hi = _GEN_772;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo_hi = _GEN_772;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo = {loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_773 = {v0_1549, v0_1548};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi_lo = _GEN_773;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi_lo = _GEN_773;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi_lo = _GEN_773;
  wire [63:0]         _GEN_774 = {v0_1551, v0_1550};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi_hi = _GEN_774;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi_hi = _GEN_774;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi_hi = _GEN_774;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi = {loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi = {loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo = {loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_775 = {v0_1553, v0_1552};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo_lo = _GEN_775;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo_lo = _GEN_775;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo_lo = _GEN_775;
  wire [63:0]         _GEN_776 = {v0_1555, v0_1554};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo_hi = _GEN_776;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo_hi = _GEN_776;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo_hi = _GEN_776;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo = {loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_777 = {v0_1557, v0_1556};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi_lo = _GEN_777;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi_lo = _GEN_777;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi_lo = _GEN_777;
  wire [63:0]         _GEN_778 = {v0_1559, v0_1558};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi_hi = _GEN_778;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi_hi = _GEN_778;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi_hi = _GEN_778;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi = {loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo = {loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_779 = {v0_1561, v0_1560};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo_lo = _GEN_779;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo_lo = _GEN_779;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo_lo = _GEN_779;
  wire [63:0]         _GEN_780 = {v0_1563, v0_1562};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo_hi = _GEN_780;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo_hi = _GEN_780;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo_hi = _GEN_780;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo = {loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_781 = {v0_1565, v0_1564};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi_lo = _GEN_781;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi_lo = _GEN_781;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi_lo = _GEN_781;
  wire [63:0]         _GEN_782 = {v0_1567, v0_1566};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi_hi = _GEN_782;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi_hi = _GEN_782;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi_hi = _GEN_782;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi = {loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi = {loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi = {loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_hi_lo_lo_lo_lo = {loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_783 = {v0_1569, v0_1568};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo_lo = _GEN_783;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo_lo = _GEN_783;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo_lo = _GEN_783;
  wire [63:0]         _GEN_784 = {v0_1571, v0_1570};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo_hi = _GEN_784;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo_hi = _GEN_784;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo_hi = _GEN_784;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo = {loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_785 = {v0_1573, v0_1572};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi_lo = _GEN_785;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi_lo = _GEN_785;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi_lo = _GEN_785;
  wire [63:0]         _GEN_786 = {v0_1575, v0_1574};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi_hi = _GEN_786;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi_hi = _GEN_786;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi_hi = _GEN_786;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi = {loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo = {loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_787 = {v0_1577, v0_1576};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo_lo = _GEN_787;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo_lo = _GEN_787;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo_lo = _GEN_787;
  wire [63:0]         _GEN_788 = {v0_1579, v0_1578};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo_hi = _GEN_788;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo_hi = _GEN_788;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo_hi = _GEN_788;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo = {loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_789 = {v0_1581, v0_1580};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi_lo = _GEN_789;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi_lo = _GEN_789;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi_lo = _GEN_789;
  wire [63:0]         _GEN_790 = {v0_1583, v0_1582};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi_hi = _GEN_790;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi_hi = _GEN_790;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi_hi = _GEN_790;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi = {loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi = {loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo = {loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_791 = {v0_1585, v0_1584};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo_lo = _GEN_791;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo_lo = _GEN_791;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo_lo = _GEN_791;
  wire [63:0]         _GEN_792 = {v0_1587, v0_1586};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo_hi = _GEN_792;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo_hi = _GEN_792;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo_hi = _GEN_792;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo = {loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_793 = {v0_1589, v0_1588};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi_lo = _GEN_793;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi_lo = _GEN_793;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi_lo = _GEN_793;
  wire [63:0]         _GEN_794 = {v0_1591, v0_1590};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi_hi = _GEN_794;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi_hi = _GEN_794;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi_hi = _GEN_794;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi = {loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo = {loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_795 = {v0_1593, v0_1592};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo_lo = _GEN_795;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo_lo = _GEN_795;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo_lo = _GEN_795;
  wire [63:0]         _GEN_796 = {v0_1595, v0_1594};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo_hi = _GEN_796;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo_hi = _GEN_796;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo_hi = _GEN_796;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo = {loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_797 = {v0_1597, v0_1596};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi_lo = _GEN_797;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi_lo = _GEN_797;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi_lo = _GEN_797;
  wire [63:0]         _GEN_798 = {v0_1599, v0_1598};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi_hi = _GEN_798;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi_hi = _GEN_798;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi_hi = _GEN_798;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi = {loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi = {loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi = {loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_hi_lo_lo_lo_hi = {loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo};
  wire [2047:0]       loadUnit_maskInput_hi_hi_lo_lo_lo = {loadUnit_maskInput_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_799 = {v0_1601, v0_1600};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo_lo = _GEN_799;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo_lo = _GEN_799;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo_lo = _GEN_799;
  wire [63:0]         _GEN_800 = {v0_1603, v0_1602};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo_hi = _GEN_800;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo_hi = _GEN_800;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo_hi = _GEN_800;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo = {loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_801 = {v0_1605, v0_1604};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi_lo = _GEN_801;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi_lo = _GEN_801;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi_lo = _GEN_801;
  wire [63:0]         _GEN_802 = {v0_1607, v0_1606};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi_hi = _GEN_802;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi_hi = _GEN_802;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi_hi = _GEN_802;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi = {loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo = {loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_803 = {v0_1609, v0_1608};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo_lo = _GEN_803;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo_lo = _GEN_803;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo_lo = _GEN_803;
  wire [63:0]         _GEN_804 = {v0_1611, v0_1610};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo_hi = _GEN_804;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo_hi = _GEN_804;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo_hi = _GEN_804;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo = {loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_805 = {v0_1613, v0_1612};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi_lo = _GEN_805;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi_lo = _GEN_805;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi_lo = _GEN_805;
  wire [63:0]         _GEN_806 = {v0_1615, v0_1614};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi_hi = _GEN_806;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi_hi = _GEN_806;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi_hi = _GEN_806;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi = {loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi = {loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo = {loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_807 = {v0_1617, v0_1616};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo_lo = _GEN_807;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo_lo = _GEN_807;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo_lo = _GEN_807;
  wire [63:0]         _GEN_808 = {v0_1619, v0_1618};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo_hi = _GEN_808;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo_hi = _GEN_808;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo_hi = _GEN_808;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo = {loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_809 = {v0_1621, v0_1620};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi_lo = _GEN_809;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi_lo = _GEN_809;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi_lo = _GEN_809;
  wire [63:0]         _GEN_810 = {v0_1623, v0_1622};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi_hi = _GEN_810;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi_hi = _GEN_810;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi_hi = _GEN_810;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi = {loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo = {loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_811 = {v0_1625, v0_1624};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo_lo = _GEN_811;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo_lo = _GEN_811;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo_lo = _GEN_811;
  wire [63:0]         _GEN_812 = {v0_1627, v0_1626};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo_hi = _GEN_812;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo_hi = _GEN_812;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo_hi = _GEN_812;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo = {loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_813 = {v0_1629, v0_1628};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi_lo = _GEN_813;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi_lo = _GEN_813;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi_lo = _GEN_813;
  wire [63:0]         _GEN_814 = {v0_1631, v0_1630};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi_hi = _GEN_814;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi_hi = _GEN_814;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi_hi = _GEN_814;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi = {loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi = {loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi = {loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_hi_lo_lo_hi_lo = {loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_815 = {v0_1633, v0_1632};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo_lo = _GEN_815;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo_lo = _GEN_815;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo_lo = _GEN_815;
  wire [63:0]         _GEN_816 = {v0_1635, v0_1634};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo_hi = _GEN_816;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo_hi = _GEN_816;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo_hi = _GEN_816;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo = {loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_817 = {v0_1637, v0_1636};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi_lo = _GEN_817;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi_lo = _GEN_817;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi_lo = _GEN_817;
  wire [63:0]         _GEN_818 = {v0_1639, v0_1638};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi_hi = _GEN_818;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi_hi = _GEN_818;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi_hi = _GEN_818;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi = {loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo = {loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_819 = {v0_1641, v0_1640};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo_lo = _GEN_819;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo_lo = _GEN_819;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo_lo = _GEN_819;
  wire [63:0]         _GEN_820 = {v0_1643, v0_1642};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo_hi = _GEN_820;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo_hi = _GEN_820;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo_hi = _GEN_820;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo = {loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_821 = {v0_1645, v0_1644};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi_lo = _GEN_821;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi_lo = _GEN_821;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi_lo = _GEN_821;
  wire [63:0]         _GEN_822 = {v0_1647, v0_1646};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi_hi = _GEN_822;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi_hi = _GEN_822;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi_hi = _GEN_822;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi = {loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi = {loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo = {loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_823 = {v0_1649, v0_1648};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo_lo = _GEN_823;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo_lo = _GEN_823;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo_lo = _GEN_823;
  wire [63:0]         _GEN_824 = {v0_1651, v0_1650};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo_hi = _GEN_824;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo_hi = _GEN_824;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo_hi = _GEN_824;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo = {loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_825 = {v0_1653, v0_1652};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi_lo = _GEN_825;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi_lo = _GEN_825;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi_lo = _GEN_825;
  wire [63:0]         _GEN_826 = {v0_1655, v0_1654};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi_hi = _GEN_826;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi_hi = _GEN_826;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi_hi = _GEN_826;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi = {loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo = {loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_827 = {v0_1657, v0_1656};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo_lo = _GEN_827;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo_lo = _GEN_827;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo_lo = _GEN_827;
  wire [63:0]         _GEN_828 = {v0_1659, v0_1658};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo_hi = _GEN_828;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo_hi = _GEN_828;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo_hi = _GEN_828;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo = {loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_829 = {v0_1661, v0_1660};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi_lo = _GEN_829;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi_lo = _GEN_829;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi_lo = _GEN_829;
  wire [63:0]         _GEN_830 = {v0_1663, v0_1662};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi_hi = _GEN_830;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi_hi = _GEN_830;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi_hi = _GEN_830;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi = {loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi = {loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi = {loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_hi_lo_lo_hi_hi = {loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo};
  wire [2047:0]       loadUnit_maskInput_hi_hi_lo_lo_hi = {loadUnit_maskInput_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_lo};
  wire [4095:0]       loadUnit_maskInput_hi_hi_lo_lo = {loadUnit_maskInput_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_831 = {v0_1665, v0_1664};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo_lo = _GEN_831;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo_lo = _GEN_831;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo_lo = _GEN_831;
  wire [63:0]         _GEN_832 = {v0_1667, v0_1666};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo_hi = _GEN_832;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo_hi = _GEN_832;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo_hi = _GEN_832;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo = {loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_833 = {v0_1669, v0_1668};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi_lo = _GEN_833;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi_lo = _GEN_833;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi_lo = _GEN_833;
  wire [63:0]         _GEN_834 = {v0_1671, v0_1670};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi_hi = _GEN_834;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi_hi = _GEN_834;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi_hi = _GEN_834;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi = {loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo = {loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_835 = {v0_1673, v0_1672};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo_lo = _GEN_835;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo_lo = _GEN_835;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo_lo = _GEN_835;
  wire [63:0]         _GEN_836 = {v0_1675, v0_1674};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo_hi = _GEN_836;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo_hi = _GEN_836;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo_hi = _GEN_836;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_837 = {v0_1677, v0_1676};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi_lo = _GEN_837;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi_lo = _GEN_837;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi_lo = _GEN_837;
  wire [63:0]         _GEN_838 = {v0_1679, v0_1678};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi_hi = _GEN_838;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi_hi = _GEN_838;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi_hi = _GEN_838;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi = {loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi = {loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo = {loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_839 = {v0_1681, v0_1680};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo_lo = _GEN_839;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo_lo = _GEN_839;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo_lo = _GEN_839;
  wire [63:0]         _GEN_840 = {v0_1683, v0_1682};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo_hi = _GEN_840;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo_hi = _GEN_840;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo_hi = _GEN_840;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo = {loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_841 = {v0_1685, v0_1684};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi_lo = _GEN_841;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi_lo = _GEN_841;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi_lo = _GEN_841;
  wire [63:0]         _GEN_842 = {v0_1687, v0_1686};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi_hi = _GEN_842;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi_hi = _GEN_842;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi_hi = _GEN_842;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi = {loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_843 = {v0_1689, v0_1688};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo_lo = _GEN_843;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo_lo = _GEN_843;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo_lo = _GEN_843;
  wire [63:0]         _GEN_844 = {v0_1691, v0_1690};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo_hi = _GEN_844;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo_hi = _GEN_844;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo_hi = _GEN_844;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_845 = {v0_1693, v0_1692};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi_lo = _GEN_845;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi_lo = _GEN_845;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi_lo = _GEN_845;
  wire [63:0]         _GEN_846 = {v0_1695, v0_1694};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi_hi = _GEN_846;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi_hi = _GEN_846;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi_hi = _GEN_846;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi = {loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi = {loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi = {loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_hi_lo_hi_lo_lo = {loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_847 = {v0_1697, v0_1696};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo_lo = _GEN_847;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo_lo = _GEN_847;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo_lo = _GEN_847;
  wire [63:0]         _GEN_848 = {v0_1699, v0_1698};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo_hi = _GEN_848;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo_hi = _GEN_848;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo_hi = _GEN_848;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo = {loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_849 = {v0_1701, v0_1700};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi_lo = _GEN_849;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi_lo = _GEN_849;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi_lo = _GEN_849;
  wire [63:0]         _GEN_850 = {v0_1703, v0_1702};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi_hi = _GEN_850;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi_hi = _GEN_850;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi_hi = _GEN_850;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi = {loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo = {loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_851 = {v0_1705, v0_1704};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo_lo = _GEN_851;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo_lo = _GEN_851;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo_lo = _GEN_851;
  wire [63:0]         _GEN_852 = {v0_1707, v0_1706};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo_hi = _GEN_852;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo_hi = _GEN_852;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo_hi = _GEN_852;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_853 = {v0_1709, v0_1708};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi_lo = _GEN_853;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi_lo = _GEN_853;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi_lo = _GEN_853;
  wire [63:0]         _GEN_854 = {v0_1711, v0_1710};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi_hi = _GEN_854;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi_hi = _GEN_854;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi_hi = _GEN_854;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi = {loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi = {loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_855 = {v0_1713, v0_1712};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo_lo = _GEN_855;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo_lo = _GEN_855;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo_lo = _GEN_855;
  wire [63:0]         _GEN_856 = {v0_1715, v0_1714};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo_hi = _GEN_856;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo_hi = _GEN_856;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo_hi = _GEN_856;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo = {loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_857 = {v0_1717, v0_1716};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi_lo = _GEN_857;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi_lo = _GEN_857;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi_lo = _GEN_857;
  wire [63:0]         _GEN_858 = {v0_1719, v0_1718};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi_hi = _GEN_858;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi_hi = _GEN_858;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi_hi = _GEN_858;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi = {loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_859 = {v0_1721, v0_1720};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo_lo = _GEN_859;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo_lo = _GEN_859;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo_lo = _GEN_859;
  wire [63:0]         _GEN_860 = {v0_1723, v0_1722};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo_hi = _GEN_860;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo_hi = _GEN_860;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo_hi = _GEN_860;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_861 = {v0_1725, v0_1724};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi_lo = _GEN_861;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi_lo = _GEN_861;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi_lo = _GEN_861;
  wire [63:0]         _GEN_862 = {v0_1727, v0_1726};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi_hi = _GEN_862;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi_hi = _GEN_862;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi_hi = _GEN_862;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi = {loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi = {loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi = {loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_hi_lo_hi_lo_hi = {loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo};
  wire [2047:0]       loadUnit_maskInput_hi_hi_lo_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_863 = {v0_1729, v0_1728};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo_lo = _GEN_863;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo_lo = _GEN_863;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo_lo = _GEN_863;
  wire [63:0]         _GEN_864 = {v0_1731, v0_1730};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo_hi = _GEN_864;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo_hi = _GEN_864;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo_hi = _GEN_864;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo = {loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_865 = {v0_1733, v0_1732};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi_lo = _GEN_865;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi_lo = _GEN_865;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi_lo = _GEN_865;
  wire [63:0]         _GEN_866 = {v0_1735, v0_1734};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi_hi = _GEN_866;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi_hi = _GEN_866;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi_hi = _GEN_866;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi = {loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo = {loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_867 = {v0_1737, v0_1736};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo_lo = _GEN_867;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo_lo = _GEN_867;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo_lo = _GEN_867;
  wire [63:0]         _GEN_868 = {v0_1739, v0_1738};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo_hi = _GEN_868;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo_hi = _GEN_868;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo_hi = _GEN_868;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_869 = {v0_1741, v0_1740};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi_lo = _GEN_869;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi_lo = _GEN_869;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi_lo = _GEN_869;
  wire [63:0]         _GEN_870 = {v0_1743, v0_1742};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi_hi = _GEN_870;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi_hi = _GEN_870;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi_hi = _GEN_870;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi = {loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi = {loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo = {loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_871 = {v0_1745, v0_1744};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo_lo = _GEN_871;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo_lo = _GEN_871;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo_lo = _GEN_871;
  wire [63:0]         _GEN_872 = {v0_1747, v0_1746};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo_hi = _GEN_872;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo_hi = _GEN_872;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo_hi = _GEN_872;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo = {loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_873 = {v0_1749, v0_1748};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi_lo = _GEN_873;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi_lo = _GEN_873;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi_lo = _GEN_873;
  wire [63:0]         _GEN_874 = {v0_1751, v0_1750};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi_hi = _GEN_874;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi_hi = _GEN_874;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi_hi = _GEN_874;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi = {loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_875 = {v0_1753, v0_1752};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo_lo = _GEN_875;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo_lo = _GEN_875;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo_lo = _GEN_875;
  wire [63:0]         _GEN_876 = {v0_1755, v0_1754};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo_hi = _GEN_876;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo_hi = _GEN_876;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo_hi = _GEN_876;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_877 = {v0_1757, v0_1756};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi_lo = _GEN_877;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi_lo = _GEN_877;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi_lo = _GEN_877;
  wire [63:0]         _GEN_878 = {v0_1759, v0_1758};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi_hi = _GEN_878;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi_hi = _GEN_878;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi_hi = _GEN_878;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi = {loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi = {loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi = {loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_hi_lo_hi_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_879 = {v0_1761, v0_1760};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo_lo = _GEN_879;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo_lo = _GEN_879;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo_lo = _GEN_879;
  wire [63:0]         _GEN_880 = {v0_1763, v0_1762};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo_hi = _GEN_880;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo_hi = _GEN_880;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo_hi = _GEN_880;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo = {loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_881 = {v0_1765, v0_1764};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi_lo = _GEN_881;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi_lo = _GEN_881;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi_lo = _GEN_881;
  wire [63:0]         _GEN_882 = {v0_1767, v0_1766};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi_hi = _GEN_882;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi_hi = _GEN_882;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi_hi = _GEN_882;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi = {loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo = {loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_883 = {v0_1769, v0_1768};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo_lo = _GEN_883;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo_lo = _GEN_883;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo_lo = _GEN_883;
  wire [63:0]         _GEN_884 = {v0_1771, v0_1770};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo_hi = _GEN_884;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo_hi = _GEN_884;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo_hi = _GEN_884;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_885 = {v0_1773, v0_1772};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi_lo = _GEN_885;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi_lo = _GEN_885;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi_lo = _GEN_885;
  wire [63:0]         _GEN_886 = {v0_1775, v0_1774};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi_hi = _GEN_886;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi_hi = _GEN_886;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi_hi = _GEN_886;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi = {loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi = {loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_887 = {v0_1777, v0_1776};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo_lo = _GEN_887;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo_lo = _GEN_887;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo_lo = _GEN_887;
  wire [63:0]         _GEN_888 = {v0_1779, v0_1778};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo_hi = _GEN_888;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo_hi = _GEN_888;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo_hi = _GEN_888;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo = {loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_889 = {v0_1781, v0_1780};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi_lo = _GEN_889;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi_lo = _GEN_889;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi_lo = _GEN_889;
  wire [63:0]         _GEN_890 = {v0_1783, v0_1782};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi_hi = _GEN_890;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi_hi = _GEN_890;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi_hi = _GEN_890;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi = {loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_891 = {v0_1785, v0_1784};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo_lo = _GEN_891;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo_lo = _GEN_891;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo_lo = _GEN_891;
  wire [63:0]         _GEN_892 = {v0_1787, v0_1786};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo_hi = _GEN_892;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo_hi = _GEN_892;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo_hi = _GEN_892;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_893 = {v0_1789, v0_1788};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi_lo = _GEN_893;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi_lo = _GEN_893;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi_lo = _GEN_893;
  wire [63:0]         _GEN_894 = {v0_1791, v0_1790};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi_hi = _GEN_894;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi_hi = _GEN_894;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi_hi = _GEN_894;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi = {loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi = {loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi = {loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_hi_lo_hi_hi_hi = {loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo};
  wire [2047:0]       loadUnit_maskInput_hi_hi_lo_hi_hi = {loadUnit_maskInput_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_lo};
  wire [4095:0]       loadUnit_maskInput_hi_hi_lo_hi = {loadUnit_maskInput_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_lo};
  wire [8191:0]       loadUnit_maskInput_hi_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_lo};
  wire [63:0]         _GEN_895 = {v0_1793, v0_1792};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo_lo = _GEN_895;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo_lo = _GEN_895;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo_lo = _GEN_895;
  wire [63:0]         _GEN_896 = {v0_1795, v0_1794};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo_hi = _GEN_896;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo_hi = _GEN_896;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo_hi = _GEN_896;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo = {loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_897 = {v0_1797, v0_1796};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi_lo = _GEN_897;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi_lo = _GEN_897;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi_lo = _GEN_897;
  wire [63:0]         _GEN_898 = {v0_1799, v0_1798};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi_hi = _GEN_898;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi_hi = _GEN_898;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi_hi = _GEN_898;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi = {loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo = {loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_899 = {v0_1801, v0_1800};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo_lo = _GEN_899;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo_lo = _GEN_899;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo_lo = _GEN_899;
  wire [63:0]         _GEN_900 = {v0_1803, v0_1802};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo_hi = _GEN_900;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo_hi = _GEN_900;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo_hi = _GEN_900;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo = {loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_901 = {v0_1805, v0_1804};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi_lo = _GEN_901;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi_lo = _GEN_901;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi_lo = _GEN_901;
  wire [63:0]         _GEN_902 = {v0_1807, v0_1806};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi_hi = _GEN_902;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi_hi = _GEN_902;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi_hi = _GEN_902;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi = {loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi = {loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo = {loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_903 = {v0_1809, v0_1808};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo_lo = _GEN_903;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo_lo = _GEN_903;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo_lo = _GEN_903;
  wire [63:0]         _GEN_904 = {v0_1811, v0_1810};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo_hi = _GEN_904;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo_hi = _GEN_904;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo_hi = _GEN_904;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo = {loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_905 = {v0_1813, v0_1812};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi_lo = _GEN_905;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi_lo = _GEN_905;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi_lo = _GEN_905;
  wire [63:0]         _GEN_906 = {v0_1815, v0_1814};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi_hi = _GEN_906;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi_hi = _GEN_906;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi_hi = _GEN_906;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi = {loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo = {loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_907 = {v0_1817, v0_1816};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo_lo = _GEN_907;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo_lo = _GEN_907;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo_lo = _GEN_907;
  wire [63:0]         _GEN_908 = {v0_1819, v0_1818};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo_hi = _GEN_908;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo_hi = _GEN_908;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo_hi = _GEN_908;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo = {loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_909 = {v0_1821, v0_1820};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi_lo = _GEN_909;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi_lo = _GEN_909;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi_lo = _GEN_909;
  wire [63:0]         _GEN_910 = {v0_1823, v0_1822};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi_hi = _GEN_910;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi_hi = _GEN_910;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi_hi = _GEN_910;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi = {loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi = {loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_hi_hi_lo_lo_lo = {loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_911 = {v0_1825, v0_1824};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo_lo = _GEN_911;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo_lo = _GEN_911;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo_lo = _GEN_911;
  wire [63:0]         _GEN_912 = {v0_1827, v0_1826};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo_hi = _GEN_912;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo_hi = _GEN_912;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo_hi = _GEN_912;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo = {loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_913 = {v0_1829, v0_1828};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi_lo = _GEN_913;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi_lo = _GEN_913;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi_lo = _GEN_913;
  wire [63:0]         _GEN_914 = {v0_1831, v0_1830};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi_hi = _GEN_914;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi_hi = _GEN_914;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi_hi = _GEN_914;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi = {loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo = {loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_915 = {v0_1833, v0_1832};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo_lo = _GEN_915;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo_lo = _GEN_915;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo_lo = _GEN_915;
  wire [63:0]         _GEN_916 = {v0_1835, v0_1834};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo_hi = _GEN_916;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo_hi = _GEN_916;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo_hi = _GEN_916;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo = {loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_917 = {v0_1837, v0_1836};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi_lo = _GEN_917;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi_lo = _GEN_917;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi_lo = _GEN_917;
  wire [63:0]         _GEN_918 = {v0_1839, v0_1838};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi_hi = _GEN_918;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi_hi = _GEN_918;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi_hi = _GEN_918;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi = {loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi = {loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo = {loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_919 = {v0_1841, v0_1840};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo_lo = _GEN_919;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo_lo = _GEN_919;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo_lo = _GEN_919;
  wire [63:0]         _GEN_920 = {v0_1843, v0_1842};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo_hi = _GEN_920;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo_hi = _GEN_920;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo_hi = _GEN_920;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo = {loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_921 = {v0_1845, v0_1844};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi_lo = _GEN_921;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi_lo = _GEN_921;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi_lo = _GEN_921;
  wire [63:0]         _GEN_922 = {v0_1847, v0_1846};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi_hi = _GEN_922;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi_hi = _GEN_922;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi_hi = _GEN_922;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi = {loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo = {loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_923 = {v0_1849, v0_1848};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo_lo = _GEN_923;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo_lo = _GEN_923;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo_lo = _GEN_923;
  wire [63:0]         _GEN_924 = {v0_1851, v0_1850};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo_hi = _GEN_924;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo_hi = _GEN_924;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo_hi = _GEN_924;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo = {loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_925 = {v0_1853, v0_1852};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi_lo = _GEN_925;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi_lo = _GEN_925;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi_lo = _GEN_925;
  wire [63:0]         _GEN_926 = {v0_1855, v0_1854};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi_hi = _GEN_926;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi_hi = _GEN_926;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi_hi = _GEN_926;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi = {loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_hi_hi_lo_lo_hi = {loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo};
  wire [2047:0]       loadUnit_maskInput_hi_hi_hi_lo_lo = {loadUnit_maskInput_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_927 = {v0_1857, v0_1856};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo_lo = _GEN_927;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo_lo = _GEN_927;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo_lo = _GEN_927;
  wire [63:0]         _GEN_928 = {v0_1859, v0_1858};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo_hi = _GEN_928;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo_hi = _GEN_928;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo_hi = _GEN_928;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo = {loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_929 = {v0_1861, v0_1860};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi_lo = _GEN_929;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi_lo = _GEN_929;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi_lo = _GEN_929;
  wire [63:0]         _GEN_930 = {v0_1863, v0_1862};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi_hi = _GEN_930;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi_hi = _GEN_930;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi_hi = _GEN_930;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi = {loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo = {loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_931 = {v0_1865, v0_1864};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo_lo = _GEN_931;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo_lo = _GEN_931;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo_lo = _GEN_931;
  wire [63:0]         _GEN_932 = {v0_1867, v0_1866};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo_hi = _GEN_932;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo_hi = _GEN_932;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo_hi = _GEN_932;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo = {loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_933 = {v0_1869, v0_1868};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi_lo = _GEN_933;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi_lo = _GEN_933;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi_lo = _GEN_933;
  wire [63:0]         _GEN_934 = {v0_1871, v0_1870};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi_hi = _GEN_934;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi_hi = _GEN_934;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi_hi = _GEN_934;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi = {loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi = {loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo = {loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_935 = {v0_1873, v0_1872};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo_lo = _GEN_935;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo_lo = _GEN_935;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo_lo = _GEN_935;
  wire [63:0]         _GEN_936 = {v0_1875, v0_1874};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo_hi = _GEN_936;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo_hi = _GEN_936;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo_hi = _GEN_936;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo = {loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_937 = {v0_1877, v0_1876};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi_lo = _GEN_937;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi_lo = _GEN_937;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi_lo = _GEN_937;
  wire [63:0]         _GEN_938 = {v0_1879, v0_1878};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi_hi = _GEN_938;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi_hi = _GEN_938;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi_hi = _GEN_938;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi = {loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo = {loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_939 = {v0_1881, v0_1880};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo_lo = _GEN_939;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo_lo = _GEN_939;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo_lo = _GEN_939;
  wire [63:0]         _GEN_940 = {v0_1883, v0_1882};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo_hi = _GEN_940;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo_hi = _GEN_940;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo_hi = _GEN_940;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo = {loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_941 = {v0_1885, v0_1884};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi_lo = _GEN_941;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi_lo = _GEN_941;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi_lo = _GEN_941;
  wire [63:0]         _GEN_942 = {v0_1887, v0_1886};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi_hi = _GEN_942;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi_hi = _GEN_942;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi_hi = _GEN_942;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi = {loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi = {loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_hi_hi_lo_hi_lo = {loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_943 = {v0_1889, v0_1888};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo_lo = _GEN_943;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo_lo = _GEN_943;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo_lo = _GEN_943;
  wire [63:0]         _GEN_944 = {v0_1891, v0_1890};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo_hi = _GEN_944;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo_hi = _GEN_944;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo_hi = _GEN_944;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo = {loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_945 = {v0_1893, v0_1892};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi_lo = _GEN_945;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi_lo = _GEN_945;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi_lo = _GEN_945;
  wire [63:0]         _GEN_946 = {v0_1895, v0_1894};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi_hi = _GEN_946;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi_hi = _GEN_946;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi_hi = _GEN_946;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi = {loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo = {loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_947 = {v0_1897, v0_1896};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo_lo = _GEN_947;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo_lo = _GEN_947;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo_lo = _GEN_947;
  wire [63:0]         _GEN_948 = {v0_1899, v0_1898};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo_hi = _GEN_948;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo_hi = _GEN_948;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo_hi = _GEN_948;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo = {loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_949 = {v0_1901, v0_1900};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi_lo = _GEN_949;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi_lo = _GEN_949;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi_lo = _GEN_949;
  wire [63:0]         _GEN_950 = {v0_1903, v0_1902};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi_hi = _GEN_950;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi_hi = _GEN_950;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi_hi = _GEN_950;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi = {loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi = {loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo = {loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_951 = {v0_1905, v0_1904};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo_lo = _GEN_951;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo_lo = _GEN_951;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo_lo = _GEN_951;
  wire [63:0]         _GEN_952 = {v0_1907, v0_1906};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo_hi = _GEN_952;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo_hi = _GEN_952;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo_hi = _GEN_952;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo = {loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_953 = {v0_1909, v0_1908};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi_lo = _GEN_953;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi_lo = _GEN_953;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi_lo = _GEN_953;
  wire [63:0]         _GEN_954 = {v0_1911, v0_1910};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi_hi = _GEN_954;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi_hi = _GEN_954;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi_hi = _GEN_954;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi = {loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo = {loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_955 = {v0_1913, v0_1912};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo_lo = _GEN_955;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo_lo = _GEN_955;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo_lo = _GEN_955;
  wire [63:0]         _GEN_956 = {v0_1915, v0_1914};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo_hi = _GEN_956;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo_hi = _GEN_956;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo_hi = _GEN_956;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo = {loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_957 = {v0_1917, v0_1916};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi_lo = _GEN_957;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi_lo = _GEN_957;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi_lo = _GEN_957;
  wire [63:0]         _GEN_958 = {v0_1919, v0_1918};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi_hi = _GEN_958;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi_hi = _GEN_958;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi_hi = _GEN_958;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_hi_hi_lo_hi_hi = {loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo};
  wire [2047:0]       loadUnit_maskInput_hi_hi_hi_lo_hi = {loadUnit_maskInput_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_lo};
  wire [4095:0]       loadUnit_maskInput_hi_hi_hi_lo = {loadUnit_maskInput_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_959 = {v0_1921, v0_1920};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo_lo = _GEN_959;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo_lo = _GEN_959;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo_lo = _GEN_959;
  wire [63:0]         _GEN_960 = {v0_1923, v0_1922};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo_hi = _GEN_960;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo_hi = _GEN_960;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo_hi = _GEN_960;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo = {loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_961 = {v0_1925, v0_1924};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi_lo = _GEN_961;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi_lo = _GEN_961;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi_lo = _GEN_961;
  wire [63:0]         _GEN_962 = {v0_1927, v0_1926};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi_hi = _GEN_962;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi_hi = _GEN_962;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi_hi = _GEN_962;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi = {loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo = {loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_963 = {v0_1929, v0_1928};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo_lo = _GEN_963;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo_lo = _GEN_963;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo_lo = _GEN_963;
  wire [63:0]         _GEN_964 = {v0_1931, v0_1930};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo_hi = _GEN_964;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo_hi = _GEN_964;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo_hi = _GEN_964;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo = {loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_965 = {v0_1933, v0_1932};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi_lo = _GEN_965;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi_lo = _GEN_965;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi_lo = _GEN_965;
  wire [63:0]         _GEN_966 = {v0_1935, v0_1934};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi_hi = _GEN_966;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi_hi = _GEN_966;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi_hi = _GEN_966;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi = {loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo = {loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_967 = {v0_1937, v0_1936};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo_lo = _GEN_967;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo_lo = _GEN_967;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo_lo = _GEN_967;
  wire [63:0]         _GEN_968 = {v0_1939, v0_1938};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo_hi = _GEN_968;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo_hi = _GEN_968;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo_hi = _GEN_968;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo = {loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_969 = {v0_1941, v0_1940};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi_lo = _GEN_969;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi_lo = _GEN_969;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi_lo = _GEN_969;
  wire [63:0]         _GEN_970 = {v0_1943, v0_1942};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi_hi = _GEN_970;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi_hi = _GEN_970;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi_hi = _GEN_970;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi = {loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo = {loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_971 = {v0_1945, v0_1944};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo_lo = _GEN_971;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo_lo = _GEN_971;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo_lo = _GEN_971;
  wire [63:0]         _GEN_972 = {v0_1947, v0_1946};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo_hi = _GEN_972;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo_hi = _GEN_972;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo_hi = _GEN_972;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo = {loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_973 = {v0_1949, v0_1948};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi_lo = _GEN_973;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi_lo = _GEN_973;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi_lo = _GEN_973;
  wire [63:0]         _GEN_974 = {v0_1951, v0_1950};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi_hi = _GEN_974;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi_hi = _GEN_974;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi_hi = _GEN_974;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi = {loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_hi_hi_hi_lo_lo = {loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_975 = {v0_1953, v0_1952};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo_lo = _GEN_975;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo_lo = _GEN_975;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo_lo = _GEN_975;
  wire [63:0]         _GEN_976 = {v0_1955, v0_1954};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo_hi = _GEN_976;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo_hi = _GEN_976;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo_hi = _GEN_976;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo = {loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_977 = {v0_1957, v0_1956};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi_lo = _GEN_977;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi_lo = _GEN_977;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi_lo = _GEN_977;
  wire [63:0]         _GEN_978 = {v0_1959, v0_1958};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi_hi = _GEN_978;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi_hi = _GEN_978;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi_hi = _GEN_978;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi = {loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo = {loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_979 = {v0_1961, v0_1960};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo_lo = _GEN_979;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo_lo = _GEN_979;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo_lo = _GEN_979;
  wire [63:0]         _GEN_980 = {v0_1963, v0_1962};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo_hi = _GEN_980;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo_hi = _GEN_980;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo_hi = _GEN_980;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo = {loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_981 = {v0_1965, v0_1964};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi_lo = _GEN_981;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi_lo = _GEN_981;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi_lo = _GEN_981;
  wire [63:0]         _GEN_982 = {v0_1967, v0_1966};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi_hi = _GEN_982;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi_hi = _GEN_982;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi_hi = _GEN_982;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi = {loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo = {loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_983 = {v0_1969, v0_1968};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo_lo = _GEN_983;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo_lo = _GEN_983;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo_lo = _GEN_983;
  wire [63:0]         _GEN_984 = {v0_1971, v0_1970};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo_hi = _GEN_984;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo_hi = _GEN_984;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo_hi = _GEN_984;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo = {loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_985 = {v0_1973, v0_1972};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi_lo = _GEN_985;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi_lo = _GEN_985;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi_lo = _GEN_985;
  wire [63:0]         _GEN_986 = {v0_1975, v0_1974};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi_hi = _GEN_986;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi_hi = _GEN_986;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi_hi = _GEN_986;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi = {loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo = {loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_987 = {v0_1977, v0_1976};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo_lo = _GEN_987;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo_lo = _GEN_987;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo_lo = _GEN_987;
  wire [63:0]         _GEN_988 = {v0_1979, v0_1978};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo_hi = _GEN_988;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo_hi = _GEN_988;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo_hi = _GEN_988;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo = {loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_989 = {v0_1981, v0_1980};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi_lo = _GEN_989;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi_lo = _GEN_989;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi_lo = _GEN_989;
  wire [63:0]         _GEN_990 = {v0_1983, v0_1982};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi_hi = _GEN_990;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi_hi = _GEN_990;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi_hi = _GEN_990;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_hi_hi_hi_lo_hi = {loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo};
  wire [2047:0]       loadUnit_maskInput_hi_hi_hi_hi_lo = {loadUnit_maskInput_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_991 = {v0_1985, v0_1984};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo_lo = _GEN_991;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo_lo = _GEN_991;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo_lo = _GEN_991;
  wire [63:0]         _GEN_992 = {v0_1987, v0_1986};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo_hi = _GEN_992;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo_hi = _GEN_992;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo_hi = _GEN_992;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo = {loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_993 = {v0_1989, v0_1988};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi_lo = _GEN_993;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi_lo = _GEN_993;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi_lo = _GEN_993;
  wire [63:0]         _GEN_994 = {v0_1991, v0_1990};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi_hi = _GEN_994;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi_hi = _GEN_994;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi_hi = _GEN_994;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi = {loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo = {loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_995 = {v0_1993, v0_1992};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo_lo = _GEN_995;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo_lo = _GEN_995;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo_lo = _GEN_995;
  wire [63:0]         _GEN_996 = {v0_1995, v0_1994};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo_hi = _GEN_996;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo_hi = _GEN_996;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo_hi = _GEN_996;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo = {loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_997 = {v0_1997, v0_1996};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi_lo = _GEN_997;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi_lo = _GEN_997;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi_lo = _GEN_997;
  wire [63:0]         _GEN_998 = {v0_1999, v0_1998};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi_hi = _GEN_998;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi_hi = _GEN_998;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi_hi = _GEN_998;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi = {loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo = {loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_999 = {v0_2001, v0_2000};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo_lo = _GEN_999;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo_lo = _GEN_999;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo_lo = _GEN_999;
  wire [63:0]         _GEN_1000 = {v0_2003, v0_2002};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo_hi = _GEN_1000;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo_hi = _GEN_1000;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo_hi = _GEN_1000;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo = {loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_1001 = {v0_2005, v0_2004};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi_lo = _GEN_1001;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi_lo = _GEN_1001;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi_lo = _GEN_1001;
  wire [63:0]         _GEN_1002 = {v0_2007, v0_2006};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi_hi = _GEN_1002;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi_hi = _GEN_1002;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi_hi = _GEN_1002;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi = {loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo = {loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_1003 = {v0_2009, v0_2008};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo_lo = _GEN_1003;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo_lo = _GEN_1003;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo_lo = _GEN_1003;
  wire [63:0]         _GEN_1004 = {v0_2011, v0_2010};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo_hi = _GEN_1004;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo_hi = _GEN_1004;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo_hi = _GEN_1004;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo = {loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_1005 = {v0_2013, v0_2012};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi_lo = _GEN_1005;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi_lo = _GEN_1005;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi_lo = _GEN_1005;
  wire [63:0]         _GEN_1006 = {v0_2015, v0_2014};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi_hi = _GEN_1006;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi_hi = _GEN_1006;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi_hi = _GEN_1006;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi = {loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_hi_hi_hi_hi_lo = {loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_1007 = {v0_2017, v0_2016};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo_lo = _GEN_1007;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo_lo = _GEN_1007;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo_lo = _GEN_1007;
  wire [63:0]         _GEN_1008 = {v0_2019, v0_2018};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo_hi = _GEN_1008;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo_hi = _GEN_1008;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo_hi = _GEN_1008;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo = {loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_1009 = {v0_2021, v0_2020};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi_lo = _GEN_1009;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi_lo = _GEN_1009;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi_lo = _GEN_1009;
  wire [63:0]         _GEN_1010 = {v0_2023, v0_2022};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi_hi = _GEN_1010;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi_hi = _GEN_1010;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi_hi = _GEN_1010;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi = {loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo = {loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_1011 = {v0_2025, v0_2024};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo_lo = _GEN_1011;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo_lo = _GEN_1011;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo_lo = _GEN_1011;
  wire [63:0]         _GEN_1012 = {v0_2027, v0_2026};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo_hi = _GEN_1012;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo_hi = _GEN_1012;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo_hi = _GEN_1012;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo = {loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_1013 = {v0_2029, v0_2028};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi_lo = _GEN_1013;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi_lo = _GEN_1013;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi_lo = _GEN_1013;
  wire [63:0]         _GEN_1014 = {v0_2031, v0_2030};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi_hi = _GEN_1014;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi_hi = _GEN_1014;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi_hi = _GEN_1014;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi = {loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo = {loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_1015 = {v0_2033, v0_2032};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo_lo = _GEN_1015;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo_lo = _GEN_1015;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo_lo = _GEN_1015;
  wire [63:0]         _GEN_1016 = {v0_2035, v0_2034};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo_hi = _GEN_1016;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo_hi = _GEN_1016;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo_hi = _GEN_1016;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo = {loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_1017 = {v0_2037, v0_2036};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi_lo = _GEN_1017;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi_lo = _GEN_1017;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi_lo = _GEN_1017;
  wire [63:0]         _GEN_1018 = {v0_2039, v0_2038};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi_hi = _GEN_1018;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi_hi = _GEN_1018;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi_hi = _GEN_1018;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi = {loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo = {loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_1019 = {v0_2041, v0_2040};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo_lo = _GEN_1019;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo_lo = _GEN_1019;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo_lo = _GEN_1019;
  wire [63:0]         _GEN_1020 = {v0_2043, v0_2042};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo_hi = _GEN_1020;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo_hi = _GEN_1020;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo_hi = _GEN_1020;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo = {loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_1021 = {v0_2045, v0_2044};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi_lo = _GEN_1021;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi_lo = _GEN_1021;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi_lo = _GEN_1021;
  wire [63:0]         _GEN_1022 = {v0_2047, v0_2046};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi_hi = _GEN_1022;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi_hi = _GEN_1022;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi_hi = _GEN_1022;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_hi_hi_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo};
  wire [2047:0]       loadUnit_maskInput_hi_hi_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_lo};
  wire [4095:0]       loadUnit_maskInput_hi_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_lo};
  wire [8191:0]       loadUnit_maskInput_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_lo};
  wire [16383:0]      loadUnit_maskInput_hi_hi = {loadUnit_maskInput_hi_hi_hi, loadUnit_maskInput_hi_hi_lo};
  wire [32767:0]      loadUnit_maskInput_hi = {loadUnit_maskInput_hi_hi, loadUnit_maskInput_hi_lo};
  wire [4095:0][15:0] _GEN_1023 =
    {{loadUnit_maskInput_hi[32767:32752]},
     {loadUnit_maskInput_hi[32751:32736]},
     {loadUnit_maskInput_hi[32735:32720]},
     {loadUnit_maskInput_hi[32719:32704]},
     {loadUnit_maskInput_hi[32703:32688]},
     {loadUnit_maskInput_hi[32687:32672]},
     {loadUnit_maskInput_hi[32671:32656]},
     {loadUnit_maskInput_hi[32655:32640]},
     {loadUnit_maskInput_hi[32639:32624]},
     {loadUnit_maskInput_hi[32623:32608]},
     {loadUnit_maskInput_hi[32607:32592]},
     {loadUnit_maskInput_hi[32591:32576]},
     {loadUnit_maskInput_hi[32575:32560]},
     {loadUnit_maskInput_hi[32559:32544]},
     {loadUnit_maskInput_hi[32543:32528]},
     {loadUnit_maskInput_hi[32527:32512]},
     {loadUnit_maskInput_hi[32511:32496]},
     {loadUnit_maskInput_hi[32495:32480]},
     {loadUnit_maskInput_hi[32479:32464]},
     {loadUnit_maskInput_hi[32463:32448]},
     {loadUnit_maskInput_hi[32447:32432]},
     {loadUnit_maskInput_hi[32431:32416]},
     {loadUnit_maskInput_hi[32415:32400]},
     {loadUnit_maskInput_hi[32399:32384]},
     {loadUnit_maskInput_hi[32383:32368]},
     {loadUnit_maskInput_hi[32367:32352]},
     {loadUnit_maskInput_hi[32351:32336]},
     {loadUnit_maskInput_hi[32335:32320]},
     {loadUnit_maskInput_hi[32319:32304]},
     {loadUnit_maskInput_hi[32303:32288]},
     {loadUnit_maskInput_hi[32287:32272]},
     {loadUnit_maskInput_hi[32271:32256]},
     {loadUnit_maskInput_hi[32255:32240]},
     {loadUnit_maskInput_hi[32239:32224]},
     {loadUnit_maskInput_hi[32223:32208]},
     {loadUnit_maskInput_hi[32207:32192]},
     {loadUnit_maskInput_hi[32191:32176]},
     {loadUnit_maskInput_hi[32175:32160]},
     {loadUnit_maskInput_hi[32159:32144]},
     {loadUnit_maskInput_hi[32143:32128]},
     {loadUnit_maskInput_hi[32127:32112]},
     {loadUnit_maskInput_hi[32111:32096]},
     {loadUnit_maskInput_hi[32095:32080]},
     {loadUnit_maskInput_hi[32079:32064]},
     {loadUnit_maskInput_hi[32063:32048]},
     {loadUnit_maskInput_hi[32047:32032]},
     {loadUnit_maskInput_hi[32031:32016]},
     {loadUnit_maskInput_hi[32015:32000]},
     {loadUnit_maskInput_hi[31999:31984]},
     {loadUnit_maskInput_hi[31983:31968]},
     {loadUnit_maskInput_hi[31967:31952]},
     {loadUnit_maskInput_hi[31951:31936]},
     {loadUnit_maskInput_hi[31935:31920]},
     {loadUnit_maskInput_hi[31919:31904]},
     {loadUnit_maskInput_hi[31903:31888]},
     {loadUnit_maskInput_hi[31887:31872]},
     {loadUnit_maskInput_hi[31871:31856]},
     {loadUnit_maskInput_hi[31855:31840]},
     {loadUnit_maskInput_hi[31839:31824]},
     {loadUnit_maskInput_hi[31823:31808]},
     {loadUnit_maskInput_hi[31807:31792]},
     {loadUnit_maskInput_hi[31791:31776]},
     {loadUnit_maskInput_hi[31775:31760]},
     {loadUnit_maskInput_hi[31759:31744]},
     {loadUnit_maskInput_hi[31743:31728]},
     {loadUnit_maskInput_hi[31727:31712]},
     {loadUnit_maskInput_hi[31711:31696]},
     {loadUnit_maskInput_hi[31695:31680]},
     {loadUnit_maskInput_hi[31679:31664]},
     {loadUnit_maskInput_hi[31663:31648]},
     {loadUnit_maskInput_hi[31647:31632]},
     {loadUnit_maskInput_hi[31631:31616]},
     {loadUnit_maskInput_hi[31615:31600]},
     {loadUnit_maskInput_hi[31599:31584]},
     {loadUnit_maskInput_hi[31583:31568]},
     {loadUnit_maskInput_hi[31567:31552]},
     {loadUnit_maskInput_hi[31551:31536]},
     {loadUnit_maskInput_hi[31535:31520]},
     {loadUnit_maskInput_hi[31519:31504]},
     {loadUnit_maskInput_hi[31503:31488]},
     {loadUnit_maskInput_hi[31487:31472]},
     {loadUnit_maskInput_hi[31471:31456]},
     {loadUnit_maskInput_hi[31455:31440]},
     {loadUnit_maskInput_hi[31439:31424]},
     {loadUnit_maskInput_hi[31423:31408]},
     {loadUnit_maskInput_hi[31407:31392]},
     {loadUnit_maskInput_hi[31391:31376]},
     {loadUnit_maskInput_hi[31375:31360]},
     {loadUnit_maskInput_hi[31359:31344]},
     {loadUnit_maskInput_hi[31343:31328]},
     {loadUnit_maskInput_hi[31327:31312]},
     {loadUnit_maskInput_hi[31311:31296]},
     {loadUnit_maskInput_hi[31295:31280]},
     {loadUnit_maskInput_hi[31279:31264]},
     {loadUnit_maskInput_hi[31263:31248]},
     {loadUnit_maskInput_hi[31247:31232]},
     {loadUnit_maskInput_hi[31231:31216]},
     {loadUnit_maskInput_hi[31215:31200]},
     {loadUnit_maskInput_hi[31199:31184]},
     {loadUnit_maskInput_hi[31183:31168]},
     {loadUnit_maskInput_hi[31167:31152]},
     {loadUnit_maskInput_hi[31151:31136]},
     {loadUnit_maskInput_hi[31135:31120]},
     {loadUnit_maskInput_hi[31119:31104]},
     {loadUnit_maskInput_hi[31103:31088]},
     {loadUnit_maskInput_hi[31087:31072]},
     {loadUnit_maskInput_hi[31071:31056]},
     {loadUnit_maskInput_hi[31055:31040]},
     {loadUnit_maskInput_hi[31039:31024]},
     {loadUnit_maskInput_hi[31023:31008]},
     {loadUnit_maskInput_hi[31007:30992]},
     {loadUnit_maskInput_hi[30991:30976]},
     {loadUnit_maskInput_hi[30975:30960]},
     {loadUnit_maskInput_hi[30959:30944]},
     {loadUnit_maskInput_hi[30943:30928]},
     {loadUnit_maskInput_hi[30927:30912]},
     {loadUnit_maskInput_hi[30911:30896]},
     {loadUnit_maskInput_hi[30895:30880]},
     {loadUnit_maskInput_hi[30879:30864]},
     {loadUnit_maskInput_hi[30863:30848]},
     {loadUnit_maskInput_hi[30847:30832]},
     {loadUnit_maskInput_hi[30831:30816]},
     {loadUnit_maskInput_hi[30815:30800]},
     {loadUnit_maskInput_hi[30799:30784]},
     {loadUnit_maskInput_hi[30783:30768]},
     {loadUnit_maskInput_hi[30767:30752]},
     {loadUnit_maskInput_hi[30751:30736]},
     {loadUnit_maskInput_hi[30735:30720]},
     {loadUnit_maskInput_hi[30719:30704]},
     {loadUnit_maskInput_hi[30703:30688]},
     {loadUnit_maskInput_hi[30687:30672]},
     {loadUnit_maskInput_hi[30671:30656]},
     {loadUnit_maskInput_hi[30655:30640]},
     {loadUnit_maskInput_hi[30639:30624]},
     {loadUnit_maskInput_hi[30623:30608]},
     {loadUnit_maskInput_hi[30607:30592]},
     {loadUnit_maskInput_hi[30591:30576]},
     {loadUnit_maskInput_hi[30575:30560]},
     {loadUnit_maskInput_hi[30559:30544]},
     {loadUnit_maskInput_hi[30543:30528]},
     {loadUnit_maskInput_hi[30527:30512]},
     {loadUnit_maskInput_hi[30511:30496]},
     {loadUnit_maskInput_hi[30495:30480]},
     {loadUnit_maskInput_hi[30479:30464]},
     {loadUnit_maskInput_hi[30463:30448]},
     {loadUnit_maskInput_hi[30447:30432]},
     {loadUnit_maskInput_hi[30431:30416]},
     {loadUnit_maskInput_hi[30415:30400]},
     {loadUnit_maskInput_hi[30399:30384]},
     {loadUnit_maskInput_hi[30383:30368]},
     {loadUnit_maskInput_hi[30367:30352]},
     {loadUnit_maskInput_hi[30351:30336]},
     {loadUnit_maskInput_hi[30335:30320]},
     {loadUnit_maskInput_hi[30319:30304]},
     {loadUnit_maskInput_hi[30303:30288]},
     {loadUnit_maskInput_hi[30287:30272]},
     {loadUnit_maskInput_hi[30271:30256]},
     {loadUnit_maskInput_hi[30255:30240]},
     {loadUnit_maskInput_hi[30239:30224]},
     {loadUnit_maskInput_hi[30223:30208]},
     {loadUnit_maskInput_hi[30207:30192]},
     {loadUnit_maskInput_hi[30191:30176]},
     {loadUnit_maskInput_hi[30175:30160]},
     {loadUnit_maskInput_hi[30159:30144]},
     {loadUnit_maskInput_hi[30143:30128]},
     {loadUnit_maskInput_hi[30127:30112]},
     {loadUnit_maskInput_hi[30111:30096]},
     {loadUnit_maskInput_hi[30095:30080]},
     {loadUnit_maskInput_hi[30079:30064]},
     {loadUnit_maskInput_hi[30063:30048]},
     {loadUnit_maskInput_hi[30047:30032]},
     {loadUnit_maskInput_hi[30031:30016]},
     {loadUnit_maskInput_hi[30015:30000]},
     {loadUnit_maskInput_hi[29999:29984]},
     {loadUnit_maskInput_hi[29983:29968]},
     {loadUnit_maskInput_hi[29967:29952]},
     {loadUnit_maskInput_hi[29951:29936]},
     {loadUnit_maskInput_hi[29935:29920]},
     {loadUnit_maskInput_hi[29919:29904]},
     {loadUnit_maskInput_hi[29903:29888]},
     {loadUnit_maskInput_hi[29887:29872]},
     {loadUnit_maskInput_hi[29871:29856]},
     {loadUnit_maskInput_hi[29855:29840]},
     {loadUnit_maskInput_hi[29839:29824]},
     {loadUnit_maskInput_hi[29823:29808]},
     {loadUnit_maskInput_hi[29807:29792]},
     {loadUnit_maskInput_hi[29791:29776]},
     {loadUnit_maskInput_hi[29775:29760]},
     {loadUnit_maskInput_hi[29759:29744]},
     {loadUnit_maskInput_hi[29743:29728]},
     {loadUnit_maskInput_hi[29727:29712]},
     {loadUnit_maskInput_hi[29711:29696]},
     {loadUnit_maskInput_hi[29695:29680]},
     {loadUnit_maskInput_hi[29679:29664]},
     {loadUnit_maskInput_hi[29663:29648]},
     {loadUnit_maskInput_hi[29647:29632]},
     {loadUnit_maskInput_hi[29631:29616]},
     {loadUnit_maskInput_hi[29615:29600]},
     {loadUnit_maskInput_hi[29599:29584]},
     {loadUnit_maskInput_hi[29583:29568]},
     {loadUnit_maskInput_hi[29567:29552]},
     {loadUnit_maskInput_hi[29551:29536]},
     {loadUnit_maskInput_hi[29535:29520]},
     {loadUnit_maskInput_hi[29519:29504]},
     {loadUnit_maskInput_hi[29503:29488]},
     {loadUnit_maskInput_hi[29487:29472]},
     {loadUnit_maskInput_hi[29471:29456]},
     {loadUnit_maskInput_hi[29455:29440]},
     {loadUnit_maskInput_hi[29439:29424]},
     {loadUnit_maskInput_hi[29423:29408]},
     {loadUnit_maskInput_hi[29407:29392]},
     {loadUnit_maskInput_hi[29391:29376]},
     {loadUnit_maskInput_hi[29375:29360]},
     {loadUnit_maskInput_hi[29359:29344]},
     {loadUnit_maskInput_hi[29343:29328]},
     {loadUnit_maskInput_hi[29327:29312]},
     {loadUnit_maskInput_hi[29311:29296]},
     {loadUnit_maskInput_hi[29295:29280]},
     {loadUnit_maskInput_hi[29279:29264]},
     {loadUnit_maskInput_hi[29263:29248]},
     {loadUnit_maskInput_hi[29247:29232]},
     {loadUnit_maskInput_hi[29231:29216]},
     {loadUnit_maskInput_hi[29215:29200]},
     {loadUnit_maskInput_hi[29199:29184]},
     {loadUnit_maskInput_hi[29183:29168]},
     {loadUnit_maskInput_hi[29167:29152]},
     {loadUnit_maskInput_hi[29151:29136]},
     {loadUnit_maskInput_hi[29135:29120]},
     {loadUnit_maskInput_hi[29119:29104]},
     {loadUnit_maskInput_hi[29103:29088]},
     {loadUnit_maskInput_hi[29087:29072]},
     {loadUnit_maskInput_hi[29071:29056]},
     {loadUnit_maskInput_hi[29055:29040]},
     {loadUnit_maskInput_hi[29039:29024]},
     {loadUnit_maskInput_hi[29023:29008]},
     {loadUnit_maskInput_hi[29007:28992]},
     {loadUnit_maskInput_hi[28991:28976]},
     {loadUnit_maskInput_hi[28975:28960]},
     {loadUnit_maskInput_hi[28959:28944]},
     {loadUnit_maskInput_hi[28943:28928]},
     {loadUnit_maskInput_hi[28927:28912]},
     {loadUnit_maskInput_hi[28911:28896]},
     {loadUnit_maskInput_hi[28895:28880]},
     {loadUnit_maskInput_hi[28879:28864]},
     {loadUnit_maskInput_hi[28863:28848]},
     {loadUnit_maskInput_hi[28847:28832]},
     {loadUnit_maskInput_hi[28831:28816]},
     {loadUnit_maskInput_hi[28815:28800]},
     {loadUnit_maskInput_hi[28799:28784]},
     {loadUnit_maskInput_hi[28783:28768]},
     {loadUnit_maskInput_hi[28767:28752]},
     {loadUnit_maskInput_hi[28751:28736]},
     {loadUnit_maskInput_hi[28735:28720]},
     {loadUnit_maskInput_hi[28719:28704]},
     {loadUnit_maskInput_hi[28703:28688]},
     {loadUnit_maskInput_hi[28687:28672]},
     {loadUnit_maskInput_hi[28671:28656]},
     {loadUnit_maskInput_hi[28655:28640]},
     {loadUnit_maskInput_hi[28639:28624]},
     {loadUnit_maskInput_hi[28623:28608]},
     {loadUnit_maskInput_hi[28607:28592]},
     {loadUnit_maskInput_hi[28591:28576]},
     {loadUnit_maskInput_hi[28575:28560]},
     {loadUnit_maskInput_hi[28559:28544]},
     {loadUnit_maskInput_hi[28543:28528]},
     {loadUnit_maskInput_hi[28527:28512]},
     {loadUnit_maskInput_hi[28511:28496]},
     {loadUnit_maskInput_hi[28495:28480]},
     {loadUnit_maskInput_hi[28479:28464]},
     {loadUnit_maskInput_hi[28463:28448]},
     {loadUnit_maskInput_hi[28447:28432]},
     {loadUnit_maskInput_hi[28431:28416]},
     {loadUnit_maskInput_hi[28415:28400]},
     {loadUnit_maskInput_hi[28399:28384]},
     {loadUnit_maskInput_hi[28383:28368]},
     {loadUnit_maskInput_hi[28367:28352]},
     {loadUnit_maskInput_hi[28351:28336]},
     {loadUnit_maskInput_hi[28335:28320]},
     {loadUnit_maskInput_hi[28319:28304]},
     {loadUnit_maskInput_hi[28303:28288]},
     {loadUnit_maskInput_hi[28287:28272]},
     {loadUnit_maskInput_hi[28271:28256]},
     {loadUnit_maskInput_hi[28255:28240]},
     {loadUnit_maskInput_hi[28239:28224]},
     {loadUnit_maskInput_hi[28223:28208]},
     {loadUnit_maskInput_hi[28207:28192]},
     {loadUnit_maskInput_hi[28191:28176]},
     {loadUnit_maskInput_hi[28175:28160]},
     {loadUnit_maskInput_hi[28159:28144]},
     {loadUnit_maskInput_hi[28143:28128]},
     {loadUnit_maskInput_hi[28127:28112]},
     {loadUnit_maskInput_hi[28111:28096]},
     {loadUnit_maskInput_hi[28095:28080]},
     {loadUnit_maskInput_hi[28079:28064]},
     {loadUnit_maskInput_hi[28063:28048]},
     {loadUnit_maskInput_hi[28047:28032]},
     {loadUnit_maskInput_hi[28031:28016]},
     {loadUnit_maskInput_hi[28015:28000]},
     {loadUnit_maskInput_hi[27999:27984]},
     {loadUnit_maskInput_hi[27983:27968]},
     {loadUnit_maskInput_hi[27967:27952]},
     {loadUnit_maskInput_hi[27951:27936]},
     {loadUnit_maskInput_hi[27935:27920]},
     {loadUnit_maskInput_hi[27919:27904]},
     {loadUnit_maskInput_hi[27903:27888]},
     {loadUnit_maskInput_hi[27887:27872]},
     {loadUnit_maskInput_hi[27871:27856]},
     {loadUnit_maskInput_hi[27855:27840]},
     {loadUnit_maskInput_hi[27839:27824]},
     {loadUnit_maskInput_hi[27823:27808]},
     {loadUnit_maskInput_hi[27807:27792]},
     {loadUnit_maskInput_hi[27791:27776]},
     {loadUnit_maskInput_hi[27775:27760]},
     {loadUnit_maskInput_hi[27759:27744]},
     {loadUnit_maskInput_hi[27743:27728]},
     {loadUnit_maskInput_hi[27727:27712]},
     {loadUnit_maskInput_hi[27711:27696]},
     {loadUnit_maskInput_hi[27695:27680]},
     {loadUnit_maskInput_hi[27679:27664]},
     {loadUnit_maskInput_hi[27663:27648]},
     {loadUnit_maskInput_hi[27647:27632]},
     {loadUnit_maskInput_hi[27631:27616]},
     {loadUnit_maskInput_hi[27615:27600]},
     {loadUnit_maskInput_hi[27599:27584]},
     {loadUnit_maskInput_hi[27583:27568]},
     {loadUnit_maskInput_hi[27567:27552]},
     {loadUnit_maskInput_hi[27551:27536]},
     {loadUnit_maskInput_hi[27535:27520]},
     {loadUnit_maskInput_hi[27519:27504]},
     {loadUnit_maskInput_hi[27503:27488]},
     {loadUnit_maskInput_hi[27487:27472]},
     {loadUnit_maskInput_hi[27471:27456]},
     {loadUnit_maskInput_hi[27455:27440]},
     {loadUnit_maskInput_hi[27439:27424]},
     {loadUnit_maskInput_hi[27423:27408]},
     {loadUnit_maskInput_hi[27407:27392]},
     {loadUnit_maskInput_hi[27391:27376]},
     {loadUnit_maskInput_hi[27375:27360]},
     {loadUnit_maskInput_hi[27359:27344]},
     {loadUnit_maskInput_hi[27343:27328]},
     {loadUnit_maskInput_hi[27327:27312]},
     {loadUnit_maskInput_hi[27311:27296]},
     {loadUnit_maskInput_hi[27295:27280]},
     {loadUnit_maskInput_hi[27279:27264]},
     {loadUnit_maskInput_hi[27263:27248]},
     {loadUnit_maskInput_hi[27247:27232]},
     {loadUnit_maskInput_hi[27231:27216]},
     {loadUnit_maskInput_hi[27215:27200]},
     {loadUnit_maskInput_hi[27199:27184]},
     {loadUnit_maskInput_hi[27183:27168]},
     {loadUnit_maskInput_hi[27167:27152]},
     {loadUnit_maskInput_hi[27151:27136]},
     {loadUnit_maskInput_hi[27135:27120]},
     {loadUnit_maskInput_hi[27119:27104]},
     {loadUnit_maskInput_hi[27103:27088]},
     {loadUnit_maskInput_hi[27087:27072]},
     {loadUnit_maskInput_hi[27071:27056]},
     {loadUnit_maskInput_hi[27055:27040]},
     {loadUnit_maskInput_hi[27039:27024]},
     {loadUnit_maskInput_hi[27023:27008]},
     {loadUnit_maskInput_hi[27007:26992]},
     {loadUnit_maskInput_hi[26991:26976]},
     {loadUnit_maskInput_hi[26975:26960]},
     {loadUnit_maskInput_hi[26959:26944]},
     {loadUnit_maskInput_hi[26943:26928]},
     {loadUnit_maskInput_hi[26927:26912]},
     {loadUnit_maskInput_hi[26911:26896]},
     {loadUnit_maskInput_hi[26895:26880]},
     {loadUnit_maskInput_hi[26879:26864]},
     {loadUnit_maskInput_hi[26863:26848]},
     {loadUnit_maskInput_hi[26847:26832]},
     {loadUnit_maskInput_hi[26831:26816]},
     {loadUnit_maskInput_hi[26815:26800]},
     {loadUnit_maskInput_hi[26799:26784]},
     {loadUnit_maskInput_hi[26783:26768]},
     {loadUnit_maskInput_hi[26767:26752]},
     {loadUnit_maskInput_hi[26751:26736]},
     {loadUnit_maskInput_hi[26735:26720]},
     {loadUnit_maskInput_hi[26719:26704]},
     {loadUnit_maskInput_hi[26703:26688]},
     {loadUnit_maskInput_hi[26687:26672]},
     {loadUnit_maskInput_hi[26671:26656]},
     {loadUnit_maskInput_hi[26655:26640]},
     {loadUnit_maskInput_hi[26639:26624]},
     {loadUnit_maskInput_hi[26623:26608]},
     {loadUnit_maskInput_hi[26607:26592]},
     {loadUnit_maskInput_hi[26591:26576]},
     {loadUnit_maskInput_hi[26575:26560]},
     {loadUnit_maskInput_hi[26559:26544]},
     {loadUnit_maskInput_hi[26543:26528]},
     {loadUnit_maskInput_hi[26527:26512]},
     {loadUnit_maskInput_hi[26511:26496]},
     {loadUnit_maskInput_hi[26495:26480]},
     {loadUnit_maskInput_hi[26479:26464]},
     {loadUnit_maskInput_hi[26463:26448]},
     {loadUnit_maskInput_hi[26447:26432]},
     {loadUnit_maskInput_hi[26431:26416]},
     {loadUnit_maskInput_hi[26415:26400]},
     {loadUnit_maskInput_hi[26399:26384]},
     {loadUnit_maskInput_hi[26383:26368]},
     {loadUnit_maskInput_hi[26367:26352]},
     {loadUnit_maskInput_hi[26351:26336]},
     {loadUnit_maskInput_hi[26335:26320]},
     {loadUnit_maskInput_hi[26319:26304]},
     {loadUnit_maskInput_hi[26303:26288]},
     {loadUnit_maskInput_hi[26287:26272]},
     {loadUnit_maskInput_hi[26271:26256]},
     {loadUnit_maskInput_hi[26255:26240]},
     {loadUnit_maskInput_hi[26239:26224]},
     {loadUnit_maskInput_hi[26223:26208]},
     {loadUnit_maskInput_hi[26207:26192]},
     {loadUnit_maskInput_hi[26191:26176]},
     {loadUnit_maskInput_hi[26175:26160]},
     {loadUnit_maskInput_hi[26159:26144]},
     {loadUnit_maskInput_hi[26143:26128]},
     {loadUnit_maskInput_hi[26127:26112]},
     {loadUnit_maskInput_hi[26111:26096]},
     {loadUnit_maskInput_hi[26095:26080]},
     {loadUnit_maskInput_hi[26079:26064]},
     {loadUnit_maskInput_hi[26063:26048]},
     {loadUnit_maskInput_hi[26047:26032]},
     {loadUnit_maskInput_hi[26031:26016]},
     {loadUnit_maskInput_hi[26015:26000]},
     {loadUnit_maskInput_hi[25999:25984]},
     {loadUnit_maskInput_hi[25983:25968]},
     {loadUnit_maskInput_hi[25967:25952]},
     {loadUnit_maskInput_hi[25951:25936]},
     {loadUnit_maskInput_hi[25935:25920]},
     {loadUnit_maskInput_hi[25919:25904]},
     {loadUnit_maskInput_hi[25903:25888]},
     {loadUnit_maskInput_hi[25887:25872]},
     {loadUnit_maskInput_hi[25871:25856]},
     {loadUnit_maskInput_hi[25855:25840]},
     {loadUnit_maskInput_hi[25839:25824]},
     {loadUnit_maskInput_hi[25823:25808]},
     {loadUnit_maskInput_hi[25807:25792]},
     {loadUnit_maskInput_hi[25791:25776]},
     {loadUnit_maskInput_hi[25775:25760]},
     {loadUnit_maskInput_hi[25759:25744]},
     {loadUnit_maskInput_hi[25743:25728]},
     {loadUnit_maskInput_hi[25727:25712]},
     {loadUnit_maskInput_hi[25711:25696]},
     {loadUnit_maskInput_hi[25695:25680]},
     {loadUnit_maskInput_hi[25679:25664]},
     {loadUnit_maskInput_hi[25663:25648]},
     {loadUnit_maskInput_hi[25647:25632]},
     {loadUnit_maskInput_hi[25631:25616]},
     {loadUnit_maskInput_hi[25615:25600]},
     {loadUnit_maskInput_hi[25599:25584]},
     {loadUnit_maskInput_hi[25583:25568]},
     {loadUnit_maskInput_hi[25567:25552]},
     {loadUnit_maskInput_hi[25551:25536]},
     {loadUnit_maskInput_hi[25535:25520]},
     {loadUnit_maskInput_hi[25519:25504]},
     {loadUnit_maskInput_hi[25503:25488]},
     {loadUnit_maskInput_hi[25487:25472]},
     {loadUnit_maskInput_hi[25471:25456]},
     {loadUnit_maskInput_hi[25455:25440]},
     {loadUnit_maskInput_hi[25439:25424]},
     {loadUnit_maskInput_hi[25423:25408]},
     {loadUnit_maskInput_hi[25407:25392]},
     {loadUnit_maskInput_hi[25391:25376]},
     {loadUnit_maskInput_hi[25375:25360]},
     {loadUnit_maskInput_hi[25359:25344]},
     {loadUnit_maskInput_hi[25343:25328]},
     {loadUnit_maskInput_hi[25327:25312]},
     {loadUnit_maskInput_hi[25311:25296]},
     {loadUnit_maskInput_hi[25295:25280]},
     {loadUnit_maskInput_hi[25279:25264]},
     {loadUnit_maskInput_hi[25263:25248]},
     {loadUnit_maskInput_hi[25247:25232]},
     {loadUnit_maskInput_hi[25231:25216]},
     {loadUnit_maskInput_hi[25215:25200]},
     {loadUnit_maskInput_hi[25199:25184]},
     {loadUnit_maskInput_hi[25183:25168]},
     {loadUnit_maskInput_hi[25167:25152]},
     {loadUnit_maskInput_hi[25151:25136]},
     {loadUnit_maskInput_hi[25135:25120]},
     {loadUnit_maskInput_hi[25119:25104]},
     {loadUnit_maskInput_hi[25103:25088]},
     {loadUnit_maskInput_hi[25087:25072]},
     {loadUnit_maskInput_hi[25071:25056]},
     {loadUnit_maskInput_hi[25055:25040]},
     {loadUnit_maskInput_hi[25039:25024]},
     {loadUnit_maskInput_hi[25023:25008]},
     {loadUnit_maskInput_hi[25007:24992]},
     {loadUnit_maskInput_hi[24991:24976]},
     {loadUnit_maskInput_hi[24975:24960]},
     {loadUnit_maskInput_hi[24959:24944]},
     {loadUnit_maskInput_hi[24943:24928]},
     {loadUnit_maskInput_hi[24927:24912]},
     {loadUnit_maskInput_hi[24911:24896]},
     {loadUnit_maskInput_hi[24895:24880]},
     {loadUnit_maskInput_hi[24879:24864]},
     {loadUnit_maskInput_hi[24863:24848]},
     {loadUnit_maskInput_hi[24847:24832]},
     {loadUnit_maskInput_hi[24831:24816]},
     {loadUnit_maskInput_hi[24815:24800]},
     {loadUnit_maskInput_hi[24799:24784]},
     {loadUnit_maskInput_hi[24783:24768]},
     {loadUnit_maskInput_hi[24767:24752]},
     {loadUnit_maskInput_hi[24751:24736]},
     {loadUnit_maskInput_hi[24735:24720]},
     {loadUnit_maskInput_hi[24719:24704]},
     {loadUnit_maskInput_hi[24703:24688]},
     {loadUnit_maskInput_hi[24687:24672]},
     {loadUnit_maskInput_hi[24671:24656]},
     {loadUnit_maskInput_hi[24655:24640]},
     {loadUnit_maskInput_hi[24639:24624]},
     {loadUnit_maskInput_hi[24623:24608]},
     {loadUnit_maskInput_hi[24607:24592]},
     {loadUnit_maskInput_hi[24591:24576]},
     {loadUnit_maskInput_hi[24575:24560]},
     {loadUnit_maskInput_hi[24559:24544]},
     {loadUnit_maskInput_hi[24543:24528]},
     {loadUnit_maskInput_hi[24527:24512]},
     {loadUnit_maskInput_hi[24511:24496]},
     {loadUnit_maskInput_hi[24495:24480]},
     {loadUnit_maskInput_hi[24479:24464]},
     {loadUnit_maskInput_hi[24463:24448]},
     {loadUnit_maskInput_hi[24447:24432]},
     {loadUnit_maskInput_hi[24431:24416]},
     {loadUnit_maskInput_hi[24415:24400]},
     {loadUnit_maskInput_hi[24399:24384]},
     {loadUnit_maskInput_hi[24383:24368]},
     {loadUnit_maskInput_hi[24367:24352]},
     {loadUnit_maskInput_hi[24351:24336]},
     {loadUnit_maskInput_hi[24335:24320]},
     {loadUnit_maskInput_hi[24319:24304]},
     {loadUnit_maskInput_hi[24303:24288]},
     {loadUnit_maskInput_hi[24287:24272]},
     {loadUnit_maskInput_hi[24271:24256]},
     {loadUnit_maskInput_hi[24255:24240]},
     {loadUnit_maskInput_hi[24239:24224]},
     {loadUnit_maskInput_hi[24223:24208]},
     {loadUnit_maskInput_hi[24207:24192]},
     {loadUnit_maskInput_hi[24191:24176]},
     {loadUnit_maskInput_hi[24175:24160]},
     {loadUnit_maskInput_hi[24159:24144]},
     {loadUnit_maskInput_hi[24143:24128]},
     {loadUnit_maskInput_hi[24127:24112]},
     {loadUnit_maskInput_hi[24111:24096]},
     {loadUnit_maskInput_hi[24095:24080]},
     {loadUnit_maskInput_hi[24079:24064]},
     {loadUnit_maskInput_hi[24063:24048]},
     {loadUnit_maskInput_hi[24047:24032]},
     {loadUnit_maskInput_hi[24031:24016]},
     {loadUnit_maskInput_hi[24015:24000]},
     {loadUnit_maskInput_hi[23999:23984]},
     {loadUnit_maskInput_hi[23983:23968]},
     {loadUnit_maskInput_hi[23967:23952]},
     {loadUnit_maskInput_hi[23951:23936]},
     {loadUnit_maskInput_hi[23935:23920]},
     {loadUnit_maskInput_hi[23919:23904]},
     {loadUnit_maskInput_hi[23903:23888]},
     {loadUnit_maskInput_hi[23887:23872]},
     {loadUnit_maskInput_hi[23871:23856]},
     {loadUnit_maskInput_hi[23855:23840]},
     {loadUnit_maskInput_hi[23839:23824]},
     {loadUnit_maskInput_hi[23823:23808]},
     {loadUnit_maskInput_hi[23807:23792]},
     {loadUnit_maskInput_hi[23791:23776]},
     {loadUnit_maskInput_hi[23775:23760]},
     {loadUnit_maskInput_hi[23759:23744]},
     {loadUnit_maskInput_hi[23743:23728]},
     {loadUnit_maskInput_hi[23727:23712]},
     {loadUnit_maskInput_hi[23711:23696]},
     {loadUnit_maskInput_hi[23695:23680]},
     {loadUnit_maskInput_hi[23679:23664]},
     {loadUnit_maskInput_hi[23663:23648]},
     {loadUnit_maskInput_hi[23647:23632]},
     {loadUnit_maskInput_hi[23631:23616]},
     {loadUnit_maskInput_hi[23615:23600]},
     {loadUnit_maskInput_hi[23599:23584]},
     {loadUnit_maskInput_hi[23583:23568]},
     {loadUnit_maskInput_hi[23567:23552]},
     {loadUnit_maskInput_hi[23551:23536]},
     {loadUnit_maskInput_hi[23535:23520]},
     {loadUnit_maskInput_hi[23519:23504]},
     {loadUnit_maskInput_hi[23503:23488]},
     {loadUnit_maskInput_hi[23487:23472]},
     {loadUnit_maskInput_hi[23471:23456]},
     {loadUnit_maskInput_hi[23455:23440]},
     {loadUnit_maskInput_hi[23439:23424]},
     {loadUnit_maskInput_hi[23423:23408]},
     {loadUnit_maskInput_hi[23407:23392]},
     {loadUnit_maskInput_hi[23391:23376]},
     {loadUnit_maskInput_hi[23375:23360]},
     {loadUnit_maskInput_hi[23359:23344]},
     {loadUnit_maskInput_hi[23343:23328]},
     {loadUnit_maskInput_hi[23327:23312]},
     {loadUnit_maskInput_hi[23311:23296]},
     {loadUnit_maskInput_hi[23295:23280]},
     {loadUnit_maskInput_hi[23279:23264]},
     {loadUnit_maskInput_hi[23263:23248]},
     {loadUnit_maskInput_hi[23247:23232]},
     {loadUnit_maskInput_hi[23231:23216]},
     {loadUnit_maskInput_hi[23215:23200]},
     {loadUnit_maskInput_hi[23199:23184]},
     {loadUnit_maskInput_hi[23183:23168]},
     {loadUnit_maskInput_hi[23167:23152]},
     {loadUnit_maskInput_hi[23151:23136]},
     {loadUnit_maskInput_hi[23135:23120]},
     {loadUnit_maskInput_hi[23119:23104]},
     {loadUnit_maskInput_hi[23103:23088]},
     {loadUnit_maskInput_hi[23087:23072]},
     {loadUnit_maskInput_hi[23071:23056]},
     {loadUnit_maskInput_hi[23055:23040]},
     {loadUnit_maskInput_hi[23039:23024]},
     {loadUnit_maskInput_hi[23023:23008]},
     {loadUnit_maskInput_hi[23007:22992]},
     {loadUnit_maskInput_hi[22991:22976]},
     {loadUnit_maskInput_hi[22975:22960]},
     {loadUnit_maskInput_hi[22959:22944]},
     {loadUnit_maskInput_hi[22943:22928]},
     {loadUnit_maskInput_hi[22927:22912]},
     {loadUnit_maskInput_hi[22911:22896]},
     {loadUnit_maskInput_hi[22895:22880]},
     {loadUnit_maskInput_hi[22879:22864]},
     {loadUnit_maskInput_hi[22863:22848]},
     {loadUnit_maskInput_hi[22847:22832]},
     {loadUnit_maskInput_hi[22831:22816]},
     {loadUnit_maskInput_hi[22815:22800]},
     {loadUnit_maskInput_hi[22799:22784]},
     {loadUnit_maskInput_hi[22783:22768]},
     {loadUnit_maskInput_hi[22767:22752]},
     {loadUnit_maskInput_hi[22751:22736]},
     {loadUnit_maskInput_hi[22735:22720]},
     {loadUnit_maskInput_hi[22719:22704]},
     {loadUnit_maskInput_hi[22703:22688]},
     {loadUnit_maskInput_hi[22687:22672]},
     {loadUnit_maskInput_hi[22671:22656]},
     {loadUnit_maskInput_hi[22655:22640]},
     {loadUnit_maskInput_hi[22639:22624]},
     {loadUnit_maskInput_hi[22623:22608]},
     {loadUnit_maskInput_hi[22607:22592]},
     {loadUnit_maskInput_hi[22591:22576]},
     {loadUnit_maskInput_hi[22575:22560]},
     {loadUnit_maskInput_hi[22559:22544]},
     {loadUnit_maskInput_hi[22543:22528]},
     {loadUnit_maskInput_hi[22527:22512]},
     {loadUnit_maskInput_hi[22511:22496]},
     {loadUnit_maskInput_hi[22495:22480]},
     {loadUnit_maskInput_hi[22479:22464]},
     {loadUnit_maskInput_hi[22463:22448]},
     {loadUnit_maskInput_hi[22447:22432]},
     {loadUnit_maskInput_hi[22431:22416]},
     {loadUnit_maskInput_hi[22415:22400]},
     {loadUnit_maskInput_hi[22399:22384]},
     {loadUnit_maskInput_hi[22383:22368]},
     {loadUnit_maskInput_hi[22367:22352]},
     {loadUnit_maskInput_hi[22351:22336]},
     {loadUnit_maskInput_hi[22335:22320]},
     {loadUnit_maskInput_hi[22319:22304]},
     {loadUnit_maskInput_hi[22303:22288]},
     {loadUnit_maskInput_hi[22287:22272]},
     {loadUnit_maskInput_hi[22271:22256]},
     {loadUnit_maskInput_hi[22255:22240]},
     {loadUnit_maskInput_hi[22239:22224]},
     {loadUnit_maskInput_hi[22223:22208]},
     {loadUnit_maskInput_hi[22207:22192]},
     {loadUnit_maskInput_hi[22191:22176]},
     {loadUnit_maskInput_hi[22175:22160]},
     {loadUnit_maskInput_hi[22159:22144]},
     {loadUnit_maskInput_hi[22143:22128]},
     {loadUnit_maskInput_hi[22127:22112]},
     {loadUnit_maskInput_hi[22111:22096]},
     {loadUnit_maskInput_hi[22095:22080]},
     {loadUnit_maskInput_hi[22079:22064]},
     {loadUnit_maskInput_hi[22063:22048]},
     {loadUnit_maskInput_hi[22047:22032]},
     {loadUnit_maskInput_hi[22031:22016]},
     {loadUnit_maskInput_hi[22015:22000]},
     {loadUnit_maskInput_hi[21999:21984]},
     {loadUnit_maskInput_hi[21983:21968]},
     {loadUnit_maskInput_hi[21967:21952]},
     {loadUnit_maskInput_hi[21951:21936]},
     {loadUnit_maskInput_hi[21935:21920]},
     {loadUnit_maskInput_hi[21919:21904]},
     {loadUnit_maskInput_hi[21903:21888]},
     {loadUnit_maskInput_hi[21887:21872]},
     {loadUnit_maskInput_hi[21871:21856]},
     {loadUnit_maskInput_hi[21855:21840]},
     {loadUnit_maskInput_hi[21839:21824]},
     {loadUnit_maskInput_hi[21823:21808]},
     {loadUnit_maskInput_hi[21807:21792]},
     {loadUnit_maskInput_hi[21791:21776]},
     {loadUnit_maskInput_hi[21775:21760]},
     {loadUnit_maskInput_hi[21759:21744]},
     {loadUnit_maskInput_hi[21743:21728]},
     {loadUnit_maskInput_hi[21727:21712]},
     {loadUnit_maskInput_hi[21711:21696]},
     {loadUnit_maskInput_hi[21695:21680]},
     {loadUnit_maskInput_hi[21679:21664]},
     {loadUnit_maskInput_hi[21663:21648]},
     {loadUnit_maskInput_hi[21647:21632]},
     {loadUnit_maskInput_hi[21631:21616]},
     {loadUnit_maskInput_hi[21615:21600]},
     {loadUnit_maskInput_hi[21599:21584]},
     {loadUnit_maskInput_hi[21583:21568]},
     {loadUnit_maskInput_hi[21567:21552]},
     {loadUnit_maskInput_hi[21551:21536]},
     {loadUnit_maskInput_hi[21535:21520]},
     {loadUnit_maskInput_hi[21519:21504]},
     {loadUnit_maskInput_hi[21503:21488]},
     {loadUnit_maskInput_hi[21487:21472]},
     {loadUnit_maskInput_hi[21471:21456]},
     {loadUnit_maskInput_hi[21455:21440]},
     {loadUnit_maskInput_hi[21439:21424]},
     {loadUnit_maskInput_hi[21423:21408]},
     {loadUnit_maskInput_hi[21407:21392]},
     {loadUnit_maskInput_hi[21391:21376]},
     {loadUnit_maskInput_hi[21375:21360]},
     {loadUnit_maskInput_hi[21359:21344]},
     {loadUnit_maskInput_hi[21343:21328]},
     {loadUnit_maskInput_hi[21327:21312]},
     {loadUnit_maskInput_hi[21311:21296]},
     {loadUnit_maskInput_hi[21295:21280]},
     {loadUnit_maskInput_hi[21279:21264]},
     {loadUnit_maskInput_hi[21263:21248]},
     {loadUnit_maskInput_hi[21247:21232]},
     {loadUnit_maskInput_hi[21231:21216]},
     {loadUnit_maskInput_hi[21215:21200]},
     {loadUnit_maskInput_hi[21199:21184]},
     {loadUnit_maskInput_hi[21183:21168]},
     {loadUnit_maskInput_hi[21167:21152]},
     {loadUnit_maskInput_hi[21151:21136]},
     {loadUnit_maskInput_hi[21135:21120]},
     {loadUnit_maskInput_hi[21119:21104]},
     {loadUnit_maskInput_hi[21103:21088]},
     {loadUnit_maskInput_hi[21087:21072]},
     {loadUnit_maskInput_hi[21071:21056]},
     {loadUnit_maskInput_hi[21055:21040]},
     {loadUnit_maskInput_hi[21039:21024]},
     {loadUnit_maskInput_hi[21023:21008]},
     {loadUnit_maskInput_hi[21007:20992]},
     {loadUnit_maskInput_hi[20991:20976]},
     {loadUnit_maskInput_hi[20975:20960]},
     {loadUnit_maskInput_hi[20959:20944]},
     {loadUnit_maskInput_hi[20943:20928]},
     {loadUnit_maskInput_hi[20927:20912]},
     {loadUnit_maskInput_hi[20911:20896]},
     {loadUnit_maskInput_hi[20895:20880]},
     {loadUnit_maskInput_hi[20879:20864]},
     {loadUnit_maskInput_hi[20863:20848]},
     {loadUnit_maskInput_hi[20847:20832]},
     {loadUnit_maskInput_hi[20831:20816]},
     {loadUnit_maskInput_hi[20815:20800]},
     {loadUnit_maskInput_hi[20799:20784]},
     {loadUnit_maskInput_hi[20783:20768]},
     {loadUnit_maskInput_hi[20767:20752]},
     {loadUnit_maskInput_hi[20751:20736]},
     {loadUnit_maskInput_hi[20735:20720]},
     {loadUnit_maskInput_hi[20719:20704]},
     {loadUnit_maskInput_hi[20703:20688]},
     {loadUnit_maskInput_hi[20687:20672]},
     {loadUnit_maskInput_hi[20671:20656]},
     {loadUnit_maskInput_hi[20655:20640]},
     {loadUnit_maskInput_hi[20639:20624]},
     {loadUnit_maskInput_hi[20623:20608]},
     {loadUnit_maskInput_hi[20607:20592]},
     {loadUnit_maskInput_hi[20591:20576]},
     {loadUnit_maskInput_hi[20575:20560]},
     {loadUnit_maskInput_hi[20559:20544]},
     {loadUnit_maskInput_hi[20543:20528]},
     {loadUnit_maskInput_hi[20527:20512]},
     {loadUnit_maskInput_hi[20511:20496]},
     {loadUnit_maskInput_hi[20495:20480]},
     {loadUnit_maskInput_hi[20479:20464]},
     {loadUnit_maskInput_hi[20463:20448]},
     {loadUnit_maskInput_hi[20447:20432]},
     {loadUnit_maskInput_hi[20431:20416]},
     {loadUnit_maskInput_hi[20415:20400]},
     {loadUnit_maskInput_hi[20399:20384]},
     {loadUnit_maskInput_hi[20383:20368]},
     {loadUnit_maskInput_hi[20367:20352]},
     {loadUnit_maskInput_hi[20351:20336]},
     {loadUnit_maskInput_hi[20335:20320]},
     {loadUnit_maskInput_hi[20319:20304]},
     {loadUnit_maskInput_hi[20303:20288]},
     {loadUnit_maskInput_hi[20287:20272]},
     {loadUnit_maskInput_hi[20271:20256]},
     {loadUnit_maskInput_hi[20255:20240]},
     {loadUnit_maskInput_hi[20239:20224]},
     {loadUnit_maskInput_hi[20223:20208]},
     {loadUnit_maskInput_hi[20207:20192]},
     {loadUnit_maskInput_hi[20191:20176]},
     {loadUnit_maskInput_hi[20175:20160]},
     {loadUnit_maskInput_hi[20159:20144]},
     {loadUnit_maskInput_hi[20143:20128]},
     {loadUnit_maskInput_hi[20127:20112]},
     {loadUnit_maskInput_hi[20111:20096]},
     {loadUnit_maskInput_hi[20095:20080]},
     {loadUnit_maskInput_hi[20079:20064]},
     {loadUnit_maskInput_hi[20063:20048]},
     {loadUnit_maskInput_hi[20047:20032]},
     {loadUnit_maskInput_hi[20031:20016]},
     {loadUnit_maskInput_hi[20015:20000]},
     {loadUnit_maskInput_hi[19999:19984]},
     {loadUnit_maskInput_hi[19983:19968]},
     {loadUnit_maskInput_hi[19967:19952]},
     {loadUnit_maskInput_hi[19951:19936]},
     {loadUnit_maskInput_hi[19935:19920]},
     {loadUnit_maskInput_hi[19919:19904]},
     {loadUnit_maskInput_hi[19903:19888]},
     {loadUnit_maskInput_hi[19887:19872]},
     {loadUnit_maskInput_hi[19871:19856]},
     {loadUnit_maskInput_hi[19855:19840]},
     {loadUnit_maskInput_hi[19839:19824]},
     {loadUnit_maskInput_hi[19823:19808]},
     {loadUnit_maskInput_hi[19807:19792]},
     {loadUnit_maskInput_hi[19791:19776]},
     {loadUnit_maskInput_hi[19775:19760]},
     {loadUnit_maskInput_hi[19759:19744]},
     {loadUnit_maskInput_hi[19743:19728]},
     {loadUnit_maskInput_hi[19727:19712]},
     {loadUnit_maskInput_hi[19711:19696]},
     {loadUnit_maskInput_hi[19695:19680]},
     {loadUnit_maskInput_hi[19679:19664]},
     {loadUnit_maskInput_hi[19663:19648]},
     {loadUnit_maskInput_hi[19647:19632]},
     {loadUnit_maskInput_hi[19631:19616]},
     {loadUnit_maskInput_hi[19615:19600]},
     {loadUnit_maskInput_hi[19599:19584]},
     {loadUnit_maskInput_hi[19583:19568]},
     {loadUnit_maskInput_hi[19567:19552]},
     {loadUnit_maskInput_hi[19551:19536]},
     {loadUnit_maskInput_hi[19535:19520]},
     {loadUnit_maskInput_hi[19519:19504]},
     {loadUnit_maskInput_hi[19503:19488]},
     {loadUnit_maskInput_hi[19487:19472]},
     {loadUnit_maskInput_hi[19471:19456]},
     {loadUnit_maskInput_hi[19455:19440]},
     {loadUnit_maskInput_hi[19439:19424]},
     {loadUnit_maskInput_hi[19423:19408]},
     {loadUnit_maskInput_hi[19407:19392]},
     {loadUnit_maskInput_hi[19391:19376]},
     {loadUnit_maskInput_hi[19375:19360]},
     {loadUnit_maskInput_hi[19359:19344]},
     {loadUnit_maskInput_hi[19343:19328]},
     {loadUnit_maskInput_hi[19327:19312]},
     {loadUnit_maskInput_hi[19311:19296]},
     {loadUnit_maskInput_hi[19295:19280]},
     {loadUnit_maskInput_hi[19279:19264]},
     {loadUnit_maskInput_hi[19263:19248]},
     {loadUnit_maskInput_hi[19247:19232]},
     {loadUnit_maskInput_hi[19231:19216]},
     {loadUnit_maskInput_hi[19215:19200]},
     {loadUnit_maskInput_hi[19199:19184]},
     {loadUnit_maskInput_hi[19183:19168]},
     {loadUnit_maskInput_hi[19167:19152]},
     {loadUnit_maskInput_hi[19151:19136]},
     {loadUnit_maskInput_hi[19135:19120]},
     {loadUnit_maskInput_hi[19119:19104]},
     {loadUnit_maskInput_hi[19103:19088]},
     {loadUnit_maskInput_hi[19087:19072]},
     {loadUnit_maskInput_hi[19071:19056]},
     {loadUnit_maskInput_hi[19055:19040]},
     {loadUnit_maskInput_hi[19039:19024]},
     {loadUnit_maskInput_hi[19023:19008]},
     {loadUnit_maskInput_hi[19007:18992]},
     {loadUnit_maskInput_hi[18991:18976]},
     {loadUnit_maskInput_hi[18975:18960]},
     {loadUnit_maskInput_hi[18959:18944]},
     {loadUnit_maskInput_hi[18943:18928]},
     {loadUnit_maskInput_hi[18927:18912]},
     {loadUnit_maskInput_hi[18911:18896]},
     {loadUnit_maskInput_hi[18895:18880]},
     {loadUnit_maskInput_hi[18879:18864]},
     {loadUnit_maskInput_hi[18863:18848]},
     {loadUnit_maskInput_hi[18847:18832]},
     {loadUnit_maskInput_hi[18831:18816]},
     {loadUnit_maskInput_hi[18815:18800]},
     {loadUnit_maskInput_hi[18799:18784]},
     {loadUnit_maskInput_hi[18783:18768]},
     {loadUnit_maskInput_hi[18767:18752]},
     {loadUnit_maskInput_hi[18751:18736]},
     {loadUnit_maskInput_hi[18735:18720]},
     {loadUnit_maskInput_hi[18719:18704]},
     {loadUnit_maskInput_hi[18703:18688]},
     {loadUnit_maskInput_hi[18687:18672]},
     {loadUnit_maskInput_hi[18671:18656]},
     {loadUnit_maskInput_hi[18655:18640]},
     {loadUnit_maskInput_hi[18639:18624]},
     {loadUnit_maskInput_hi[18623:18608]},
     {loadUnit_maskInput_hi[18607:18592]},
     {loadUnit_maskInput_hi[18591:18576]},
     {loadUnit_maskInput_hi[18575:18560]},
     {loadUnit_maskInput_hi[18559:18544]},
     {loadUnit_maskInput_hi[18543:18528]},
     {loadUnit_maskInput_hi[18527:18512]},
     {loadUnit_maskInput_hi[18511:18496]},
     {loadUnit_maskInput_hi[18495:18480]},
     {loadUnit_maskInput_hi[18479:18464]},
     {loadUnit_maskInput_hi[18463:18448]},
     {loadUnit_maskInput_hi[18447:18432]},
     {loadUnit_maskInput_hi[18431:18416]},
     {loadUnit_maskInput_hi[18415:18400]},
     {loadUnit_maskInput_hi[18399:18384]},
     {loadUnit_maskInput_hi[18383:18368]},
     {loadUnit_maskInput_hi[18367:18352]},
     {loadUnit_maskInput_hi[18351:18336]},
     {loadUnit_maskInput_hi[18335:18320]},
     {loadUnit_maskInput_hi[18319:18304]},
     {loadUnit_maskInput_hi[18303:18288]},
     {loadUnit_maskInput_hi[18287:18272]},
     {loadUnit_maskInput_hi[18271:18256]},
     {loadUnit_maskInput_hi[18255:18240]},
     {loadUnit_maskInput_hi[18239:18224]},
     {loadUnit_maskInput_hi[18223:18208]},
     {loadUnit_maskInput_hi[18207:18192]},
     {loadUnit_maskInput_hi[18191:18176]},
     {loadUnit_maskInput_hi[18175:18160]},
     {loadUnit_maskInput_hi[18159:18144]},
     {loadUnit_maskInput_hi[18143:18128]},
     {loadUnit_maskInput_hi[18127:18112]},
     {loadUnit_maskInput_hi[18111:18096]},
     {loadUnit_maskInput_hi[18095:18080]},
     {loadUnit_maskInput_hi[18079:18064]},
     {loadUnit_maskInput_hi[18063:18048]},
     {loadUnit_maskInput_hi[18047:18032]},
     {loadUnit_maskInput_hi[18031:18016]},
     {loadUnit_maskInput_hi[18015:18000]},
     {loadUnit_maskInput_hi[17999:17984]},
     {loadUnit_maskInput_hi[17983:17968]},
     {loadUnit_maskInput_hi[17967:17952]},
     {loadUnit_maskInput_hi[17951:17936]},
     {loadUnit_maskInput_hi[17935:17920]},
     {loadUnit_maskInput_hi[17919:17904]},
     {loadUnit_maskInput_hi[17903:17888]},
     {loadUnit_maskInput_hi[17887:17872]},
     {loadUnit_maskInput_hi[17871:17856]},
     {loadUnit_maskInput_hi[17855:17840]},
     {loadUnit_maskInput_hi[17839:17824]},
     {loadUnit_maskInput_hi[17823:17808]},
     {loadUnit_maskInput_hi[17807:17792]},
     {loadUnit_maskInput_hi[17791:17776]},
     {loadUnit_maskInput_hi[17775:17760]},
     {loadUnit_maskInput_hi[17759:17744]},
     {loadUnit_maskInput_hi[17743:17728]},
     {loadUnit_maskInput_hi[17727:17712]},
     {loadUnit_maskInput_hi[17711:17696]},
     {loadUnit_maskInput_hi[17695:17680]},
     {loadUnit_maskInput_hi[17679:17664]},
     {loadUnit_maskInput_hi[17663:17648]},
     {loadUnit_maskInput_hi[17647:17632]},
     {loadUnit_maskInput_hi[17631:17616]},
     {loadUnit_maskInput_hi[17615:17600]},
     {loadUnit_maskInput_hi[17599:17584]},
     {loadUnit_maskInput_hi[17583:17568]},
     {loadUnit_maskInput_hi[17567:17552]},
     {loadUnit_maskInput_hi[17551:17536]},
     {loadUnit_maskInput_hi[17535:17520]},
     {loadUnit_maskInput_hi[17519:17504]},
     {loadUnit_maskInput_hi[17503:17488]},
     {loadUnit_maskInput_hi[17487:17472]},
     {loadUnit_maskInput_hi[17471:17456]},
     {loadUnit_maskInput_hi[17455:17440]},
     {loadUnit_maskInput_hi[17439:17424]},
     {loadUnit_maskInput_hi[17423:17408]},
     {loadUnit_maskInput_hi[17407:17392]},
     {loadUnit_maskInput_hi[17391:17376]},
     {loadUnit_maskInput_hi[17375:17360]},
     {loadUnit_maskInput_hi[17359:17344]},
     {loadUnit_maskInput_hi[17343:17328]},
     {loadUnit_maskInput_hi[17327:17312]},
     {loadUnit_maskInput_hi[17311:17296]},
     {loadUnit_maskInput_hi[17295:17280]},
     {loadUnit_maskInput_hi[17279:17264]},
     {loadUnit_maskInput_hi[17263:17248]},
     {loadUnit_maskInput_hi[17247:17232]},
     {loadUnit_maskInput_hi[17231:17216]},
     {loadUnit_maskInput_hi[17215:17200]},
     {loadUnit_maskInput_hi[17199:17184]},
     {loadUnit_maskInput_hi[17183:17168]},
     {loadUnit_maskInput_hi[17167:17152]},
     {loadUnit_maskInput_hi[17151:17136]},
     {loadUnit_maskInput_hi[17135:17120]},
     {loadUnit_maskInput_hi[17119:17104]},
     {loadUnit_maskInput_hi[17103:17088]},
     {loadUnit_maskInput_hi[17087:17072]},
     {loadUnit_maskInput_hi[17071:17056]},
     {loadUnit_maskInput_hi[17055:17040]},
     {loadUnit_maskInput_hi[17039:17024]},
     {loadUnit_maskInput_hi[17023:17008]},
     {loadUnit_maskInput_hi[17007:16992]},
     {loadUnit_maskInput_hi[16991:16976]},
     {loadUnit_maskInput_hi[16975:16960]},
     {loadUnit_maskInput_hi[16959:16944]},
     {loadUnit_maskInput_hi[16943:16928]},
     {loadUnit_maskInput_hi[16927:16912]},
     {loadUnit_maskInput_hi[16911:16896]},
     {loadUnit_maskInput_hi[16895:16880]},
     {loadUnit_maskInput_hi[16879:16864]},
     {loadUnit_maskInput_hi[16863:16848]},
     {loadUnit_maskInput_hi[16847:16832]},
     {loadUnit_maskInput_hi[16831:16816]},
     {loadUnit_maskInput_hi[16815:16800]},
     {loadUnit_maskInput_hi[16799:16784]},
     {loadUnit_maskInput_hi[16783:16768]},
     {loadUnit_maskInput_hi[16767:16752]},
     {loadUnit_maskInput_hi[16751:16736]},
     {loadUnit_maskInput_hi[16735:16720]},
     {loadUnit_maskInput_hi[16719:16704]},
     {loadUnit_maskInput_hi[16703:16688]},
     {loadUnit_maskInput_hi[16687:16672]},
     {loadUnit_maskInput_hi[16671:16656]},
     {loadUnit_maskInput_hi[16655:16640]},
     {loadUnit_maskInput_hi[16639:16624]},
     {loadUnit_maskInput_hi[16623:16608]},
     {loadUnit_maskInput_hi[16607:16592]},
     {loadUnit_maskInput_hi[16591:16576]},
     {loadUnit_maskInput_hi[16575:16560]},
     {loadUnit_maskInput_hi[16559:16544]},
     {loadUnit_maskInput_hi[16543:16528]},
     {loadUnit_maskInput_hi[16527:16512]},
     {loadUnit_maskInput_hi[16511:16496]},
     {loadUnit_maskInput_hi[16495:16480]},
     {loadUnit_maskInput_hi[16479:16464]},
     {loadUnit_maskInput_hi[16463:16448]},
     {loadUnit_maskInput_hi[16447:16432]},
     {loadUnit_maskInput_hi[16431:16416]},
     {loadUnit_maskInput_hi[16415:16400]},
     {loadUnit_maskInput_hi[16399:16384]},
     {loadUnit_maskInput_hi[16383:16368]},
     {loadUnit_maskInput_hi[16367:16352]},
     {loadUnit_maskInput_hi[16351:16336]},
     {loadUnit_maskInput_hi[16335:16320]},
     {loadUnit_maskInput_hi[16319:16304]},
     {loadUnit_maskInput_hi[16303:16288]},
     {loadUnit_maskInput_hi[16287:16272]},
     {loadUnit_maskInput_hi[16271:16256]},
     {loadUnit_maskInput_hi[16255:16240]},
     {loadUnit_maskInput_hi[16239:16224]},
     {loadUnit_maskInput_hi[16223:16208]},
     {loadUnit_maskInput_hi[16207:16192]},
     {loadUnit_maskInput_hi[16191:16176]},
     {loadUnit_maskInput_hi[16175:16160]},
     {loadUnit_maskInput_hi[16159:16144]},
     {loadUnit_maskInput_hi[16143:16128]},
     {loadUnit_maskInput_hi[16127:16112]},
     {loadUnit_maskInput_hi[16111:16096]},
     {loadUnit_maskInput_hi[16095:16080]},
     {loadUnit_maskInput_hi[16079:16064]},
     {loadUnit_maskInput_hi[16063:16048]},
     {loadUnit_maskInput_hi[16047:16032]},
     {loadUnit_maskInput_hi[16031:16016]},
     {loadUnit_maskInput_hi[16015:16000]},
     {loadUnit_maskInput_hi[15999:15984]},
     {loadUnit_maskInput_hi[15983:15968]},
     {loadUnit_maskInput_hi[15967:15952]},
     {loadUnit_maskInput_hi[15951:15936]},
     {loadUnit_maskInput_hi[15935:15920]},
     {loadUnit_maskInput_hi[15919:15904]},
     {loadUnit_maskInput_hi[15903:15888]},
     {loadUnit_maskInput_hi[15887:15872]},
     {loadUnit_maskInput_hi[15871:15856]},
     {loadUnit_maskInput_hi[15855:15840]},
     {loadUnit_maskInput_hi[15839:15824]},
     {loadUnit_maskInput_hi[15823:15808]},
     {loadUnit_maskInput_hi[15807:15792]},
     {loadUnit_maskInput_hi[15791:15776]},
     {loadUnit_maskInput_hi[15775:15760]},
     {loadUnit_maskInput_hi[15759:15744]},
     {loadUnit_maskInput_hi[15743:15728]},
     {loadUnit_maskInput_hi[15727:15712]},
     {loadUnit_maskInput_hi[15711:15696]},
     {loadUnit_maskInput_hi[15695:15680]},
     {loadUnit_maskInput_hi[15679:15664]},
     {loadUnit_maskInput_hi[15663:15648]},
     {loadUnit_maskInput_hi[15647:15632]},
     {loadUnit_maskInput_hi[15631:15616]},
     {loadUnit_maskInput_hi[15615:15600]},
     {loadUnit_maskInput_hi[15599:15584]},
     {loadUnit_maskInput_hi[15583:15568]},
     {loadUnit_maskInput_hi[15567:15552]},
     {loadUnit_maskInput_hi[15551:15536]},
     {loadUnit_maskInput_hi[15535:15520]},
     {loadUnit_maskInput_hi[15519:15504]},
     {loadUnit_maskInput_hi[15503:15488]},
     {loadUnit_maskInput_hi[15487:15472]},
     {loadUnit_maskInput_hi[15471:15456]},
     {loadUnit_maskInput_hi[15455:15440]},
     {loadUnit_maskInput_hi[15439:15424]},
     {loadUnit_maskInput_hi[15423:15408]},
     {loadUnit_maskInput_hi[15407:15392]},
     {loadUnit_maskInput_hi[15391:15376]},
     {loadUnit_maskInput_hi[15375:15360]},
     {loadUnit_maskInput_hi[15359:15344]},
     {loadUnit_maskInput_hi[15343:15328]},
     {loadUnit_maskInput_hi[15327:15312]},
     {loadUnit_maskInput_hi[15311:15296]},
     {loadUnit_maskInput_hi[15295:15280]},
     {loadUnit_maskInput_hi[15279:15264]},
     {loadUnit_maskInput_hi[15263:15248]},
     {loadUnit_maskInput_hi[15247:15232]},
     {loadUnit_maskInput_hi[15231:15216]},
     {loadUnit_maskInput_hi[15215:15200]},
     {loadUnit_maskInput_hi[15199:15184]},
     {loadUnit_maskInput_hi[15183:15168]},
     {loadUnit_maskInput_hi[15167:15152]},
     {loadUnit_maskInput_hi[15151:15136]},
     {loadUnit_maskInput_hi[15135:15120]},
     {loadUnit_maskInput_hi[15119:15104]},
     {loadUnit_maskInput_hi[15103:15088]},
     {loadUnit_maskInput_hi[15087:15072]},
     {loadUnit_maskInput_hi[15071:15056]},
     {loadUnit_maskInput_hi[15055:15040]},
     {loadUnit_maskInput_hi[15039:15024]},
     {loadUnit_maskInput_hi[15023:15008]},
     {loadUnit_maskInput_hi[15007:14992]},
     {loadUnit_maskInput_hi[14991:14976]},
     {loadUnit_maskInput_hi[14975:14960]},
     {loadUnit_maskInput_hi[14959:14944]},
     {loadUnit_maskInput_hi[14943:14928]},
     {loadUnit_maskInput_hi[14927:14912]},
     {loadUnit_maskInput_hi[14911:14896]},
     {loadUnit_maskInput_hi[14895:14880]},
     {loadUnit_maskInput_hi[14879:14864]},
     {loadUnit_maskInput_hi[14863:14848]},
     {loadUnit_maskInput_hi[14847:14832]},
     {loadUnit_maskInput_hi[14831:14816]},
     {loadUnit_maskInput_hi[14815:14800]},
     {loadUnit_maskInput_hi[14799:14784]},
     {loadUnit_maskInput_hi[14783:14768]},
     {loadUnit_maskInput_hi[14767:14752]},
     {loadUnit_maskInput_hi[14751:14736]},
     {loadUnit_maskInput_hi[14735:14720]},
     {loadUnit_maskInput_hi[14719:14704]},
     {loadUnit_maskInput_hi[14703:14688]},
     {loadUnit_maskInput_hi[14687:14672]},
     {loadUnit_maskInput_hi[14671:14656]},
     {loadUnit_maskInput_hi[14655:14640]},
     {loadUnit_maskInput_hi[14639:14624]},
     {loadUnit_maskInput_hi[14623:14608]},
     {loadUnit_maskInput_hi[14607:14592]},
     {loadUnit_maskInput_hi[14591:14576]},
     {loadUnit_maskInput_hi[14575:14560]},
     {loadUnit_maskInput_hi[14559:14544]},
     {loadUnit_maskInput_hi[14543:14528]},
     {loadUnit_maskInput_hi[14527:14512]},
     {loadUnit_maskInput_hi[14511:14496]},
     {loadUnit_maskInput_hi[14495:14480]},
     {loadUnit_maskInput_hi[14479:14464]},
     {loadUnit_maskInput_hi[14463:14448]},
     {loadUnit_maskInput_hi[14447:14432]},
     {loadUnit_maskInput_hi[14431:14416]},
     {loadUnit_maskInput_hi[14415:14400]},
     {loadUnit_maskInput_hi[14399:14384]},
     {loadUnit_maskInput_hi[14383:14368]},
     {loadUnit_maskInput_hi[14367:14352]},
     {loadUnit_maskInput_hi[14351:14336]},
     {loadUnit_maskInput_hi[14335:14320]},
     {loadUnit_maskInput_hi[14319:14304]},
     {loadUnit_maskInput_hi[14303:14288]},
     {loadUnit_maskInput_hi[14287:14272]},
     {loadUnit_maskInput_hi[14271:14256]},
     {loadUnit_maskInput_hi[14255:14240]},
     {loadUnit_maskInput_hi[14239:14224]},
     {loadUnit_maskInput_hi[14223:14208]},
     {loadUnit_maskInput_hi[14207:14192]},
     {loadUnit_maskInput_hi[14191:14176]},
     {loadUnit_maskInput_hi[14175:14160]},
     {loadUnit_maskInput_hi[14159:14144]},
     {loadUnit_maskInput_hi[14143:14128]},
     {loadUnit_maskInput_hi[14127:14112]},
     {loadUnit_maskInput_hi[14111:14096]},
     {loadUnit_maskInput_hi[14095:14080]},
     {loadUnit_maskInput_hi[14079:14064]},
     {loadUnit_maskInput_hi[14063:14048]},
     {loadUnit_maskInput_hi[14047:14032]},
     {loadUnit_maskInput_hi[14031:14016]},
     {loadUnit_maskInput_hi[14015:14000]},
     {loadUnit_maskInput_hi[13999:13984]},
     {loadUnit_maskInput_hi[13983:13968]},
     {loadUnit_maskInput_hi[13967:13952]},
     {loadUnit_maskInput_hi[13951:13936]},
     {loadUnit_maskInput_hi[13935:13920]},
     {loadUnit_maskInput_hi[13919:13904]},
     {loadUnit_maskInput_hi[13903:13888]},
     {loadUnit_maskInput_hi[13887:13872]},
     {loadUnit_maskInput_hi[13871:13856]},
     {loadUnit_maskInput_hi[13855:13840]},
     {loadUnit_maskInput_hi[13839:13824]},
     {loadUnit_maskInput_hi[13823:13808]},
     {loadUnit_maskInput_hi[13807:13792]},
     {loadUnit_maskInput_hi[13791:13776]},
     {loadUnit_maskInput_hi[13775:13760]},
     {loadUnit_maskInput_hi[13759:13744]},
     {loadUnit_maskInput_hi[13743:13728]},
     {loadUnit_maskInput_hi[13727:13712]},
     {loadUnit_maskInput_hi[13711:13696]},
     {loadUnit_maskInput_hi[13695:13680]},
     {loadUnit_maskInput_hi[13679:13664]},
     {loadUnit_maskInput_hi[13663:13648]},
     {loadUnit_maskInput_hi[13647:13632]},
     {loadUnit_maskInput_hi[13631:13616]},
     {loadUnit_maskInput_hi[13615:13600]},
     {loadUnit_maskInput_hi[13599:13584]},
     {loadUnit_maskInput_hi[13583:13568]},
     {loadUnit_maskInput_hi[13567:13552]},
     {loadUnit_maskInput_hi[13551:13536]},
     {loadUnit_maskInput_hi[13535:13520]},
     {loadUnit_maskInput_hi[13519:13504]},
     {loadUnit_maskInput_hi[13503:13488]},
     {loadUnit_maskInput_hi[13487:13472]},
     {loadUnit_maskInput_hi[13471:13456]},
     {loadUnit_maskInput_hi[13455:13440]},
     {loadUnit_maskInput_hi[13439:13424]},
     {loadUnit_maskInput_hi[13423:13408]},
     {loadUnit_maskInput_hi[13407:13392]},
     {loadUnit_maskInput_hi[13391:13376]},
     {loadUnit_maskInput_hi[13375:13360]},
     {loadUnit_maskInput_hi[13359:13344]},
     {loadUnit_maskInput_hi[13343:13328]},
     {loadUnit_maskInput_hi[13327:13312]},
     {loadUnit_maskInput_hi[13311:13296]},
     {loadUnit_maskInput_hi[13295:13280]},
     {loadUnit_maskInput_hi[13279:13264]},
     {loadUnit_maskInput_hi[13263:13248]},
     {loadUnit_maskInput_hi[13247:13232]},
     {loadUnit_maskInput_hi[13231:13216]},
     {loadUnit_maskInput_hi[13215:13200]},
     {loadUnit_maskInput_hi[13199:13184]},
     {loadUnit_maskInput_hi[13183:13168]},
     {loadUnit_maskInput_hi[13167:13152]},
     {loadUnit_maskInput_hi[13151:13136]},
     {loadUnit_maskInput_hi[13135:13120]},
     {loadUnit_maskInput_hi[13119:13104]},
     {loadUnit_maskInput_hi[13103:13088]},
     {loadUnit_maskInput_hi[13087:13072]},
     {loadUnit_maskInput_hi[13071:13056]},
     {loadUnit_maskInput_hi[13055:13040]},
     {loadUnit_maskInput_hi[13039:13024]},
     {loadUnit_maskInput_hi[13023:13008]},
     {loadUnit_maskInput_hi[13007:12992]},
     {loadUnit_maskInput_hi[12991:12976]},
     {loadUnit_maskInput_hi[12975:12960]},
     {loadUnit_maskInput_hi[12959:12944]},
     {loadUnit_maskInput_hi[12943:12928]},
     {loadUnit_maskInput_hi[12927:12912]},
     {loadUnit_maskInput_hi[12911:12896]},
     {loadUnit_maskInput_hi[12895:12880]},
     {loadUnit_maskInput_hi[12879:12864]},
     {loadUnit_maskInput_hi[12863:12848]},
     {loadUnit_maskInput_hi[12847:12832]},
     {loadUnit_maskInput_hi[12831:12816]},
     {loadUnit_maskInput_hi[12815:12800]},
     {loadUnit_maskInput_hi[12799:12784]},
     {loadUnit_maskInput_hi[12783:12768]},
     {loadUnit_maskInput_hi[12767:12752]},
     {loadUnit_maskInput_hi[12751:12736]},
     {loadUnit_maskInput_hi[12735:12720]},
     {loadUnit_maskInput_hi[12719:12704]},
     {loadUnit_maskInput_hi[12703:12688]},
     {loadUnit_maskInput_hi[12687:12672]},
     {loadUnit_maskInput_hi[12671:12656]},
     {loadUnit_maskInput_hi[12655:12640]},
     {loadUnit_maskInput_hi[12639:12624]},
     {loadUnit_maskInput_hi[12623:12608]},
     {loadUnit_maskInput_hi[12607:12592]},
     {loadUnit_maskInput_hi[12591:12576]},
     {loadUnit_maskInput_hi[12575:12560]},
     {loadUnit_maskInput_hi[12559:12544]},
     {loadUnit_maskInput_hi[12543:12528]},
     {loadUnit_maskInput_hi[12527:12512]},
     {loadUnit_maskInput_hi[12511:12496]},
     {loadUnit_maskInput_hi[12495:12480]},
     {loadUnit_maskInput_hi[12479:12464]},
     {loadUnit_maskInput_hi[12463:12448]},
     {loadUnit_maskInput_hi[12447:12432]},
     {loadUnit_maskInput_hi[12431:12416]},
     {loadUnit_maskInput_hi[12415:12400]},
     {loadUnit_maskInput_hi[12399:12384]},
     {loadUnit_maskInput_hi[12383:12368]},
     {loadUnit_maskInput_hi[12367:12352]},
     {loadUnit_maskInput_hi[12351:12336]},
     {loadUnit_maskInput_hi[12335:12320]},
     {loadUnit_maskInput_hi[12319:12304]},
     {loadUnit_maskInput_hi[12303:12288]},
     {loadUnit_maskInput_hi[12287:12272]},
     {loadUnit_maskInput_hi[12271:12256]},
     {loadUnit_maskInput_hi[12255:12240]},
     {loadUnit_maskInput_hi[12239:12224]},
     {loadUnit_maskInput_hi[12223:12208]},
     {loadUnit_maskInput_hi[12207:12192]},
     {loadUnit_maskInput_hi[12191:12176]},
     {loadUnit_maskInput_hi[12175:12160]},
     {loadUnit_maskInput_hi[12159:12144]},
     {loadUnit_maskInput_hi[12143:12128]},
     {loadUnit_maskInput_hi[12127:12112]},
     {loadUnit_maskInput_hi[12111:12096]},
     {loadUnit_maskInput_hi[12095:12080]},
     {loadUnit_maskInput_hi[12079:12064]},
     {loadUnit_maskInput_hi[12063:12048]},
     {loadUnit_maskInput_hi[12047:12032]},
     {loadUnit_maskInput_hi[12031:12016]},
     {loadUnit_maskInput_hi[12015:12000]},
     {loadUnit_maskInput_hi[11999:11984]},
     {loadUnit_maskInput_hi[11983:11968]},
     {loadUnit_maskInput_hi[11967:11952]},
     {loadUnit_maskInput_hi[11951:11936]},
     {loadUnit_maskInput_hi[11935:11920]},
     {loadUnit_maskInput_hi[11919:11904]},
     {loadUnit_maskInput_hi[11903:11888]},
     {loadUnit_maskInput_hi[11887:11872]},
     {loadUnit_maskInput_hi[11871:11856]},
     {loadUnit_maskInput_hi[11855:11840]},
     {loadUnit_maskInput_hi[11839:11824]},
     {loadUnit_maskInput_hi[11823:11808]},
     {loadUnit_maskInput_hi[11807:11792]},
     {loadUnit_maskInput_hi[11791:11776]},
     {loadUnit_maskInput_hi[11775:11760]},
     {loadUnit_maskInput_hi[11759:11744]},
     {loadUnit_maskInput_hi[11743:11728]},
     {loadUnit_maskInput_hi[11727:11712]},
     {loadUnit_maskInput_hi[11711:11696]},
     {loadUnit_maskInput_hi[11695:11680]},
     {loadUnit_maskInput_hi[11679:11664]},
     {loadUnit_maskInput_hi[11663:11648]},
     {loadUnit_maskInput_hi[11647:11632]},
     {loadUnit_maskInput_hi[11631:11616]},
     {loadUnit_maskInput_hi[11615:11600]},
     {loadUnit_maskInput_hi[11599:11584]},
     {loadUnit_maskInput_hi[11583:11568]},
     {loadUnit_maskInput_hi[11567:11552]},
     {loadUnit_maskInput_hi[11551:11536]},
     {loadUnit_maskInput_hi[11535:11520]},
     {loadUnit_maskInput_hi[11519:11504]},
     {loadUnit_maskInput_hi[11503:11488]},
     {loadUnit_maskInput_hi[11487:11472]},
     {loadUnit_maskInput_hi[11471:11456]},
     {loadUnit_maskInput_hi[11455:11440]},
     {loadUnit_maskInput_hi[11439:11424]},
     {loadUnit_maskInput_hi[11423:11408]},
     {loadUnit_maskInput_hi[11407:11392]},
     {loadUnit_maskInput_hi[11391:11376]},
     {loadUnit_maskInput_hi[11375:11360]},
     {loadUnit_maskInput_hi[11359:11344]},
     {loadUnit_maskInput_hi[11343:11328]},
     {loadUnit_maskInput_hi[11327:11312]},
     {loadUnit_maskInput_hi[11311:11296]},
     {loadUnit_maskInput_hi[11295:11280]},
     {loadUnit_maskInput_hi[11279:11264]},
     {loadUnit_maskInput_hi[11263:11248]},
     {loadUnit_maskInput_hi[11247:11232]},
     {loadUnit_maskInput_hi[11231:11216]},
     {loadUnit_maskInput_hi[11215:11200]},
     {loadUnit_maskInput_hi[11199:11184]},
     {loadUnit_maskInput_hi[11183:11168]},
     {loadUnit_maskInput_hi[11167:11152]},
     {loadUnit_maskInput_hi[11151:11136]},
     {loadUnit_maskInput_hi[11135:11120]},
     {loadUnit_maskInput_hi[11119:11104]},
     {loadUnit_maskInput_hi[11103:11088]},
     {loadUnit_maskInput_hi[11087:11072]},
     {loadUnit_maskInput_hi[11071:11056]},
     {loadUnit_maskInput_hi[11055:11040]},
     {loadUnit_maskInput_hi[11039:11024]},
     {loadUnit_maskInput_hi[11023:11008]},
     {loadUnit_maskInput_hi[11007:10992]},
     {loadUnit_maskInput_hi[10991:10976]},
     {loadUnit_maskInput_hi[10975:10960]},
     {loadUnit_maskInput_hi[10959:10944]},
     {loadUnit_maskInput_hi[10943:10928]},
     {loadUnit_maskInput_hi[10927:10912]},
     {loadUnit_maskInput_hi[10911:10896]},
     {loadUnit_maskInput_hi[10895:10880]},
     {loadUnit_maskInput_hi[10879:10864]},
     {loadUnit_maskInput_hi[10863:10848]},
     {loadUnit_maskInput_hi[10847:10832]},
     {loadUnit_maskInput_hi[10831:10816]},
     {loadUnit_maskInput_hi[10815:10800]},
     {loadUnit_maskInput_hi[10799:10784]},
     {loadUnit_maskInput_hi[10783:10768]},
     {loadUnit_maskInput_hi[10767:10752]},
     {loadUnit_maskInput_hi[10751:10736]},
     {loadUnit_maskInput_hi[10735:10720]},
     {loadUnit_maskInput_hi[10719:10704]},
     {loadUnit_maskInput_hi[10703:10688]},
     {loadUnit_maskInput_hi[10687:10672]},
     {loadUnit_maskInput_hi[10671:10656]},
     {loadUnit_maskInput_hi[10655:10640]},
     {loadUnit_maskInput_hi[10639:10624]},
     {loadUnit_maskInput_hi[10623:10608]},
     {loadUnit_maskInput_hi[10607:10592]},
     {loadUnit_maskInput_hi[10591:10576]},
     {loadUnit_maskInput_hi[10575:10560]},
     {loadUnit_maskInput_hi[10559:10544]},
     {loadUnit_maskInput_hi[10543:10528]},
     {loadUnit_maskInput_hi[10527:10512]},
     {loadUnit_maskInput_hi[10511:10496]},
     {loadUnit_maskInput_hi[10495:10480]},
     {loadUnit_maskInput_hi[10479:10464]},
     {loadUnit_maskInput_hi[10463:10448]},
     {loadUnit_maskInput_hi[10447:10432]},
     {loadUnit_maskInput_hi[10431:10416]},
     {loadUnit_maskInput_hi[10415:10400]},
     {loadUnit_maskInput_hi[10399:10384]},
     {loadUnit_maskInput_hi[10383:10368]},
     {loadUnit_maskInput_hi[10367:10352]},
     {loadUnit_maskInput_hi[10351:10336]},
     {loadUnit_maskInput_hi[10335:10320]},
     {loadUnit_maskInput_hi[10319:10304]},
     {loadUnit_maskInput_hi[10303:10288]},
     {loadUnit_maskInput_hi[10287:10272]},
     {loadUnit_maskInput_hi[10271:10256]},
     {loadUnit_maskInput_hi[10255:10240]},
     {loadUnit_maskInput_hi[10239:10224]},
     {loadUnit_maskInput_hi[10223:10208]},
     {loadUnit_maskInput_hi[10207:10192]},
     {loadUnit_maskInput_hi[10191:10176]},
     {loadUnit_maskInput_hi[10175:10160]},
     {loadUnit_maskInput_hi[10159:10144]},
     {loadUnit_maskInput_hi[10143:10128]},
     {loadUnit_maskInput_hi[10127:10112]},
     {loadUnit_maskInput_hi[10111:10096]},
     {loadUnit_maskInput_hi[10095:10080]},
     {loadUnit_maskInput_hi[10079:10064]},
     {loadUnit_maskInput_hi[10063:10048]},
     {loadUnit_maskInput_hi[10047:10032]},
     {loadUnit_maskInput_hi[10031:10016]},
     {loadUnit_maskInput_hi[10015:10000]},
     {loadUnit_maskInput_hi[9999:9984]},
     {loadUnit_maskInput_hi[9983:9968]},
     {loadUnit_maskInput_hi[9967:9952]},
     {loadUnit_maskInput_hi[9951:9936]},
     {loadUnit_maskInput_hi[9935:9920]},
     {loadUnit_maskInput_hi[9919:9904]},
     {loadUnit_maskInput_hi[9903:9888]},
     {loadUnit_maskInput_hi[9887:9872]},
     {loadUnit_maskInput_hi[9871:9856]},
     {loadUnit_maskInput_hi[9855:9840]},
     {loadUnit_maskInput_hi[9839:9824]},
     {loadUnit_maskInput_hi[9823:9808]},
     {loadUnit_maskInput_hi[9807:9792]},
     {loadUnit_maskInput_hi[9791:9776]},
     {loadUnit_maskInput_hi[9775:9760]},
     {loadUnit_maskInput_hi[9759:9744]},
     {loadUnit_maskInput_hi[9743:9728]},
     {loadUnit_maskInput_hi[9727:9712]},
     {loadUnit_maskInput_hi[9711:9696]},
     {loadUnit_maskInput_hi[9695:9680]},
     {loadUnit_maskInput_hi[9679:9664]},
     {loadUnit_maskInput_hi[9663:9648]},
     {loadUnit_maskInput_hi[9647:9632]},
     {loadUnit_maskInput_hi[9631:9616]},
     {loadUnit_maskInput_hi[9615:9600]},
     {loadUnit_maskInput_hi[9599:9584]},
     {loadUnit_maskInput_hi[9583:9568]},
     {loadUnit_maskInput_hi[9567:9552]},
     {loadUnit_maskInput_hi[9551:9536]},
     {loadUnit_maskInput_hi[9535:9520]},
     {loadUnit_maskInput_hi[9519:9504]},
     {loadUnit_maskInput_hi[9503:9488]},
     {loadUnit_maskInput_hi[9487:9472]},
     {loadUnit_maskInput_hi[9471:9456]},
     {loadUnit_maskInput_hi[9455:9440]},
     {loadUnit_maskInput_hi[9439:9424]},
     {loadUnit_maskInput_hi[9423:9408]},
     {loadUnit_maskInput_hi[9407:9392]},
     {loadUnit_maskInput_hi[9391:9376]},
     {loadUnit_maskInput_hi[9375:9360]},
     {loadUnit_maskInput_hi[9359:9344]},
     {loadUnit_maskInput_hi[9343:9328]},
     {loadUnit_maskInput_hi[9327:9312]},
     {loadUnit_maskInput_hi[9311:9296]},
     {loadUnit_maskInput_hi[9295:9280]},
     {loadUnit_maskInput_hi[9279:9264]},
     {loadUnit_maskInput_hi[9263:9248]},
     {loadUnit_maskInput_hi[9247:9232]},
     {loadUnit_maskInput_hi[9231:9216]},
     {loadUnit_maskInput_hi[9215:9200]},
     {loadUnit_maskInput_hi[9199:9184]},
     {loadUnit_maskInput_hi[9183:9168]},
     {loadUnit_maskInput_hi[9167:9152]},
     {loadUnit_maskInput_hi[9151:9136]},
     {loadUnit_maskInput_hi[9135:9120]},
     {loadUnit_maskInput_hi[9119:9104]},
     {loadUnit_maskInput_hi[9103:9088]},
     {loadUnit_maskInput_hi[9087:9072]},
     {loadUnit_maskInput_hi[9071:9056]},
     {loadUnit_maskInput_hi[9055:9040]},
     {loadUnit_maskInput_hi[9039:9024]},
     {loadUnit_maskInput_hi[9023:9008]},
     {loadUnit_maskInput_hi[9007:8992]},
     {loadUnit_maskInput_hi[8991:8976]},
     {loadUnit_maskInput_hi[8975:8960]},
     {loadUnit_maskInput_hi[8959:8944]},
     {loadUnit_maskInput_hi[8943:8928]},
     {loadUnit_maskInput_hi[8927:8912]},
     {loadUnit_maskInput_hi[8911:8896]},
     {loadUnit_maskInput_hi[8895:8880]},
     {loadUnit_maskInput_hi[8879:8864]},
     {loadUnit_maskInput_hi[8863:8848]},
     {loadUnit_maskInput_hi[8847:8832]},
     {loadUnit_maskInput_hi[8831:8816]},
     {loadUnit_maskInput_hi[8815:8800]},
     {loadUnit_maskInput_hi[8799:8784]},
     {loadUnit_maskInput_hi[8783:8768]},
     {loadUnit_maskInput_hi[8767:8752]},
     {loadUnit_maskInput_hi[8751:8736]},
     {loadUnit_maskInput_hi[8735:8720]},
     {loadUnit_maskInput_hi[8719:8704]},
     {loadUnit_maskInput_hi[8703:8688]},
     {loadUnit_maskInput_hi[8687:8672]},
     {loadUnit_maskInput_hi[8671:8656]},
     {loadUnit_maskInput_hi[8655:8640]},
     {loadUnit_maskInput_hi[8639:8624]},
     {loadUnit_maskInput_hi[8623:8608]},
     {loadUnit_maskInput_hi[8607:8592]},
     {loadUnit_maskInput_hi[8591:8576]},
     {loadUnit_maskInput_hi[8575:8560]},
     {loadUnit_maskInput_hi[8559:8544]},
     {loadUnit_maskInput_hi[8543:8528]},
     {loadUnit_maskInput_hi[8527:8512]},
     {loadUnit_maskInput_hi[8511:8496]},
     {loadUnit_maskInput_hi[8495:8480]},
     {loadUnit_maskInput_hi[8479:8464]},
     {loadUnit_maskInput_hi[8463:8448]},
     {loadUnit_maskInput_hi[8447:8432]},
     {loadUnit_maskInput_hi[8431:8416]},
     {loadUnit_maskInput_hi[8415:8400]},
     {loadUnit_maskInput_hi[8399:8384]},
     {loadUnit_maskInput_hi[8383:8368]},
     {loadUnit_maskInput_hi[8367:8352]},
     {loadUnit_maskInput_hi[8351:8336]},
     {loadUnit_maskInput_hi[8335:8320]},
     {loadUnit_maskInput_hi[8319:8304]},
     {loadUnit_maskInput_hi[8303:8288]},
     {loadUnit_maskInput_hi[8287:8272]},
     {loadUnit_maskInput_hi[8271:8256]},
     {loadUnit_maskInput_hi[8255:8240]},
     {loadUnit_maskInput_hi[8239:8224]},
     {loadUnit_maskInput_hi[8223:8208]},
     {loadUnit_maskInput_hi[8207:8192]},
     {loadUnit_maskInput_hi[8191:8176]},
     {loadUnit_maskInput_hi[8175:8160]},
     {loadUnit_maskInput_hi[8159:8144]},
     {loadUnit_maskInput_hi[8143:8128]},
     {loadUnit_maskInput_hi[8127:8112]},
     {loadUnit_maskInput_hi[8111:8096]},
     {loadUnit_maskInput_hi[8095:8080]},
     {loadUnit_maskInput_hi[8079:8064]},
     {loadUnit_maskInput_hi[8063:8048]},
     {loadUnit_maskInput_hi[8047:8032]},
     {loadUnit_maskInput_hi[8031:8016]},
     {loadUnit_maskInput_hi[8015:8000]},
     {loadUnit_maskInput_hi[7999:7984]},
     {loadUnit_maskInput_hi[7983:7968]},
     {loadUnit_maskInput_hi[7967:7952]},
     {loadUnit_maskInput_hi[7951:7936]},
     {loadUnit_maskInput_hi[7935:7920]},
     {loadUnit_maskInput_hi[7919:7904]},
     {loadUnit_maskInput_hi[7903:7888]},
     {loadUnit_maskInput_hi[7887:7872]},
     {loadUnit_maskInput_hi[7871:7856]},
     {loadUnit_maskInput_hi[7855:7840]},
     {loadUnit_maskInput_hi[7839:7824]},
     {loadUnit_maskInput_hi[7823:7808]},
     {loadUnit_maskInput_hi[7807:7792]},
     {loadUnit_maskInput_hi[7791:7776]},
     {loadUnit_maskInput_hi[7775:7760]},
     {loadUnit_maskInput_hi[7759:7744]},
     {loadUnit_maskInput_hi[7743:7728]},
     {loadUnit_maskInput_hi[7727:7712]},
     {loadUnit_maskInput_hi[7711:7696]},
     {loadUnit_maskInput_hi[7695:7680]},
     {loadUnit_maskInput_hi[7679:7664]},
     {loadUnit_maskInput_hi[7663:7648]},
     {loadUnit_maskInput_hi[7647:7632]},
     {loadUnit_maskInput_hi[7631:7616]},
     {loadUnit_maskInput_hi[7615:7600]},
     {loadUnit_maskInput_hi[7599:7584]},
     {loadUnit_maskInput_hi[7583:7568]},
     {loadUnit_maskInput_hi[7567:7552]},
     {loadUnit_maskInput_hi[7551:7536]},
     {loadUnit_maskInput_hi[7535:7520]},
     {loadUnit_maskInput_hi[7519:7504]},
     {loadUnit_maskInput_hi[7503:7488]},
     {loadUnit_maskInput_hi[7487:7472]},
     {loadUnit_maskInput_hi[7471:7456]},
     {loadUnit_maskInput_hi[7455:7440]},
     {loadUnit_maskInput_hi[7439:7424]},
     {loadUnit_maskInput_hi[7423:7408]},
     {loadUnit_maskInput_hi[7407:7392]},
     {loadUnit_maskInput_hi[7391:7376]},
     {loadUnit_maskInput_hi[7375:7360]},
     {loadUnit_maskInput_hi[7359:7344]},
     {loadUnit_maskInput_hi[7343:7328]},
     {loadUnit_maskInput_hi[7327:7312]},
     {loadUnit_maskInput_hi[7311:7296]},
     {loadUnit_maskInput_hi[7295:7280]},
     {loadUnit_maskInput_hi[7279:7264]},
     {loadUnit_maskInput_hi[7263:7248]},
     {loadUnit_maskInput_hi[7247:7232]},
     {loadUnit_maskInput_hi[7231:7216]},
     {loadUnit_maskInput_hi[7215:7200]},
     {loadUnit_maskInput_hi[7199:7184]},
     {loadUnit_maskInput_hi[7183:7168]},
     {loadUnit_maskInput_hi[7167:7152]},
     {loadUnit_maskInput_hi[7151:7136]},
     {loadUnit_maskInput_hi[7135:7120]},
     {loadUnit_maskInput_hi[7119:7104]},
     {loadUnit_maskInput_hi[7103:7088]},
     {loadUnit_maskInput_hi[7087:7072]},
     {loadUnit_maskInput_hi[7071:7056]},
     {loadUnit_maskInput_hi[7055:7040]},
     {loadUnit_maskInput_hi[7039:7024]},
     {loadUnit_maskInput_hi[7023:7008]},
     {loadUnit_maskInput_hi[7007:6992]},
     {loadUnit_maskInput_hi[6991:6976]},
     {loadUnit_maskInput_hi[6975:6960]},
     {loadUnit_maskInput_hi[6959:6944]},
     {loadUnit_maskInput_hi[6943:6928]},
     {loadUnit_maskInput_hi[6927:6912]},
     {loadUnit_maskInput_hi[6911:6896]},
     {loadUnit_maskInput_hi[6895:6880]},
     {loadUnit_maskInput_hi[6879:6864]},
     {loadUnit_maskInput_hi[6863:6848]},
     {loadUnit_maskInput_hi[6847:6832]},
     {loadUnit_maskInput_hi[6831:6816]},
     {loadUnit_maskInput_hi[6815:6800]},
     {loadUnit_maskInput_hi[6799:6784]},
     {loadUnit_maskInput_hi[6783:6768]},
     {loadUnit_maskInput_hi[6767:6752]},
     {loadUnit_maskInput_hi[6751:6736]},
     {loadUnit_maskInput_hi[6735:6720]},
     {loadUnit_maskInput_hi[6719:6704]},
     {loadUnit_maskInput_hi[6703:6688]},
     {loadUnit_maskInput_hi[6687:6672]},
     {loadUnit_maskInput_hi[6671:6656]},
     {loadUnit_maskInput_hi[6655:6640]},
     {loadUnit_maskInput_hi[6639:6624]},
     {loadUnit_maskInput_hi[6623:6608]},
     {loadUnit_maskInput_hi[6607:6592]},
     {loadUnit_maskInput_hi[6591:6576]},
     {loadUnit_maskInput_hi[6575:6560]},
     {loadUnit_maskInput_hi[6559:6544]},
     {loadUnit_maskInput_hi[6543:6528]},
     {loadUnit_maskInput_hi[6527:6512]},
     {loadUnit_maskInput_hi[6511:6496]},
     {loadUnit_maskInput_hi[6495:6480]},
     {loadUnit_maskInput_hi[6479:6464]},
     {loadUnit_maskInput_hi[6463:6448]},
     {loadUnit_maskInput_hi[6447:6432]},
     {loadUnit_maskInput_hi[6431:6416]},
     {loadUnit_maskInput_hi[6415:6400]},
     {loadUnit_maskInput_hi[6399:6384]},
     {loadUnit_maskInput_hi[6383:6368]},
     {loadUnit_maskInput_hi[6367:6352]},
     {loadUnit_maskInput_hi[6351:6336]},
     {loadUnit_maskInput_hi[6335:6320]},
     {loadUnit_maskInput_hi[6319:6304]},
     {loadUnit_maskInput_hi[6303:6288]},
     {loadUnit_maskInput_hi[6287:6272]},
     {loadUnit_maskInput_hi[6271:6256]},
     {loadUnit_maskInput_hi[6255:6240]},
     {loadUnit_maskInput_hi[6239:6224]},
     {loadUnit_maskInput_hi[6223:6208]},
     {loadUnit_maskInput_hi[6207:6192]},
     {loadUnit_maskInput_hi[6191:6176]},
     {loadUnit_maskInput_hi[6175:6160]},
     {loadUnit_maskInput_hi[6159:6144]},
     {loadUnit_maskInput_hi[6143:6128]},
     {loadUnit_maskInput_hi[6127:6112]},
     {loadUnit_maskInput_hi[6111:6096]},
     {loadUnit_maskInput_hi[6095:6080]},
     {loadUnit_maskInput_hi[6079:6064]},
     {loadUnit_maskInput_hi[6063:6048]},
     {loadUnit_maskInput_hi[6047:6032]},
     {loadUnit_maskInput_hi[6031:6016]},
     {loadUnit_maskInput_hi[6015:6000]},
     {loadUnit_maskInput_hi[5999:5984]},
     {loadUnit_maskInput_hi[5983:5968]},
     {loadUnit_maskInput_hi[5967:5952]},
     {loadUnit_maskInput_hi[5951:5936]},
     {loadUnit_maskInput_hi[5935:5920]},
     {loadUnit_maskInput_hi[5919:5904]},
     {loadUnit_maskInput_hi[5903:5888]},
     {loadUnit_maskInput_hi[5887:5872]},
     {loadUnit_maskInput_hi[5871:5856]},
     {loadUnit_maskInput_hi[5855:5840]},
     {loadUnit_maskInput_hi[5839:5824]},
     {loadUnit_maskInput_hi[5823:5808]},
     {loadUnit_maskInput_hi[5807:5792]},
     {loadUnit_maskInput_hi[5791:5776]},
     {loadUnit_maskInput_hi[5775:5760]},
     {loadUnit_maskInput_hi[5759:5744]},
     {loadUnit_maskInput_hi[5743:5728]},
     {loadUnit_maskInput_hi[5727:5712]},
     {loadUnit_maskInput_hi[5711:5696]},
     {loadUnit_maskInput_hi[5695:5680]},
     {loadUnit_maskInput_hi[5679:5664]},
     {loadUnit_maskInput_hi[5663:5648]},
     {loadUnit_maskInput_hi[5647:5632]},
     {loadUnit_maskInput_hi[5631:5616]},
     {loadUnit_maskInput_hi[5615:5600]},
     {loadUnit_maskInput_hi[5599:5584]},
     {loadUnit_maskInput_hi[5583:5568]},
     {loadUnit_maskInput_hi[5567:5552]},
     {loadUnit_maskInput_hi[5551:5536]},
     {loadUnit_maskInput_hi[5535:5520]},
     {loadUnit_maskInput_hi[5519:5504]},
     {loadUnit_maskInput_hi[5503:5488]},
     {loadUnit_maskInput_hi[5487:5472]},
     {loadUnit_maskInput_hi[5471:5456]},
     {loadUnit_maskInput_hi[5455:5440]},
     {loadUnit_maskInput_hi[5439:5424]},
     {loadUnit_maskInput_hi[5423:5408]},
     {loadUnit_maskInput_hi[5407:5392]},
     {loadUnit_maskInput_hi[5391:5376]},
     {loadUnit_maskInput_hi[5375:5360]},
     {loadUnit_maskInput_hi[5359:5344]},
     {loadUnit_maskInput_hi[5343:5328]},
     {loadUnit_maskInput_hi[5327:5312]},
     {loadUnit_maskInput_hi[5311:5296]},
     {loadUnit_maskInput_hi[5295:5280]},
     {loadUnit_maskInput_hi[5279:5264]},
     {loadUnit_maskInput_hi[5263:5248]},
     {loadUnit_maskInput_hi[5247:5232]},
     {loadUnit_maskInput_hi[5231:5216]},
     {loadUnit_maskInput_hi[5215:5200]},
     {loadUnit_maskInput_hi[5199:5184]},
     {loadUnit_maskInput_hi[5183:5168]},
     {loadUnit_maskInput_hi[5167:5152]},
     {loadUnit_maskInput_hi[5151:5136]},
     {loadUnit_maskInput_hi[5135:5120]},
     {loadUnit_maskInput_hi[5119:5104]},
     {loadUnit_maskInput_hi[5103:5088]},
     {loadUnit_maskInput_hi[5087:5072]},
     {loadUnit_maskInput_hi[5071:5056]},
     {loadUnit_maskInput_hi[5055:5040]},
     {loadUnit_maskInput_hi[5039:5024]},
     {loadUnit_maskInput_hi[5023:5008]},
     {loadUnit_maskInput_hi[5007:4992]},
     {loadUnit_maskInput_hi[4991:4976]},
     {loadUnit_maskInput_hi[4975:4960]},
     {loadUnit_maskInput_hi[4959:4944]},
     {loadUnit_maskInput_hi[4943:4928]},
     {loadUnit_maskInput_hi[4927:4912]},
     {loadUnit_maskInput_hi[4911:4896]},
     {loadUnit_maskInput_hi[4895:4880]},
     {loadUnit_maskInput_hi[4879:4864]},
     {loadUnit_maskInput_hi[4863:4848]},
     {loadUnit_maskInput_hi[4847:4832]},
     {loadUnit_maskInput_hi[4831:4816]},
     {loadUnit_maskInput_hi[4815:4800]},
     {loadUnit_maskInput_hi[4799:4784]},
     {loadUnit_maskInput_hi[4783:4768]},
     {loadUnit_maskInput_hi[4767:4752]},
     {loadUnit_maskInput_hi[4751:4736]},
     {loadUnit_maskInput_hi[4735:4720]},
     {loadUnit_maskInput_hi[4719:4704]},
     {loadUnit_maskInput_hi[4703:4688]},
     {loadUnit_maskInput_hi[4687:4672]},
     {loadUnit_maskInput_hi[4671:4656]},
     {loadUnit_maskInput_hi[4655:4640]},
     {loadUnit_maskInput_hi[4639:4624]},
     {loadUnit_maskInput_hi[4623:4608]},
     {loadUnit_maskInput_hi[4607:4592]},
     {loadUnit_maskInput_hi[4591:4576]},
     {loadUnit_maskInput_hi[4575:4560]},
     {loadUnit_maskInput_hi[4559:4544]},
     {loadUnit_maskInput_hi[4543:4528]},
     {loadUnit_maskInput_hi[4527:4512]},
     {loadUnit_maskInput_hi[4511:4496]},
     {loadUnit_maskInput_hi[4495:4480]},
     {loadUnit_maskInput_hi[4479:4464]},
     {loadUnit_maskInput_hi[4463:4448]},
     {loadUnit_maskInput_hi[4447:4432]},
     {loadUnit_maskInput_hi[4431:4416]},
     {loadUnit_maskInput_hi[4415:4400]},
     {loadUnit_maskInput_hi[4399:4384]},
     {loadUnit_maskInput_hi[4383:4368]},
     {loadUnit_maskInput_hi[4367:4352]},
     {loadUnit_maskInput_hi[4351:4336]},
     {loadUnit_maskInput_hi[4335:4320]},
     {loadUnit_maskInput_hi[4319:4304]},
     {loadUnit_maskInput_hi[4303:4288]},
     {loadUnit_maskInput_hi[4287:4272]},
     {loadUnit_maskInput_hi[4271:4256]},
     {loadUnit_maskInput_hi[4255:4240]},
     {loadUnit_maskInput_hi[4239:4224]},
     {loadUnit_maskInput_hi[4223:4208]},
     {loadUnit_maskInput_hi[4207:4192]},
     {loadUnit_maskInput_hi[4191:4176]},
     {loadUnit_maskInput_hi[4175:4160]},
     {loadUnit_maskInput_hi[4159:4144]},
     {loadUnit_maskInput_hi[4143:4128]},
     {loadUnit_maskInput_hi[4127:4112]},
     {loadUnit_maskInput_hi[4111:4096]},
     {loadUnit_maskInput_hi[4095:4080]},
     {loadUnit_maskInput_hi[4079:4064]},
     {loadUnit_maskInput_hi[4063:4048]},
     {loadUnit_maskInput_hi[4047:4032]},
     {loadUnit_maskInput_hi[4031:4016]},
     {loadUnit_maskInput_hi[4015:4000]},
     {loadUnit_maskInput_hi[3999:3984]},
     {loadUnit_maskInput_hi[3983:3968]},
     {loadUnit_maskInput_hi[3967:3952]},
     {loadUnit_maskInput_hi[3951:3936]},
     {loadUnit_maskInput_hi[3935:3920]},
     {loadUnit_maskInput_hi[3919:3904]},
     {loadUnit_maskInput_hi[3903:3888]},
     {loadUnit_maskInput_hi[3887:3872]},
     {loadUnit_maskInput_hi[3871:3856]},
     {loadUnit_maskInput_hi[3855:3840]},
     {loadUnit_maskInput_hi[3839:3824]},
     {loadUnit_maskInput_hi[3823:3808]},
     {loadUnit_maskInput_hi[3807:3792]},
     {loadUnit_maskInput_hi[3791:3776]},
     {loadUnit_maskInput_hi[3775:3760]},
     {loadUnit_maskInput_hi[3759:3744]},
     {loadUnit_maskInput_hi[3743:3728]},
     {loadUnit_maskInput_hi[3727:3712]},
     {loadUnit_maskInput_hi[3711:3696]},
     {loadUnit_maskInput_hi[3695:3680]},
     {loadUnit_maskInput_hi[3679:3664]},
     {loadUnit_maskInput_hi[3663:3648]},
     {loadUnit_maskInput_hi[3647:3632]},
     {loadUnit_maskInput_hi[3631:3616]},
     {loadUnit_maskInput_hi[3615:3600]},
     {loadUnit_maskInput_hi[3599:3584]},
     {loadUnit_maskInput_hi[3583:3568]},
     {loadUnit_maskInput_hi[3567:3552]},
     {loadUnit_maskInput_hi[3551:3536]},
     {loadUnit_maskInput_hi[3535:3520]},
     {loadUnit_maskInput_hi[3519:3504]},
     {loadUnit_maskInput_hi[3503:3488]},
     {loadUnit_maskInput_hi[3487:3472]},
     {loadUnit_maskInput_hi[3471:3456]},
     {loadUnit_maskInput_hi[3455:3440]},
     {loadUnit_maskInput_hi[3439:3424]},
     {loadUnit_maskInput_hi[3423:3408]},
     {loadUnit_maskInput_hi[3407:3392]},
     {loadUnit_maskInput_hi[3391:3376]},
     {loadUnit_maskInput_hi[3375:3360]},
     {loadUnit_maskInput_hi[3359:3344]},
     {loadUnit_maskInput_hi[3343:3328]},
     {loadUnit_maskInput_hi[3327:3312]},
     {loadUnit_maskInput_hi[3311:3296]},
     {loadUnit_maskInput_hi[3295:3280]},
     {loadUnit_maskInput_hi[3279:3264]},
     {loadUnit_maskInput_hi[3263:3248]},
     {loadUnit_maskInput_hi[3247:3232]},
     {loadUnit_maskInput_hi[3231:3216]},
     {loadUnit_maskInput_hi[3215:3200]},
     {loadUnit_maskInput_hi[3199:3184]},
     {loadUnit_maskInput_hi[3183:3168]},
     {loadUnit_maskInput_hi[3167:3152]},
     {loadUnit_maskInput_hi[3151:3136]},
     {loadUnit_maskInput_hi[3135:3120]},
     {loadUnit_maskInput_hi[3119:3104]},
     {loadUnit_maskInput_hi[3103:3088]},
     {loadUnit_maskInput_hi[3087:3072]},
     {loadUnit_maskInput_hi[3071:3056]},
     {loadUnit_maskInput_hi[3055:3040]},
     {loadUnit_maskInput_hi[3039:3024]},
     {loadUnit_maskInput_hi[3023:3008]},
     {loadUnit_maskInput_hi[3007:2992]},
     {loadUnit_maskInput_hi[2991:2976]},
     {loadUnit_maskInput_hi[2975:2960]},
     {loadUnit_maskInput_hi[2959:2944]},
     {loadUnit_maskInput_hi[2943:2928]},
     {loadUnit_maskInput_hi[2927:2912]},
     {loadUnit_maskInput_hi[2911:2896]},
     {loadUnit_maskInput_hi[2895:2880]},
     {loadUnit_maskInput_hi[2879:2864]},
     {loadUnit_maskInput_hi[2863:2848]},
     {loadUnit_maskInput_hi[2847:2832]},
     {loadUnit_maskInput_hi[2831:2816]},
     {loadUnit_maskInput_hi[2815:2800]},
     {loadUnit_maskInput_hi[2799:2784]},
     {loadUnit_maskInput_hi[2783:2768]},
     {loadUnit_maskInput_hi[2767:2752]},
     {loadUnit_maskInput_hi[2751:2736]},
     {loadUnit_maskInput_hi[2735:2720]},
     {loadUnit_maskInput_hi[2719:2704]},
     {loadUnit_maskInput_hi[2703:2688]},
     {loadUnit_maskInput_hi[2687:2672]},
     {loadUnit_maskInput_hi[2671:2656]},
     {loadUnit_maskInput_hi[2655:2640]},
     {loadUnit_maskInput_hi[2639:2624]},
     {loadUnit_maskInput_hi[2623:2608]},
     {loadUnit_maskInput_hi[2607:2592]},
     {loadUnit_maskInput_hi[2591:2576]},
     {loadUnit_maskInput_hi[2575:2560]},
     {loadUnit_maskInput_hi[2559:2544]},
     {loadUnit_maskInput_hi[2543:2528]},
     {loadUnit_maskInput_hi[2527:2512]},
     {loadUnit_maskInput_hi[2511:2496]},
     {loadUnit_maskInput_hi[2495:2480]},
     {loadUnit_maskInput_hi[2479:2464]},
     {loadUnit_maskInput_hi[2463:2448]},
     {loadUnit_maskInput_hi[2447:2432]},
     {loadUnit_maskInput_hi[2431:2416]},
     {loadUnit_maskInput_hi[2415:2400]},
     {loadUnit_maskInput_hi[2399:2384]},
     {loadUnit_maskInput_hi[2383:2368]},
     {loadUnit_maskInput_hi[2367:2352]},
     {loadUnit_maskInput_hi[2351:2336]},
     {loadUnit_maskInput_hi[2335:2320]},
     {loadUnit_maskInput_hi[2319:2304]},
     {loadUnit_maskInput_hi[2303:2288]},
     {loadUnit_maskInput_hi[2287:2272]},
     {loadUnit_maskInput_hi[2271:2256]},
     {loadUnit_maskInput_hi[2255:2240]},
     {loadUnit_maskInput_hi[2239:2224]},
     {loadUnit_maskInput_hi[2223:2208]},
     {loadUnit_maskInput_hi[2207:2192]},
     {loadUnit_maskInput_hi[2191:2176]},
     {loadUnit_maskInput_hi[2175:2160]},
     {loadUnit_maskInput_hi[2159:2144]},
     {loadUnit_maskInput_hi[2143:2128]},
     {loadUnit_maskInput_hi[2127:2112]},
     {loadUnit_maskInput_hi[2111:2096]},
     {loadUnit_maskInput_hi[2095:2080]},
     {loadUnit_maskInput_hi[2079:2064]},
     {loadUnit_maskInput_hi[2063:2048]},
     {loadUnit_maskInput_hi[2047:2032]},
     {loadUnit_maskInput_hi[2031:2016]},
     {loadUnit_maskInput_hi[2015:2000]},
     {loadUnit_maskInput_hi[1999:1984]},
     {loadUnit_maskInput_hi[1983:1968]},
     {loadUnit_maskInput_hi[1967:1952]},
     {loadUnit_maskInput_hi[1951:1936]},
     {loadUnit_maskInput_hi[1935:1920]},
     {loadUnit_maskInput_hi[1919:1904]},
     {loadUnit_maskInput_hi[1903:1888]},
     {loadUnit_maskInput_hi[1887:1872]},
     {loadUnit_maskInput_hi[1871:1856]},
     {loadUnit_maskInput_hi[1855:1840]},
     {loadUnit_maskInput_hi[1839:1824]},
     {loadUnit_maskInput_hi[1823:1808]},
     {loadUnit_maskInput_hi[1807:1792]},
     {loadUnit_maskInput_hi[1791:1776]},
     {loadUnit_maskInput_hi[1775:1760]},
     {loadUnit_maskInput_hi[1759:1744]},
     {loadUnit_maskInput_hi[1743:1728]},
     {loadUnit_maskInput_hi[1727:1712]},
     {loadUnit_maskInput_hi[1711:1696]},
     {loadUnit_maskInput_hi[1695:1680]},
     {loadUnit_maskInput_hi[1679:1664]},
     {loadUnit_maskInput_hi[1663:1648]},
     {loadUnit_maskInput_hi[1647:1632]},
     {loadUnit_maskInput_hi[1631:1616]},
     {loadUnit_maskInput_hi[1615:1600]},
     {loadUnit_maskInput_hi[1599:1584]},
     {loadUnit_maskInput_hi[1583:1568]},
     {loadUnit_maskInput_hi[1567:1552]},
     {loadUnit_maskInput_hi[1551:1536]},
     {loadUnit_maskInput_hi[1535:1520]},
     {loadUnit_maskInput_hi[1519:1504]},
     {loadUnit_maskInput_hi[1503:1488]},
     {loadUnit_maskInput_hi[1487:1472]},
     {loadUnit_maskInput_hi[1471:1456]},
     {loadUnit_maskInput_hi[1455:1440]},
     {loadUnit_maskInput_hi[1439:1424]},
     {loadUnit_maskInput_hi[1423:1408]},
     {loadUnit_maskInput_hi[1407:1392]},
     {loadUnit_maskInput_hi[1391:1376]},
     {loadUnit_maskInput_hi[1375:1360]},
     {loadUnit_maskInput_hi[1359:1344]},
     {loadUnit_maskInput_hi[1343:1328]},
     {loadUnit_maskInput_hi[1327:1312]},
     {loadUnit_maskInput_hi[1311:1296]},
     {loadUnit_maskInput_hi[1295:1280]},
     {loadUnit_maskInput_hi[1279:1264]},
     {loadUnit_maskInput_hi[1263:1248]},
     {loadUnit_maskInput_hi[1247:1232]},
     {loadUnit_maskInput_hi[1231:1216]},
     {loadUnit_maskInput_hi[1215:1200]},
     {loadUnit_maskInput_hi[1199:1184]},
     {loadUnit_maskInput_hi[1183:1168]},
     {loadUnit_maskInput_hi[1167:1152]},
     {loadUnit_maskInput_hi[1151:1136]},
     {loadUnit_maskInput_hi[1135:1120]},
     {loadUnit_maskInput_hi[1119:1104]},
     {loadUnit_maskInput_hi[1103:1088]},
     {loadUnit_maskInput_hi[1087:1072]},
     {loadUnit_maskInput_hi[1071:1056]},
     {loadUnit_maskInput_hi[1055:1040]},
     {loadUnit_maskInput_hi[1039:1024]},
     {loadUnit_maskInput_hi[1023:1008]},
     {loadUnit_maskInput_hi[1007:992]},
     {loadUnit_maskInput_hi[991:976]},
     {loadUnit_maskInput_hi[975:960]},
     {loadUnit_maskInput_hi[959:944]},
     {loadUnit_maskInput_hi[943:928]},
     {loadUnit_maskInput_hi[927:912]},
     {loadUnit_maskInput_hi[911:896]},
     {loadUnit_maskInput_hi[895:880]},
     {loadUnit_maskInput_hi[879:864]},
     {loadUnit_maskInput_hi[863:848]},
     {loadUnit_maskInput_hi[847:832]},
     {loadUnit_maskInput_hi[831:816]},
     {loadUnit_maskInput_hi[815:800]},
     {loadUnit_maskInput_hi[799:784]},
     {loadUnit_maskInput_hi[783:768]},
     {loadUnit_maskInput_hi[767:752]},
     {loadUnit_maskInput_hi[751:736]},
     {loadUnit_maskInput_hi[735:720]},
     {loadUnit_maskInput_hi[719:704]},
     {loadUnit_maskInput_hi[703:688]},
     {loadUnit_maskInput_hi[687:672]},
     {loadUnit_maskInput_hi[671:656]},
     {loadUnit_maskInput_hi[655:640]},
     {loadUnit_maskInput_hi[639:624]},
     {loadUnit_maskInput_hi[623:608]},
     {loadUnit_maskInput_hi[607:592]},
     {loadUnit_maskInput_hi[591:576]},
     {loadUnit_maskInput_hi[575:560]},
     {loadUnit_maskInput_hi[559:544]},
     {loadUnit_maskInput_hi[543:528]},
     {loadUnit_maskInput_hi[527:512]},
     {loadUnit_maskInput_hi[511:496]},
     {loadUnit_maskInput_hi[495:480]},
     {loadUnit_maskInput_hi[479:464]},
     {loadUnit_maskInput_hi[463:448]},
     {loadUnit_maskInput_hi[447:432]},
     {loadUnit_maskInput_hi[431:416]},
     {loadUnit_maskInput_hi[415:400]},
     {loadUnit_maskInput_hi[399:384]},
     {loadUnit_maskInput_hi[383:368]},
     {loadUnit_maskInput_hi[367:352]},
     {loadUnit_maskInput_hi[351:336]},
     {loadUnit_maskInput_hi[335:320]},
     {loadUnit_maskInput_hi[319:304]},
     {loadUnit_maskInput_hi[303:288]},
     {loadUnit_maskInput_hi[287:272]},
     {loadUnit_maskInput_hi[271:256]},
     {loadUnit_maskInput_hi[255:240]},
     {loadUnit_maskInput_hi[239:224]},
     {loadUnit_maskInput_hi[223:208]},
     {loadUnit_maskInput_hi[207:192]},
     {loadUnit_maskInput_hi[191:176]},
     {loadUnit_maskInput_hi[175:160]},
     {loadUnit_maskInput_hi[159:144]},
     {loadUnit_maskInput_hi[143:128]},
     {loadUnit_maskInput_hi[127:112]},
     {loadUnit_maskInput_hi[111:96]},
     {loadUnit_maskInput_hi[95:80]},
     {loadUnit_maskInput_hi[79:64]},
     {loadUnit_maskInput_hi[63:48]},
     {loadUnit_maskInput_hi[47:32]},
     {loadUnit_maskInput_hi[31:16]},
     {loadUnit_maskInput_hi[15:0]},
     {loadUnit_maskInput_lo[32767:32752]},
     {loadUnit_maskInput_lo[32751:32736]},
     {loadUnit_maskInput_lo[32735:32720]},
     {loadUnit_maskInput_lo[32719:32704]},
     {loadUnit_maskInput_lo[32703:32688]},
     {loadUnit_maskInput_lo[32687:32672]},
     {loadUnit_maskInput_lo[32671:32656]},
     {loadUnit_maskInput_lo[32655:32640]},
     {loadUnit_maskInput_lo[32639:32624]},
     {loadUnit_maskInput_lo[32623:32608]},
     {loadUnit_maskInput_lo[32607:32592]},
     {loadUnit_maskInput_lo[32591:32576]},
     {loadUnit_maskInput_lo[32575:32560]},
     {loadUnit_maskInput_lo[32559:32544]},
     {loadUnit_maskInput_lo[32543:32528]},
     {loadUnit_maskInput_lo[32527:32512]},
     {loadUnit_maskInput_lo[32511:32496]},
     {loadUnit_maskInput_lo[32495:32480]},
     {loadUnit_maskInput_lo[32479:32464]},
     {loadUnit_maskInput_lo[32463:32448]},
     {loadUnit_maskInput_lo[32447:32432]},
     {loadUnit_maskInput_lo[32431:32416]},
     {loadUnit_maskInput_lo[32415:32400]},
     {loadUnit_maskInput_lo[32399:32384]},
     {loadUnit_maskInput_lo[32383:32368]},
     {loadUnit_maskInput_lo[32367:32352]},
     {loadUnit_maskInput_lo[32351:32336]},
     {loadUnit_maskInput_lo[32335:32320]},
     {loadUnit_maskInput_lo[32319:32304]},
     {loadUnit_maskInput_lo[32303:32288]},
     {loadUnit_maskInput_lo[32287:32272]},
     {loadUnit_maskInput_lo[32271:32256]},
     {loadUnit_maskInput_lo[32255:32240]},
     {loadUnit_maskInput_lo[32239:32224]},
     {loadUnit_maskInput_lo[32223:32208]},
     {loadUnit_maskInput_lo[32207:32192]},
     {loadUnit_maskInput_lo[32191:32176]},
     {loadUnit_maskInput_lo[32175:32160]},
     {loadUnit_maskInput_lo[32159:32144]},
     {loadUnit_maskInput_lo[32143:32128]},
     {loadUnit_maskInput_lo[32127:32112]},
     {loadUnit_maskInput_lo[32111:32096]},
     {loadUnit_maskInput_lo[32095:32080]},
     {loadUnit_maskInput_lo[32079:32064]},
     {loadUnit_maskInput_lo[32063:32048]},
     {loadUnit_maskInput_lo[32047:32032]},
     {loadUnit_maskInput_lo[32031:32016]},
     {loadUnit_maskInput_lo[32015:32000]},
     {loadUnit_maskInput_lo[31999:31984]},
     {loadUnit_maskInput_lo[31983:31968]},
     {loadUnit_maskInput_lo[31967:31952]},
     {loadUnit_maskInput_lo[31951:31936]},
     {loadUnit_maskInput_lo[31935:31920]},
     {loadUnit_maskInput_lo[31919:31904]},
     {loadUnit_maskInput_lo[31903:31888]},
     {loadUnit_maskInput_lo[31887:31872]},
     {loadUnit_maskInput_lo[31871:31856]},
     {loadUnit_maskInput_lo[31855:31840]},
     {loadUnit_maskInput_lo[31839:31824]},
     {loadUnit_maskInput_lo[31823:31808]},
     {loadUnit_maskInput_lo[31807:31792]},
     {loadUnit_maskInput_lo[31791:31776]},
     {loadUnit_maskInput_lo[31775:31760]},
     {loadUnit_maskInput_lo[31759:31744]},
     {loadUnit_maskInput_lo[31743:31728]},
     {loadUnit_maskInput_lo[31727:31712]},
     {loadUnit_maskInput_lo[31711:31696]},
     {loadUnit_maskInput_lo[31695:31680]},
     {loadUnit_maskInput_lo[31679:31664]},
     {loadUnit_maskInput_lo[31663:31648]},
     {loadUnit_maskInput_lo[31647:31632]},
     {loadUnit_maskInput_lo[31631:31616]},
     {loadUnit_maskInput_lo[31615:31600]},
     {loadUnit_maskInput_lo[31599:31584]},
     {loadUnit_maskInput_lo[31583:31568]},
     {loadUnit_maskInput_lo[31567:31552]},
     {loadUnit_maskInput_lo[31551:31536]},
     {loadUnit_maskInput_lo[31535:31520]},
     {loadUnit_maskInput_lo[31519:31504]},
     {loadUnit_maskInput_lo[31503:31488]},
     {loadUnit_maskInput_lo[31487:31472]},
     {loadUnit_maskInput_lo[31471:31456]},
     {loadUnit_maskInput_lo[31455:31440]},
     {loadUnit_maskInput_lo[31439:31424]},
     {loadUnit_maskInput_lo[31423:31408]},
     {loadUnit_maskInput_lo[31407:31392]},
     {loadUnit_maskInput_lo[31391:31376]},
     {loadUnit_maskInput_lo[31375:31360]},
     {loadUnit_maskInput_lo[31359:31344]},
     {loadUnit_maskInput_lo[31343:31328]},
     {loadUnit_maskInput_lo[31327:31312]},
     {loadUnit_maskInput_lo[31311:31296]},
     {loadUnit_maskInput_lo[31295:31280]},
     {loadUnit_maskInput_lo[31279:31264]},
     {loadUnit_maskInput_lo[31263:31248]},
     {loadUnit_maskInput_lo[31247:31232]},
     {loadUnit_maskInput_lo[31231:31216]},
     {loadUnit_maskInput_lo[31215:31200]},
     {loadUnit_maskInput_lo[31199:31184]},
     {loadUnit_maskInput_lo[31183:31168]},
     {loadUnit_maskInput_lo[31167:31152]},
     {loadUnit_maskInput_lo[31151:31136]},
     {loadUnit_maskInput_lo[31135:31120]},
     {loadUnit_maskInput_lo[31119:31104]},
     {loadUnit_maskInput_lo[31103:31088]},
     {loadUnit_maskInput_lo[31087:31072]},
     {loadUnit_maskInput_lo[31071:31056]},
     {loadUnit_maskInput_lo[31055:31040]},
     {loadUnit_maskInput_lo[31039:31024]},
     {loadUnit_maskInput_lo[31023:31008]},
     {loadUnit_maskInput_lo[31007:30992]},
     {loadUnit_maskInput_lo[30991:30976]},
     {loadUnit_maskInput_lo[30975:30960]},
     {loadUnit_maskInput_lo[30959:30944]},
     {loadUnit_maskInput_lo[30943:30928]},
     {loadUnit_maskInput_lo[30927:30912]},
     {loadUnit_maskInput_lo[30911:30896]},
     {loadUnit_maskInput_lo[30895:30880]},
     {loadUnit_maskInput_lo[30879:30864]},
     {loadUnit_maskInput_lo[30863:30848]},
     {loadUnit_maskInput_lo[30847:30832]},
     {loadUnit_maskInput_lo[30831:30816]},
     {loadUnit_maskInput_lo[30815:30800]},
     {loadUnit_maskInput_lo[30799:30784]},
     {loadUnit_maskInput_lo[30783:30768]},
     {loadUnit_maskInput_lo[30767:30752]},
     {loadUnit_maskInput_lo[30751:30736]},
     {loadUnit_maskInput_lo[30735:30720]},
     {loadUnit_maskInput_lo[30719:30704]},
     {loadUnit_maskInput_lo[30703:30688]},
     {loadUnit_maskInput_lo[30687:30672]},
     {loadUnit_maskInput_lo[30671:30656]},
     {loadUnit_maskInput_lo[30655:30640]},
     {loadUnit_maskInput_lo[30639:30624]},
     {loadUnit_maskInput_lo[30623:30608]},
     {loadUnit_maskInput_lo[30607:30592]},
     {loadUnit_maskInput_lo[30591:30576]},
     {loadUnit_maskInput_lo[30575:30560]},
     {loadUnit_maskInput_lo[30559:30544]},
     {loadUnit_maskInput_lo[30543:30528]},
     {loadUnit_maskInput_lo[30527:30512]},
     {loadUnit_maskInput_lo[30511:30496]},
     {loadUnit_maskInput_lo[30495:30480]},
     {loadUnit_maskInput_lo[30479:30464]},
     {loadUnit_maskInput_lo[30463:30448]},
     {loadUnit_maskInput_lo[30447:30432]},
     {loadUnit_maskInput_lo[30431:30416]},
     {loadUnit_maskInput_lo[30415:30400]},
     {loadUnit_maskInput_lo[30399:30384]},
     {loadUnit_maskInput_lo[30383:30368]},
     {loadUnit_maskInput_lo[30367:30352]},
     {loadUnit_maskInput_lo[30351:30336]},
     {loadUnit_maskInput_lo[30335:30320]},
     {loadUnit_maskInput_lo[30319:30304]},
     {loadUnit_maskInput_lo[30303:30288]},
     {loadUnit_maskInput_lo[30287:30272]},
     {loadUnit_maskInput_lo[30271:30256]},
     {loadUnit_maskInput_lo[30255:30240]},
     {loadUnit_maskInput_lo[30239:30224]},
     {loadUnit_maskInput_lo[30223:30208]},
     {loadUnit_maskInput_lo[30207:30192]},
     {loadUnit_maskInput_lo[30191:30176]},
     {loadUnit_maskInput_lo[30175:30160]},
     {loadUnit_maskInput_lo[30159:30144]},
     {loadUnit_maskInput_lo[30143:30128]},
     {loadUnit_maskInput_lo[30127:30112]},
     {loadUnit_maskInput_lo[30111:30096]},
     {loadUnit_maskInput_lo[30095:30080]},
     {loadUnit_maskInput_lo[30079:30064]},
     {loadUnit_maskInput_lo[30063:30048]},
     {loadUnit_maskInput_lo[30047:30032]},
     {loadUnit_maskInput_lo[30031:30016]},
     {loadUnit_maskInput_lo[30015:30000]},
     {loadUnit_maskInput_lo[29999:29984]},
     {loadUnit_maskInput_lo[29983:29968]},
     {loadUnit_maskInput_lo[29967:29952]},
     {loadUnit_maskInput_lo[29951:29936]},
     {loadUnit_maskInput_lo[29935:29920]},
     {loadUnit_maskInput_lo[29919:29904]},
     {loadUnit_maskInput_lo[29903:29888]},
     {loadUnit_maskInput_lo[29887:29872]},
     {loadUnit_maskInput_lo[29871:29856]},
     {loadUnit_maskInput_lo[29855:29840]},
     {loadUnit_maskInput_lo[29839:29824]},
     {loadUnit_maskInput_lo[29823:29808]},
     {loadUnit_maskInput_lo[29807:29792]},
     {loadUnit_maskInput_lo[29791:29776]},
     {loadUnit_maskInput_lo[29775:29760]},
     {loadUnit_maskInput_lo[29759:29744]},
     {loadUnit_maskInput_lo[29743:29728]},
     {loadUnit_maskInput_lo[29727:29712]},
     {loadUnit_maskInput_lo[29711:29696]},
     {loadUnit_maskInput_lo[29695:29680]},
     {loadUnit_maskInput_lo[29679:29664]},
     {loadUnit_maskInput_lo[29663:29648]},
     {loadUnit_maskInput_lo[29647:29632]},
     {loadUnit_maskInput_lo[29631:29616]},
     {loadUnit_maskInput_lo[29615:29600]},
     {loadUnit_maskInput_lo[29599:29584]},
     {loadUnit_maskInput_lo[29583:29568]},
     {loadUnit_maskInput_lo[29567:29552]},
     {loadUnit_maskInput_lo[29551:29536]},
     {loadUnit_maskInput_lo[29535:29520]},
     {loadUnit_maskInput_lo[29519:29504]},
     {loadUnit_maskInput_lo[29503:29488]},
     {loadUnit_maskInput_lo[29487:29472]},
     {loadUnit_maskInput_lo[29471:29456]},
     {loadUnit_maskInput_lo[29455:29440]},
     {loadUnit_maskInput_lo[29439:29424]},
     {loadUnit_maskInput_lo[29423:29408]},
     {loadUnit_maskInput_lo[29407:29392]},
     {loadUnit_maskInput_lo[29391:29376]},
     {loadUnit_maskInput_lo[29375:29360]},
     {loadUnit_maskInput_lo[29359:29344]},
     {loadUnit_maskInput_lo[29343:29328]},
     {loadUnit_maskInput_lo[29327:29312]},
     {loadUnit_maskInput_lo[29311:29296]},
     {loadUnit_maskInput_lo[29295:29280]},
     {loadUnit_maskInput_lo[29279:29264]},
     {loadUnit_maskInput_lo[29263:29248]},
     {loadUnit_maskInput_lo[29247:29232]},
     {loadUnit_maskInput_lo[29231:29216]},
     {loadUnit_maskInput_lo[29215:29200]},
     {loadUnit_maskInput_lo[29199:29184]},
     {loadUnit_maskInput_lo[29183:29168]},
     {loadUnit_maskInput_lo[29167:29152]},
     {loadUnit_maskInput_lo[29151:29136]},
     {loadUnit_maskInput_lo[29135:29120]},
     {loadUnit_maskInput_lo[29119:29104]},
     {loadUnit_maskInput_lo[29103:29088]},
     {loadUnit_maskInput_lo[29087:29072]},
     {loadUnit_maskInput_lo[29071:29056]},
     {loadUnit_maskInput_lo[29055:29040]},
     {loadUnit_maskInput_lo[29039:29024]},
     {loadUnit_maskInput_lo[29023:29008]},
     {loadUnit_maskInput_lo[29007:28992]},
     {loadUnit_maskInput_lo[28991:28976]},
     {loadUnit_maskInput_lo[28975:28960]},
     {loadUnit_maskInput_lo[28959:28944]},
     {loadUnit_maskInput_lo[28943:28928]},
     {loadUnit_maskInput_lo[28927:28912]},
     {loadUnit_maskInput_lo[28911:28896]},
     {loadUnit_maskInput_lo[28895:28880]},
     {loadUnit_maskInput_lo[28879:28864]},
     {loadUnit_maskInput_lo[28863:28848]},
     {loadUnit_maskInput_lo[28847:28832]},
     {loadUnit_maskInput_lo[28831:28816]},
     {loadUnit_maskInput_lo[28815:28800]},
     {loadUnit_maskInput_lo[28799:28784]},
     {loadUnit_maskInput_lo[28783:28768]},
     {loadUnit_maskInput_lo[28767:28752]},
     {loadUnit_maskInput_lo[28751:28736]},
     {loadUnit_maskInput_lo[28735:28720]},
     {loadUnit_maskInput_lo[28719:28704]},
     {loadUnit_maskInput_lo[28703:28688]},
     {loadUnit_maskInput_lo[28687:28672]},
     {loadUnit_maskInput_lo[28671:28656]},
     {loadUnit_maskInput_lo[28655:28640]},
     {loadUnit_maskInput_lo[28639:28624]},
     {loadUnit_maskInput_lo[28623:28608]},
     {loadUnit_maskInput_lo[28607:28592]},
     {loadUnit_maskInput_lo[28591:28576]},
     {loadUnit_maskInput_lo[28575:28560]},
     {loadUnit_maskInput_lo[28559:28544]},
     {loadUnit_maskInput_lo[28543:28528]},
     {loadUnit_maskInput_lo[28527:28512]},
     {loadUnit_maskInput_lo[28511:28496]},
     {loadUnit_maskInput_lo[28495:28480]},
     {loadUnit_maskInput_lo[28479:28464]},
     {loadUnit_maskInput_lo[28463:28448]},
     {loadUnit_maskInput_lo[28447:28432]},
     {loadUnit_maskInput_lo[28431:28416]},
     {loadUnit_maskInput_lo[28415:28400]},
     {loadUnit_maskInput_lo[28399:28384]},
     {loadUnit_maskInput_lo[28383:28368]},
     {loadUnit_maskInput_lo[28367:28352]},
     {loadUnit_maskInput_lo[28351:28336]},
     {loadUnit_maskInput_lo[28335:28320]},
     {loadUnit_maskInput_lo[28319:28304]},
     {loadUnit_maskInput_lo[28303:28288]},
     {loadUnit_maskInput_lo[28287:28272]},
     {loadUnit_maskInput_lo[28271:28256]},
     {loadUnit_maskInput_lo[28255:28240]},
     {loadUnit_maskInput_lo[28239:28224]},
     {loadUnit_maskInput_lo[28223:28208]},
     {loadUnit_maskInput_lo[28207:28192]},
     {loadUnit_maskInput_lo[28191:28176]},
     {loadUnit_maskInput_lo[28175:28160]},
     {loadUnit_maskInput_lo[28159:28144]},
     {loadUnit_maskInput_lo[28143:28128]},
     {loadUnit_maskInput_lo[28127:28112]},
     {loadUnit_maskInput_lo[28111:28096]},
     {loadUnit_maskInput_lo[28095:28080]},
     {loadUnit_maskInput_lo[28079:28064]},
     {loadUnit_maskInput_lo[28063:28048]},
     {loadUnit_maskInput_lo[28047:28032]},
     {loadUnit_maskInput_lo[28031:28016]},
     {loadUnit_maskInput_lo[28015:28000]},
     {loadUnit_maskInput_lo[27999:27984]},
     {loadUnit_maskInput_lo[27983:27968]},
     {loadUnit_maskInput_lo[27967:27952]},
     {loadUnit_maskInput_lo[27951:27936]},
     {loadUnit_maskInput_lo[27935:27920]},
     {loadUnit_maskInput_lo[27919:27904]},
     {loadUnit_maskInput_lo[27903:27888]},
     {loadUnit_maskInput_lo[27887:27872]},
     {loadUnit_maskInput_lo[27871:27856]},
     {loadUnit_maskInput_lo[27855:27840]},
     {loadUnit_maskInput_lo[27839:27824]},
     {loadUnit_maskInput_lo[27823:27808]},
     {loadUnit_maskInput_lo[27807:27792]},
     {loadUnit_maskInput_lo[27791:27776]},
     {loadUnit_maskInput_lo[27775:27760]},
     {loadUnit_maskInput_lo[27759:27744]},
     {loadUnit_maskInput_lo[27743:27728]},
     {loadUnit_maskInput_lo[27727:27712]},
     {loadUnit_maskInput_lo[27711:27696]},
     {loadUnit_maskInput_lo[27695:27680]},
     {loadUnit_maskInput_lo[27679:27664]},
     {loadUnit_maskInput_lo[27663:27648]},
     {loadUnit_maskInput_lo[27647:27632]},
     {loadUnit_maskInput_lo[27631:27616]},
     {loadUnit_maskInput_lo[27615:27600]},
     {loadUnit_maskInput_lo[27599:27584]},
     {loadUnit_maskInput_lo[27583:27568]},
     {loadUnit_maskInput_lo[27567:27552]},
     {loadUnit_maskInput_lo[27551:27536]},
     {loadUnit_maskInput_lo[27535:27520]},
     {loadUnit_maskInput_lo[27519:27504]},
     {loadUnit_maskInput_lo[27503:27488]},
     {loadUnit_maskInput_lo[27487:27472]},
     {loadUnit_maskInput_lo[27471:27456]},
     {loadUnit_maskInput_lo[27455:27440]},
     {loadUnit_maskInput_lo[27439:27424]},
     {loadUnit_maskInput_lo[27423:27408]},
     {loadUnit_maskInput_lo[27407:27392]},
     {loadUnit_maskInput_lo[27391:27376]},
     {loadUnit_maskInput_lo[27375:27360]},
     {loadUnit_maskInput_lo[27359:27344]},
     {loadUnit_maskInput_lo[27343:27328]},
     {loadUnit_maskInput_lo[27327:27312]},
     {loadUnit_maskInput_lo[27311:27296]},
     {loadUnit_maskInput_lo[27295:27280]},
     {loadUnit_maskInput_lo[27279:27264]},
     {loadUnit_maskInput_lo[27263:27248]},
     {loadUnit_maskInput_lo[27247:27232]},
     {loadUnit_maskInput_lo[27231:27216]},
     {loadUnit_maskInput_lo[27215:27200]},
     {loadUnit_maskInput_lo[27199:27184]},
     {loadUnit_maskInput_lo[27183:27168]},
     {loadUnit_maskInput_lo[27167:27152]},
     {loadUnit_maskInput_lo[27151:27136]},
     {loadUnit_maskInput_lo[27135:27120]},
     {loadUnit_maskInput_lo[27119:27104]},
     {loadUnit_maskInput_lo[27103:27088]},
     {loadUnit_maskInput_lo[27087:27072]},
     {loadUnit_maskInput_lo[27071:27056]},
     {loadUnit_maskInput_lo[27055:27040]},
     {loadUnit_maskInput_lo[27039:27024]},
     {loadUnit_maskInput_lo[27023:27008]},
     {loadUnit_maskInput_lo[27007:26992]},
     {loadUnit_maskInput_lo[26991:26976]},
     {loadUnit_maskInput_lo[26975:26960]},
     {loadUnit_maskInput_lo[26959:26944]},
     {loadUnit_maskInput_lo[26943:26928]},
     {loadUnit_maskInput_lo[26927:26912]},
     {loadUnit_maskInput_lo[26911:26896]},
     {loadUnit_maskInput_lo[26895:26880]},
     {loadUnit_maskInput_lo[26879:26864]},
     {loadUnit_maskInput_lo[26863:26848]},
     {loadUnit_maskInput_lo[26847:26832]},
     {loadUnit_maskInput_lo[26831:26816]},
     {loadUnit_maskInput_lo[26815:26800]},
     {loadUnit_maskInput_lo[26799:26784]},
     {loadUnit_maskInput_lo[26783:26768]},
     {loadUnit_maskInput_lo[26767:26752]},
     {loadUnit_maskInput_lo[26751:26736]},
     {loadUnit_maskInput_lo[26735:26720]},
     {loadUnit_maskInput_lo[26719:26704]},
     {loadUnit_maskInput_lo[26703:26688]},
     {loadUnit_maskInput_lo[26687:26672]},
     {loadUnit_maskInput_lo[26671:26656]},
     {loadUnit_maskInput_lo[26655:26640]},
     {loadUnit_maskInput_lo[26639:26624]},
     {loadUnit_maskInput_lo[26623:26608]},
     {loadUnit_maskInput_lo[26607:26592]},
     {loadUnit_maskInput_lo[26591:26576]},
     {loadUnit_maskInput_lo[26575:26560]},
     {loadUnit_maskInput_lo[26559:26544]},
     {loadUnit_maskInput_lo[26543:26528]},
     {loadUnit_maskInput_lo[26527:26512]},
     {loadUnit_maskInput_lo[26511:26496]},
     {loadUnit_maskInput_lo[26495:26480]},
     {loadUnit_maskInput_lo[26479:26464]},
     {loadUnit_maskInput_lo[26463:26448]},
     {loadUnit_maskInput_lo[26447:26432]},
     {loadUnit_maskInput_lo[26431:26416]},
     {loadUnit_maskInput_lo[26415:26400]},
     {loadUnit_maskInput_lo[26399:26384]},
     {loadUnit_maskInput_lo[26383:26368]},
     {loadUnit_maskInput_lo[26367:26352]},
     {loadUnit_maskInput_lo[26351:26336]},
     {loadUnit_maskInput_lo[26335:26320]},
     {loadUnit_maskInput_lo[26319:26304]},
     {loadUnit_maskInput_lo[26303:26288]},
     {loadUnit_maskInput_lo[26287:26272]},
     {loadUnit_maskInput_lo[26271:26256]},
     {loadUnit_maskInput_lo[26255:26240]},
     {loadUnit_maskInput_lo[26239:26224]},
     {loadUnit_maskInput_lo[26223:26208]},
     {loadUnit_maskInput_lo[26207:26192]},
     {loadUnit_maskInput_lo[26191:26176]},
     {loadUnit_maskInput_lo[26175:26160]},
     {loadUnit_maskInput_lo[26159:26144]},
     {loadUnit_maskInput_lo[26143:26128]},
     {loadUnit_maskInput_lo[26127:26112]},
     {loadUnit_maskInput_lo[26111:26096]},
     {loadUnit_maskInput_lo[26095:26080]},
     {loadUnit_maskInput_lo[26079:26064]},
     {loadUnit_maskInput_lo[26063:26048]},
     {loadUnit_maskInput_lo[26047:26032]},
     {loadUnit_maskInput_lo[26031:26016]},
     {loadUnit_maskInput_lo[26015:26000]},
     {loadUnit_maskInput_lo[25999:25984]},
     {loadUnit_maskInput_lo[25983:25968]},
     {loadUnit_maskInput_lo[25967:25952]},
     {loadUnit_maskInput_lo[25951:25936]},
     {loadUnit_maskInput_lo[25935:25920]},
     {loadUnit_maskInput_lo[25919:25904]},
     {loadUnit_maskInput_lo[25903:25888]},
     {loadUnit_maskInput_lo[25887:25872]},
     {loadUnit_maskInput_lo[25871:25856]},
     {loadUnit_maskInput_lo[25855:25840]},
     {loadUnit_maskInput_lo[25839:25824]},
     {loadUnit_maskInput_lo[25823:25808]},
     {loadUnit_maskInput_lo[25807:25792]},
     {loadUnit_maskInput_lo[25791:25776]},
     {loadUnit_maskInput_lo[25775:25760]},
     {loadUnit_maskInput_lo[25759:25744]},
     {loadUnit_maskInput_lo[25743:25728]},
     {loadUnit_maskInput_lo[25727:25712]},
     {loadUnit_maskInput_lo[25711:25696]},
     {loadUnit_maskInput_lo[25695:25680]},
     {loadUnit_maskInput_lo[25679:25664]},
     {loadUnit_maskInput_lo[25663:25648]},
     {loadUnit_maskInput_lo[25647:25632]},
     {loadUnit_maskInput_lo[25631:25616]},
     {loadUnit_maskInput_lo[25615:25600]},
     {loadUnit_maskInput_lo[25599:25584]},
     {loadUnit_maskInput_lo[25583:25568]},
     {loadUnit_maskInput_lo[25567:25552]},
     {loadUnit_maskInput_lo[25551:25536]},
     {loadUnit_maskInput_lo[25535:25520]},
     {loadUnit_maskInput_lo[25519:25504]},
     {loadUnit_maskInput_lo[25503:25488]},
     {loadUnit_maskInput_lo[25487:25472]},
     {loadUnit_maskInput_lo[25471:25456]},
     {loadUnit_maskInput_lo[25455:25440]},
     {loadUnit_maskInput_lo[25439:25424]},
     {loadUnit_maskInput_lo[25423:25408]},
     {loadUnit_maskInput_lo[25407:25392]},
     {loadUnit_maskInput_lo[25391:25376]},
     {loadUnit_maskInput_lo[25375:25360]},
     {loadUnit_maskInput_lo[25359:25344]},
     {loadUnit_maskInput_lo[25343:25328]},
     {loadUnit_maskInput_lo[25327:25312]},
     {loadUnit_maskInput_lo[25311:25296]},
     {loadUnit_maskInput_lo[25295:25280]},
     {loadUnit_maskInput_lo[25279:25264]},
     {loadUnit_maskInput_lo[25263:25248]},
     {loadUnit_maskInput_lo[25247:25232]},
     {loadUnit_maskInput_lo[25231:25216]},
     {loadUnit_maskInput_lo[25215:25200]},
     {loadUnit_maskInput_lo[25199:25184]},
     {loadUnit_maskInput_lo[25183:25168]},
     {loadUnit_maskInput_lo[25167:25152]},
     {loadUnit_maskInput_lo[25151:25136]},
     {loadUnit_maskInput_lo[25135:25120]},
     {loadUnit_maskInput_lo[25119:25104]},
     {loadUnit_maskInput_lo[25103:25088]},
     {loadUnit_maskInput_lo[25087:25072]},
     {loadUnit_maskInput_lo[25071:25056]},
     {loadUnit_maskInput_lo[25055:25040]},
     {loadUnit_maskInput_lo[25039:25024]},
     {loadUnit_maskInput_lo[25023:25008]},
     {loadUnit_maskInput_lo[25007:24992]},
     {loadUnit_maskInput_lo[24991:24976]},
     {loadUnit_maskInput_lo[24975:24960]},
     {loadUnit_maskInput_lo[24959:24944]},
     {loadUnit_maskInput_lo[24943:24928]},
     {loadUnit_maskInput_lo[24927:24912]},
     {loadUnit_maskInput_lo[24911:24896]},
     {loadUnit_maskInput_lo[24895:24880]},
     {loadUnit_maskInput_lo[24879:24864]},
     {loadUnit_maskInput_lo[24863:24848]},
     {loadUnit_maskInput_lo[24847:24832]},
     {loadUnit_maskInput_lo[24831:24816]},
     {loadUnit_maskInput_lo[24815:24800]},
     {loadUnit_maskInput_lo[24799:24784]},
     {loadUnit_maskInput_lo[24783:24768]},
     {loadUnit_maskInput_lo[24767:24752]},
     {loadUnit_maskInput_lo[24751:24736]},
     {loadUnit_maskInput_lo[24735:24720]},
     {loadUnit_maskInput_lo[24719:24704]},
     {loadUnit_maskInput_lo[24703:24688]},
     {loadUnit_maskInput_lo[24687:24672]},
     {loadUnit_maskInput_lo[24671:24656]},
     {loadUnit_maskInput_lo[24655:24640]},
     {loadUnit_maskInput_lo[24639:24624]},
     {loadUnit_maskInput_lo[24623:24608]},
     {loadUnit_maskInput_lo[24607:24592]},
     {loadUnit_maskInput_lo[24591:24576]},
     {loadUnit_maskInput_lo[24575:24560]},
     {loadUnit_maskInput_lo[24559:24544]},
     {loadUnit_maskInput_lo[24543:24528]},
     {loadUnit_maskInput_lo[24527:24512]},
     {loadUnit_maskInput_lo[24511:24496]},
     {loadUnit_maskInput_lo[24495:24480]},
     {loadUnit_maskInput_lo[24479:24464]},
     {loadUnit_maskInput_lo[24463:24448]},
     {loadUnit_maskInput_lo[24447:24432]},
     {loadUnit_maskInput_lo[24431:24416]},
     {loadUnit_maskInput_lo[24415:24400]},
     {loadUnit_maskInput_lo[24399:24384]},
     {loadUnit_maskInput_lo[24383:24368]},
     {loadUnit_maskInput_lo[24367:24352]},
     {loadUnit_maskInput_lo[24351:24336]},
     {loadUnit_maskInput_lo[24335:24320]},
     {loadUnit_maskInput_lo[24319:24304]},
     {loadUnit_maskInput_lo[24303:24288]},
     {loadUnit_maskInput_lo[24287:24272]},
     {loadUnit_maskInput_lo[24271:24256]},
     {loadUnit_maskInput_lo[24255:24240]},
     {loadUnit_maskInput_lo[24239:24224]},
     {loadUnit_maskInput_lo[24223:24208]},
     {loadUnit_maskInput_lo[24207:24192]},
     {loadUnit_maskInput_lo[24191:24176]},
     {loadUnit_maskInput_lo[24175:24160]},
     {loadUnit_maskInput_lo[24159:24144]},
     {loadUnit_maskInput_lo[24143:24128]},
     {loadUnit_maskInput_lo[24127:24112]},
     {loadUnit_maskInput_lo[24111:24096]},
     {loadUnit_maskInput_lo[24095:24080]},
     {loadUnit_maskInput_lo[24079:24064]},
     {loadUnit_maskInput_lo[24063:24048]},
     {loadUnit_maskInput_lo[24047:24032]},
     {loadUnit_maskInput_lo[24031:24016]},
     {loadUnit_maskInput_lo[24015:24000]},
     {loadUnit_maskInput_lo[23999:23984]},
     {loadUnit_maskInput_lo[23983:23968]},
     {loadUnit_maskInput_lo[23967:23952]},
     {loadUnit_maskInput_lo[23951:23936]},
     {loadUnit_maskInput_lo[23935:23920]},
     {loadUnit_maskInput_lo[23919:23904]},
     {loadUnit_maskInput_lo[23903:23888]},
     {loadUnit_maskInput_lo[23887:23872]},
     {loadUnit_maskInput_lo[23871:23856]},
     {loadUnit_maskInput_lo[23855:23840]},
     {loadUnit_maskInput_lo[23839:23824]},
     {loadUnit_maskInput_lo[23823:23808]},
     {loadUnit_maskInput_lo[23807:23792]},
     {loadUnit_maskInput_lo[23791:23776]},
     {loadUnit_maskInput_lo[23775:23760]},
     {loadUnit_maskInput_lo[23759:23744]},
     {loadUnit_maskInput_lo[23743:23728]},
     {loadUnit_maskInput_lo[23727:23712]},
     {loadUnit_maskInput_lo[23711:23696]},
     {loadUnit_maskInput_lo[23695:23680]},
     {loadUnit_maskInput_lo[23679:23664]},
     {loadUnit_maskInput_lo[23663:23648]},
     {loadUnit_maskInput_lo[23647:23632]},
     {loadUnit_maskInput_lo[23631:23616]},
     {loadUnit_maskInput_lo[23615:23600]},
     {loadUnit_maskInput_lo[23599:23584]},
     {loadUnit_maskInput_lo[23583:23568]},
     {loadUnit_maskInput_lo[23567:23552]},
     {loadUnit_maskInput_lo[23551:23536]},
     {loadUnit_maskInput_lo[23535:23520]},
     {loadUnit_maskInput_lo[23519:23504]},
     {loadUnit_maskInput_lo[23503:23488]},
     {loadUnit_maskInput_lo[23487:23472]},
     {loadUnit_maskInput_lo[23471:23456]},
     {loadUnit_maskInput_lo[23455:23440]},
     {loadUnit_maskInput_lo[23439:23424]},
     {loadUnit_maskInput_lo[23423:23408]},
     {loadUnit_maskInput_lo[23407:23392]},
     {loadUnit_maskInput_lo[23391:23376]},
     {loadUnit_maskInput_lo[23375:23360]},
     {loadUnit_maskInput_lo[23359:23344]},
     {loadUnit_maskInput_lo[23343:23328]},
     {loadUnit_maskInput_lo[23327:23312]},
     {loadUnit_maskInput_lo[23311:23296]},
     {loadUnit_maskInput_lo[23295:23280]},
     {loadUnit_maskInput_lo[23279:23264]},
     {loadUnit_maskInput_lo[23263:23248]},
     {loadUnit_maskInput_lo[23247:23232]},
     {loadUnit_maskInput_lo[23231:23216]},
     {loadUnit_maskInput_lo[23215:23200]},
     {loadUnit_maskInput_lo[23199:23184]},
     {loadUnit_maskInput_lo[23183:23168]},
     {loadUnit_maskInput_lo[23167:23152]},
     {loadUnit_maskInput_lo[23151:23136]},
     {loadUnit_maskInput_lo[23135:23120]},
     {loadUnit_maskInput_lo[23119:23104]},
     {loadUnit_maskInput_lo[23103:23088]},
     {loadUnit_maskInput_lo[23087:23072]},
     {loadUnit_maskInput_lo[23071:23056]},
     {loadUnit_maskInput_lo[23055:23040]},
     {loadUnit_maskInput_lo[23039:23024]},
     {loadUnit_maskInput_lo[23023:23008]},
     {loadUnit_maskInput_lo[23007:22992]},
     {loadUnit_maskInput_lo[22991:22976]},
     {loadUnit_maskInput_lo[22975:22960]},
     {loadUnit_maskInput_lo[22959:22944]},
     {loadUnit_maskInput_lo[22943:22928]},
     {loadUnit_maskInput_lo[22927:22912]},
     {loadUnit_maskInput_lo[22911:22896]},
     {loadUnit_maskInput_lo[22895:22880]},
     {loadUnit_maskInput_lo[22879:22864]},
     {loadUnit_maskInput_lo[22863:22848]},
     {loadUnit_maskInput_lo[22847:22832]},
     {loadUnit_maskInput_lo[22831:22816]},
     {loadUnit_maskInput_lo[22815:22800]},
     {loadUnit_maskInput_lo[22799:22784]},
     {loadUnit_maskInput_lo[22783:22768]},
     {loadUnit_maskInput_lo[22767:22752]},
     {loadUnit_maskInput_lo[22751:22736]},
     {loadUnit_maskInput_lo[22735:22720]},
     {loadUnit_maskInput_lo[22719:22704]},
     {loadUnit_maskInput_lo[22703:22688]},
     {loadUnit_maskInput_lo[22687:22672]},
     {loadUnit_maskInput_lo[22671:22656]},
     {loadUnit_maskInput_lo[22655:22640]},
     {loadUnit_maskInput_lo[22639:22624]},
     {loadUnit_maskInput_lo[22623:22608]},
     {loadUnit_maskInput_lo[22607:22592]},
     {loadUnit_maskInput_lo[22591:22576]},
     {loadUnit_maskInput_lo[22575:22560]},
     {loadUnit_maskInput_lo[22559:22544]},
     {loadUnit_maskInput_lo[22543:22528]},
     {loadUnit_maskInput_lo[22527:22512]},
     {loadUnit_maskInput_lo[22511:22496]},
     {loadUnit_maskInput_lo[22495:22480]},
     {loadUnit_maskInput_lo[22479:22464]},
     {loadUnit_maskInput_lo[22463:22448]},
     {loadUnit_maskInput_lo[22447:22432]},
     {loadUnit_maskInput_lo[22431:22416]},
     {loadUnit_maskInput_lo[22415:22400]},
     {loadUnit_maskInput_lo[22399:22384]},
     {loadUnit_maskInput_lo[22383:22368]},
     {loadUnit_maskInput_lo[22367:22352]},
     {loadUnit_maskInput_lo[22351:22336]},
     {loadUnit_maskInput_lo[22335:22320]},
     {loadUnit_maskInput_lo[22319:22304]},
     {loadUnit_maskInput_lo[22303:22288]},
     {loadUnit_maskInput_lo[22287:22272]},
     {loadUnit_maskInput_lo[22271:22256]},
     {loadUnit_maskInput_lo[22255:22240]},
     {loadUnit_maskInput_lo[22239:22224]},
     {loadUnit_maskInput_lo[22223:22208]},
     {loadUnit_maskInput_lo[22207:22192]},
     {loadUnit_maskInput_lo[22191:22176]},
     {loadUnit_maskInput_lo[22175:22160]},
     {loadUnit_maskInput_lo[22159:22144]},
     {loadUnit_maskInput_lo[22143:22128]},
     {loadUnit_maskInput_lo[22127:22112]},
     {loadUnit_maskInput_lo[22111:22096]},
     {loadUnit_maskInput_lo[22095:22080]},
     {loadUnit_maskInput_lo[22079:22064]},
     {loadUnit_maskInput_lo[22063:22048]},
     {loadUnit_maskInput_lo[22047:22032]},
     {loadUnit_maskInput_lo[22031:22016]},
     {loadUnit_maskInput_lo[22015:22000]},
     {loadUnit_maskInput_lo[21999:21984]},
     {loadUnit_maskInput_lo[21983:21968]},
     {loadUnit_maskInput_lo[21967:21952]},
     {loadUnit_maskInput_lo[21951:21936]},
     {loadUnit_maskInput_lo[21935:21920]},
     {loadUnit_maskInput_lo[21919:21904]},
     {loadUnit_maskInput_lo[21903:21888]},
     {loadUnit_maskInput_lo[21887:21872]},
     {loadUnit_maskInput_lo[21871:21856]},
     {loadUnit_maskInput_lo[21855:21840]},
     {loadUnit_maskInput_lo[21839:21824]},
     {loadUnit_maskInput_lo[21823:21808]},
     {loadUnit_maskInput_lo[21807:21792]},
     {loadUnit_maskInput_lo[21791:21776]},
     {loadUnit_maskInput_lo[21775:21760]},
     {loadUnit_maskInput_lo[21759:21744]},
     {loadUnit_maskInput_lo[21743:21728]},
     {loadUnit_maskInput_lo[21727:21712]},
     {loadUnit_maskInput_lo[21711:21696]},
     {loadUnit_maskInput_lo[21695:21680]},
     {loadUnit_maskInput_lo[21679:21664]},
     {loadUnit_maskInput_lo[21663:21648]},
     {loadUnit_maskInput_lo[21647:21632]},
     {loadUnit_maskInput_lo[21631:21616]},
     {loadUnit_maskInput_lo[21615:21600]},
     {loadUnit_maskInput_lo[21599:21584]},
     {loadUnit_maskInput_lo[21583:21568]},
     {loadUnit_maskInput_lo[21567:21552]},
     {loadUnit_maskInput_lo[21551:21536]},
     {loadUnit_maskInput_lo[21535:21520]},
     {loadUnit_maskInput_lo[21519:21504]},
     {loadUnit_maskInput_lo[21503:21488]},
     {loadUnit_maskInput_lo[21487:21472]},
     {loadUnit_maskInput_lo[21471:21456]},
     {loadUnit_maskInput_lo[21455:21440]},
     {loadUnit_maskInput_lo[21439:21424]},
     {loadUnit_maskInput_lo[21423:21408]},
     {loadUnit_maskInput_lo[21407:21392]},
     {loadUnit_maskInput_lo[21391:21376]},
     {loadUnit_maskInput_lo[21375:21360]},
     {loadUnit_maskInput_lo[21359:21344]},
     {loadUnit_maskInput_lo[21343:21328]},
     {loadUnit_maskInput_lo[21327:21312]},
     {loadUnit_maskInput_lo[21311:21296]},
     {loadUnit_maskInput_lo[21295:21280]},
     {loadUnit_maskInput_lo[21279:21264]},
     {loadUnit_maskInput_lo[21263:21248]},
     {loadUnit_maskInput_lo[21247:21232]},
     {loadUnit_maskInput_lo[21231:21216]},
     {loadUnit_maskInput_lo[21215:21200]},
     {loadUnit_maskInput_lo[21199:21184]},
     {loadUnit_maskInput_lo[21183:21168]},
     {loadUnit_maskInput_lo[21167:21152]},
     {loadUnit_maskInput_lo[21151:21136]},
     {loadUnit_maskInput_lo[21135:21120]},
     {loadUnit_maskInput_lo[21119:21104]},
     {loadUnit_maskInput_lo[21103:21088]},
     {loadUnit_maskInput_lo[21087:21072]},
     {loadUnit_maskInput_lo[21071:21056]},
     {loadUnit_maskInput_lo[21055:21040]},
     {loadUnit_maskInput_lo[21039:21024]},
     {loadUnit_maskInput_lo[21023:21008]},
     {loadUnit_maskInput_lo[21007:20992]},
     {loadUnit_maskInput_lo[20991:20976]},
     {loadUnit_maskInput_lo[20975:20960]},
     {loadUnit_maskInput_lo[20959:20944]},
     {loadUnit_maskInput_lo[20943:20928]},
     {loadUnit_maskInput_lo[20927:20912]},
     {loadUnit_maskInput_lo[20911:20896]},
     {loadUnit_maskInput_lo[20895:20880]},
     {loadUnit_maskInput_lo[20879:20864]},
     {loadUnit_maskInput_lo[20863:20848]},
     {loadUnit_maskInput_lo[20847:20832]},
     {loadUnit_maskInput_lo[20831:20816]},
     {loadUnit_maskInput_lo[20815:20800]},
     {loadUnit_maskInput_lo[20799:20784]},
     {loadUnit_maskInput_lo[20783:20768]},
     {loadUnit_maskInput_lo[20767:20752]},
     {loadUnit_maskInput_lo[20751:20736]},
     {loadUnit_maskInput_lo[20735:20720]},
     {loadUnit_maskInput_lo[20719:20704]},
     {loadUnit_maskInput_lo[20703:20688]},
     {loadUnit_maskInput_lo[20687:20672]},
     {loadUnit_maskInput_lo[20671:20656]},
     {loadUnit_maskInput_lo[20655:20640]},
     {loadUnit_maskInput_lo[20639:20624]},
     {loadUnit_maskInput_lo[20623:20608]},
     {loadUnit_maskInput_lo[20607:20592]},
     {loadUnit_maskInput_lo[20591:20576]},
     {loadUnit_maskInput_lo[20575:20560]},
     {loadUnit_maskInput_lo[20559:20544]},
     {loadUnit_maskInput_lo[20543:20528]},
     {loadUnit_maskInput_lo[20527:20512]},
     {loadUnit_maskInput_lo[20511:20496]},
     {loadUnit_maskInput_lo[20495:20480]},
     {loadUnit_maskInput_lo[20479:20464]},
     {loadUnit_maskInput_lo[20463:20448]},
     {loadUnit_maskInput_lo[20447:20432]},
     {loadUnit_maskInput_lo[20431:20416]},
     {loadUnit_maskInput_lo[20415:20400]},
     {loadUnit_maskInput_lo[20399:20384]},
     {loadUnit_maskInput_lo[20383:20368]},
     {loadUnit_maskInput_lo[20367:20352]},
     {loadUnit_maskInput_lo[20351:20336]},
     {loadUnit_maskInput_lo[20335:20320]},
     {loadUnit_maskInput_lo[20319:20304]},
     {loadUnit_maskInput_lo[20303:20288]},
     {loadUnit_maskInput_lo[20287:20272]},
     {loadUnit_maskInput_lo[20271:20256]},
     {loadUnit_maskInput_lo[20255:20240]},
     {loadUnit_maskInput_lo[20239:20224]},
     {loadUnit_maskInput_lo[20223:20208]},
     {loadUnit_maskInput_lo[20207:20192]},
     {loadUnit_maskInput_lo[20191:20176]},
     {loadUnit_maskInput_lo[20175:20160]},
     {loadUnit_maskInput_lo[20159:20144]},
     {loadUnit_maskInput_lo[20143:20128]},
     {loadUnit_maskInput_lo[20127:20112]},
     {loadUnit_maskInput_lo[20111:20096]},
     {loadUnit_maskInput_lo[20095:20080]},
     {loadUnit_maskInput_lo[20079:20064]},
     {loadUnit_maskInput_lo[20063:20048]},
     {loadUnit_maskInput_lo[20047:20032]},
     {loadUnit_maskInput_lo[20031:20016]},
     {loadUnit_maskInput_lo[20015:20000]},
     {loadUnit_maskInput_lo[19999:19984]},
     {loadUnit_maskInput_lo[19983:19968]},
     {loadUnit_maskInput_lo[19967:19952]},
     {loadUnit_maskInput_lo[19951:19936]},
     {loadUnit_maskInput_lo[19935:19920]},
     {loadUnit_maskInput_lo[19919:19904]},
     {loadUnit_maskInput_lo[19903:19888]},
     {loadUnit_maskInput_lo[19887:19872]},
     {loadUnit_maskInput_lo[19871:19856]},
     {loadUnit_maskInput_lo[19855:19840]},
     {loadUnit_maskInput_lo[19839:19824]},
     {loadUnit_maskInput_lo[19823:19808]},
     {loadUnit_maskInput_lo[19807:19792]},
     {loadUnit_maskInput_lo[19791:19776]},
     {loadUnit_maskInput_lo[19775:19760]},
     {loadUnit_maskInput_lo[19759:19744]},
     {loadUnit_maskInput_lo[19743:19728]},
     {loadUnit_maskInput_lo[19727:19712]},
     {loadUnit_maskInput_lo[19711:19696]},
     {loadUnit_maskInput_lo[19695:19680]},
     {loadUnit_maskInput_lo[19679:19664]},
     {loadUnit_maskInput_lo[19663:19648]},
     {loadUnit_maskInput_lo[19647:19632]},
     {loadUnit_maskInput_lo[19631:19616]},
     {loadUnit_maskInput_lo[19615:19600]},
     {loadUnit_maskInput_lo[19599:19584]},
     {loadUnit_maskInput_lo[19583:19568]},
     {loadUnit_maskInput_lo[19567:19552]},
     {loadUnit_maskInput_lo[19551:19536]},
     {loadUnit_maskInput_lo[19535:19520]},
     {loadUnit_maskInput_lo[19519:19504]},
     {loadUnit_maskInput_lo[19503:19488]},
     {loadUnit_maskInput_lo[19487:19472]},
     {loadUnit_maskInput_lo[19471:19456]},
     {loadUnit_maskInput_lo[19455:19440]},
     {loadUnit_maskInput_lo[19439:19424]},
     {loadUnit_maskInput_lo[19423:19408]},
     {loadUnit_maskInput_lo[19407:19392]},
     {loadUnit_maskInput_lo[19391:19376]},
     {loadUnit_maskInput_lo[19375:19360]},
     {loadUnit_maskInput_lo[19359:19344]},
     {loadUnit_maskInput_lo[19343:19328]},
     {loadUnit_maskInput_lo[19327:19312]},
     {loadUnit_maskInput_lo[19311:19296]},
     {loadUnit_maskInput_lo[19295:19280]},
     {loadUnit_maskInput_lo[19279:19264]},
     {loadUnit_maskInput_lo[19263:19248]},
     {loadUnit_maskInput_lo[19247:19232]},
     {loadUnit_maskInput_lo[19231:19216]},
     {loadUnit_maskInput_lo[19215:19200]},
     {loadUnit_maskInput_lo[19199:19184]},
     {loadUnit_maskInput_lo[19183:19168]},
     {loadUnit_maskInput_lo[19167:19152]},
     {loadUnit_maskInput_lo[19151:19136]},
     {loadUnit_maskInput_lo[19135:19120]},
     {loadUnit_maskInput_lo[19119:19104]},
     {loadUnit_maskInput_lo[19103:19088]},
     {loadUnit_maskInput_lo[19087:19072]},
     {loadUnit_maskInput_lo[19071:19056]},
     {loadUnit_maskInput_lo[19055:19040]},
     {loadUnit_maskInput_lo[19039:19024]},
     {loadUnit_maskInput_lo[19023:19008]},
     {loadUnit_maskInput_lo[19007:18992]},
     {loadUnit_maskInput_lo[18991:18976]},
     {loadUnit_maskInput_lo[18975:18960]},
     {loadUnit_maskInput_lo[18959:18944]},
     {loadUnit_maskInput_lo[18943:18928]},
     {loadUnit_maskInput_lo[18927:18912]},
     {loadUnit_maskInput_lo[18911:18896]},
     {loadUnit_maskInput_lo[18895:18880]},
     {loadUnit_maskInput_lo[18879:18864]},
     {loadUnit_maskInput_lo[18863:18848]},
     {loadUnit_maskInput_lo[18847:18832]},
     {loadUnit_maskInput_lo[18831:18816]},
     {loadUnit_maskInput_lo[18815:18800]},
     {loadUnit_maskInput_lo[18799:18784]},
     {loadUnit_maskInput_lo[18783:18768]},
     {loadUnit_maskInput_lo[18767:18752]},
     {loadUnit_maskInput_lo[18751:18736]},
     {loadUnit_maskInput_lo[18735:18720]},
     {loadUnit_maskInput_lo[18719:18704]},
     {loadUnit_maskInput_lo[18703:18688]},
     {loadUnit_maskInput_lo[18687:18672]},
     {loadUnit_maskInput_lo[18671:18656]},
     {loadUnit_maskInput_lo[18655:18640]},
     {loadUnit_maskInput_lo[18639:18624]},
     {loadUnit_maskInput_lo[18623:18608]},
     {loadUnit_maskInput_lo[18607:18592]},
     {loadUnit_maskInput_lo[18591:18576]},
     {loadUnit_maskInput_lo[18575:18560]},
     {loadUnit_maskInput_lo[18559:18544]},
     {loadUnit_maskInput_lo[18543:18528]},
     {loadUnit_maskInput_lo[18527:18512]},
     {loadUnit_maskInput_lo[18511:18496]},
     {loadUnit_maskInput_lo[18495:18480]},
     {loadUnit_maskInput_lo[18479:18464]},
     {loadUnit_maskInput_lo[18463:18448]},
     {loadUnit_maskInput_lo[18447:18432]},
     {loadUnit_maskInput_lo[18431:18416]},
     {loadUnit_maskInput_lo[18415:18400]},
     {loadUnit_maskInput_lo[18399:18384]},
     {loadUnit_maskInput_lo[18383:18368]},
     {loadUnit_maskInput_lo[18367:18352]},
     {loadUnit_maskInput_lo[18351:18336]},
     {loadUnit_maskInput_lo[18335:18320]},
     {loadUnit_maskInput_lo[18319:18304]},
     {loadUnit_maskInput_lo[18303:18288]},
     {loadUnit_maskInput_lo[18287:18272]},
     {loadUnit_maskInput_lo[18271:18256]},
     {loadUnit_maskInput_lo[18255:18240]},
     {loadUnit_maskInput_lo[18239:18224]},
     {loadUnit_maskInput_lo[18223:18208]},
     {loadUnit_maskInput_lo[18207:18192]},
     {loadUnit_maskInput_lo[18191:18176]},
     {loadUnit_maskInput_lo[18175:18160]},
     {loadUnit_maskInput_lo[18159:18144]},
     {loadUnit_maskInput_lo[18143:18128]},
     {loadUnit_maskInput_lo[18127:18112]},
     {loadUnit_maskInput_lo[18111:18096]},
     {loadUnit_maskInput_lo[18095:18080]},
     {loadUnit_maskInput_lo[18079:18064]},
     {loadUnit_maskInput_lo[18063:18048]},
     {loadUnit_maskInput_lo[18047:18032]},
     {loadUnit_maskInput_lo[18031:18016]},
     {loadUnit_maskInput_lo[18015:18000]},
     {loadUnit_maskInput_lo[17999:17984]},
     {loadUnit_maskInput_lo[17983:17968]},
     {loadUnit_maskInput_lo[17967:17952]},
     {loadUnit_maskInput_lo[17951:17936]},
     {loadUnit_maskInput_lo[17935:17920]},
     {loadUnit_maskInput_lo[17919:17904]},
     {loadUnit_maskInput_lo[17903:17888]},
     {loadUnit_maskInput_lo[17887:17872]},
     {loadUnit_maskInput_lo[17871:17856]},
     {loadUnit_maskInput_lo[17855:17840]},
     {loadUnit_maskInput_lo[17839:17824]},
     {loadUnit_maskInput_lo[17823:17808]},
     {loadUnit_maskInput_lo[17807:17792]},
     {loadUnit_maskInput_lo[17791:17776]},
     {loadUnit_maskInput_lo[17775:17760]},
     {loadUnit_maskInput_lo[17759:17744]},
     {loadUnit_maskInput_lo[17743:17728]},
     {loadUnit_maskInput_lo[17727:17712]},
     {loadUnit_maskInput_lo[17711:17696]},
     {loadUnit_maskInput_lo[17695:17680]},
     {loadUnit_maskInput_lo[17679:17664]},
     {loadUnit_maskInput_lo[17663:17648]},
     {loadUnit_maskInput_lo[17647:17632]},
     {loadUnit_maskInput_lo[17631:17616]},
     {loadUnit_maskInput_lo[17615:17600]},
     {loadUnit_maskInput_lo[17599:17584]},
     {loadUnit_maskInput_lo[17583:17568]},
     {loadUnit_maskInput_lo[17567:17552]},
     {loadUnit_maskInput_lo[17551:17536]},
     {loadUnit_maskInput_lo[17535:17520]},
     {loadUnit_maskInput_lo[17519:17504]},
     {loadUnit_maskInput_lo[17503:17488]},
     {loadUnit_maskInput_lo[17487:17472]},
     {loadUnit_maskInput_lo[17471:17456]},
     {loadUnit_maskInput_lo[17455:17440]},
     {loadUnit_maskInput_lo[17439:17424]},
     {loadUnit_maskInput_lo[17423:17408]},
     {loadUnit_maskInput_lo[17407:17392]},
     {loadUnit_maskInput_lo[17391:17376]},
     {loadUnit_maskInput_lo[17375:17360]},
     {loadUnit_maskInput_lo[17359:17344]},
     {loadUnit_maskInput_lo[17343:17328]},
     {loadUnit_maskInput_lo[17327:17312]},
     {loadUnit_maskInput_lo[17311:17296]},
     {loadUnit_maskInput_lo[17295:17280]},
     {loadUnit_maskInput_lo[17279:17264]},
     {loadUnit_maskInput_lo[17263:17248]},
     {loadUnit_maskInput_lo[17247:17232]},
     {loadUnit_maskInput_lo[17231:17216]},
     {loadUnit_maskInput_lo[17215:17200]},
     {loadUnit_maskInput_lo[17199:17184]},
     {loadUnit_maskInput_lo[17183:17168]},
     {loadUnit_maskInput_lo[17167:17152]},
     {loadUnit_maskInput_lo[17151:17136]},
     {loadUnit_maskInput_lo[17135:17120]},
     {loadUnit_maskInput_lo[17119:17104]},
     {loadUnit_maskInput_lo[17103:17088]},
     {loadUnit_maskInput_lo[17087:17072]},
     {loadUnit_maskInput_lo[17071:17056]},
     {loadUnit_maskInput_lo[17055:17040]},
     {loadUnit_maskInput_lo[17039:17024]},
     {loadUnit_maskInput_lo[17023:17008]},
     {loadUnit_maskInput_lo[17007:16992]},
     {loadUnit_maskInput_lo[16991:16976]},
     {loadUnit_maskInput_lo[16975:16960]},
     {loadUnit_maskInput_lo[16959:16944]},
     {loadUnit_maskInput_lo[16943:16928]},
     {loadUnit_maskInput_lo[16927:16912]},
     {loadUnit_maskInput_lo[16911:16896]},
     {loadUnit_maskInput_lo[16895:16880]},
     {loadUnit_maskInput_lo[16879:16864]},
     {loadUnit_maskInput_lo[16863:16848]},
     {loadUnit_maskInput_lo[16847:16832]},
     {loadUnit_maskInput_lo[16831:16816]},
     {loadUnit_maskInput_lo[16815:16800]},
     {loadUnit_maskInput_lo[16799:16784]},
     {loadUnit_maskInput_lo[16783:16768]},
     {loadUnit_maskInput_lo[16767:16752]},
     {loadUnit_maskInput_lo[16751:16736]},
     {loadUnit_maskInput_lo[16735:16720]},
     {loadUnit_maskInput_lo[16719:16704]},
     {loadUnit_maskInput_lo[16703:16688]},
     {loadUnit_maskInput_lo[16687:16672]},
     {loadUnit_maskInput_lo[16671:16656]},
     {loadUnit_maskInput_lo[16655:16640]},
     {loadUnit_maskInput_lo[16639:16624]},
     {loadUnit_maskInput_lo[16623:16608]},
     {loadUnit_maskInput_lo[16607:16592]},
     {loadUnit_maskInput_lo[16591:16576]},
     {loadUnit_maskInput_lo[16575:16560]},
     {loadUnit_maskInput_lo[16559:16544]},
     {loadUnit_maskInput_lo[16543:16528]},
     {loadUnit_maskInput_lo[16527:16512]},
     {loadUnit_maskInput_lo[16511:16496]},
     {loadUnit_maskInput_lo[16495:16480]},
     {loadUnit_maskInput_lo[16479:16464]},
     {loadUnit_maskInput_lo[16463:16448]},
     {loadUnit_maskInput_lo[16447:16432]},
     {loadUnit_maskInput_lo[16431:16416]},
     {loadUnit_maskInput_lo[16415:16400]},
     {loadUnit_maskInput_lo[16399:16384]},
     {loadUnit_maskInput_lo[16383:16368]},
     {loadUnit_maskInput_lo[16367:16352]},
     {loadUnit_maskInput_lo[16351:16336]},
     {loadUnit_maskInput_lo[16335:16320]},
     {loadUnit_maskInput_lo[16319:16304]},
     {loadUnit_maskInput_lo[16303:16288]},
     {loadUnit_maskInput_lo[16287:16272]},
     {loadUnit_maskInput_lo[16271:16256]},
     {loadUnit_maskInput_lo[16255:16240]},
     {loadUnit_maskInput_lo[16239:16224]},
     {loadUnit_maskInput_lo[16223:16208]},
     {loadUnit_maskInput_lo[16207:16192]},
     {loadUnit_maskInput_lo[16191:16176]},
     {loadUnit_maskInput_lo[16175:16160]},
     {loadUnit_maskInput_lo[16159:16144]},
     {loadUnit_maskInput_lo[16143:16128]},
     {loadUnit_maskInput_lo[16127:16112]},
     {loadUnit_maskInput_lo[16111:16096]},
     {loadUnit_maskInput_lo[16095:16080]},
     {loadUnit_maskInput_lo[16079:16064]},
     {loadUnit_maskInput_lo[16063:16048]},
     {loadUnit_maskInput_lo[16047:16032]},
     {loadUnit_maskInput_lo[16031:16016]},
     {loadUnit_maskInput_lo[16015:16000]},
     {loadUnit_maskInput_lo[15999:15984]},
     {loadUnit_maskInput_lo[15983:15968]},
     {loadUnit_maskInput_lo[15967:15952]},
     {loadUnit_maskInput_lo[15951:15936]},
     {loadUnit_maskInput_lo[15935:15920]},
     {loadUnit_maskInput_lo[15919:15904]},
     {loadUnit_maskInput_lo[15903:15888]},
     {loadUnit_maskInput_lo[15887:15872]},
     {loadUnit_maskInput_lo[15871:15856]},
     {loadUnit_maskInput_lo[15855:15840]},
     {loadUnit_maskInput_lo[15839:15824]},
     {loadUnit_maskInput_lo[15823:15808]},
     {loadUnit_maskInput_lo[15807:15792]},
     {loadUnit_maskInput_lo[15791:15776]},
     {loadUnit_maskInput_lo[15775:15760]},
     {loadUnit_maskInput_lo[15759:15744]},
     {loadUnit_maskInput_lo[15743:15728]},
     {loadUnit_maskInput_lo[15727:15712]},
     {loadUnit_maskInput_lo[15711:15696]},
     {loadUnit_maskInput_lo[15695:15680]},
     {loadUnit_maskInput_lo[15679:15664]},
     {loadUnit_maskInput_lo[15663:15648]},
     {loadUnit_maskInput_lo[15647:15632]},
     {loadUnit_maskInput_lo[15631:15616]},
     {loadUnit_maskInput_lo[15615:15600]},
     {loadUnit_maskInput_lo[15599:15584]},
     {loadUnit_maskInput_lo[15583:15568]},
     {loadUnit_maskInput_lo[15567:15552]},
     {loadUnit_maskInput_lo[15551:15536]},
     {loadUnit_maskInput_lo[15535:15520]},
     {loadUnit_maskInput_lo[15519:15504]},
     {loadUnit_maskInput_lo[15503:15488]},
     {loadUnit_maskInput_lo[15487:15472]},
     {loadUnit_maskInput_lo[15471:15456]},
     {loadUnit_maskInput_lo[15455:15440]},
     {loadUnit_maskInput_lo[15439:15424]},
     {loadUnit_maskInput_lo[15423:15408]},
     {loadUnit_maskInput_lo[15407:15392]},
     {loadUnit_maskInput_lo[15391:15376]},
     {loadUnit_maskInput_lo[15375:15360]},
     {loadUnit_maskInput_lo[15359:15344]},
     {loadUnit_maskInput_lo[15343:15328]},
     {loadUnit_maskInput_lo[15327:15312]},
     {loadUnit_maskInput_lo[15311:15296]},
     {loadUnit_maskInput_lo[15295:15280]},
     {loadUnit_maskInput_lo[15279:15264]},
     {loadUnit_maskInput_lo[15263:15248]},
     {loadUnit_maskInput_lo[15247:15232]},
     {loadUnit_maskInput_lo[15231:15216]},
     {loadUnit_maskInput_lo[15215:15200]},
     {loadUnit_maskInput_lo[15199:15184]},
     {loadUnit_maskInput_lo[15183:15168]},
     {loadUnit_maskInput_lo[15167:15152]},
     {loadUnit_maskInput_lo[15151:15136]},
     {loadUnit_maskInput_lo[15135:15120]},
     {loadUnit_maskInput_lo[15119:15104]},
     {loadUnit_maskInput_lo[15103:15088]},
     {loadUnit_maskInput_lo[15087:15072]},
     {loadUnit_maskInput_lo[15071:15056]},
     {loadUnit_maskInput_lo[15055:15040]},
     {loadUnit_maskInput_lo[15039:15024]},
     {loadUnit_maskInput_lo[15023:15008]},
     {loadUnit_maskInput_lo[15007:14992]},
     {loadUnit_maskInput_lo[14991:14976]},
     {loadUnit_maskInput_lo[14975:14960]},
     {loadUnit_maskInput_lo[14959:14944]},
     {loadUnit_maskInput_lo[14943:14928]},
     {loadUnit_maskInput_lo[14927:14912]},
     {loadUnit_maskInput_lo[14911:14896]},
     {loadUnit_maskInput_lo[14895:14880]},
     {loadUnit_maskInput_lo[14879:14864]},
     {loadUnit_maskInput_lo[14863:14848]},
     {loadUnit_maskInput_lo[14847:14832]},
     {loadUnit_maskInput_lo[14831:14816]},
     {loadUnit_maskInput_lo[14815:14800]},
     {loadUnit_maskInput_lo[14799:14784]},
     {loadUnit_maskInput_lo[14783:14768]},
     {loadUnit_maskInput_lo[14767:14752]},
     {loadUnit_maskInput_lo[14751:14736]},
     {loadUnit_maskInput_lo[14735:14720]},
     {loadUnit_maskInput_lo[14719:14704]},
     {loadUnit_maskInput_lo[14703:14688]},
     {loadUnit_maskInput_lo[14687:14672]},
     {loadUnit_maskInput_lo[14671:14656]},
     {loadUnit_maskInput_lo[14655:14640]},
     {loadUnit_maskInput_lo[14639:14624]},
     {loadUnit_maskInput_lo[14623:14608]},
     {loadUnit_maskInput_lo[14607:14592]},
     {loadUnit_maskInput_lo[14591:14576]},
     {loadUnit_maskInput_lo[14575:14560]},
     {loadUnit_maskInput_lo[14559:14544]},
     {loadUnit_maskInput_lo[14543:14528]},
     {loadUnit_maskInput_lo[14527:14512]},
     {loadUnit_maskInput_lo[14511:14496]},
     {loadUnit_maskInput_lo[14495:14480]},
     {loadUnit_maskInput_lo[14479:14464]},
     {loadUnit_maskInput_lo[14463:14448]},
     {loadUnit_maskInput_lo[14447:14432]},
     {loadUnit_maskInput_lo[14431:14416]},
     {loadUnit_maskInput_lo[14415:14400]},
     {loadUnit_maskInput_lo[14399:14384]},
     {loadUnit_maskInput_lo[14383:14368]},
     {loadUnit_maskInput_lo[14367:14352]},
     {loadUnit_maskInput_lo[14351:14336]},
     {loadUnit_maskInput_lo[14335:14320]},
     {loadUnit_maskInput_lo[14319:14304]},
     {loadUnit_maskInput_lo[14303:14288]},
     {loadUnit_maskInput_lo[14287:14272]},
     {loadUnit_maskInput_lo[14271:14256]},
     {loadUnit_maskInput_lo[14255:14240]},
     {loadUnit_maskInput_lo[14239:14224]},
     {loadUnit_maskInput_lo[14223:14208]},
     {loadUnit_maskInput_lo[14207:14192]},
     {loadUnit_maskInput_lo[14191:14176]},
     {loadUnit_maskInput_lo[14175:14160]},
     {loadUnit_maskInput_lo[14159:14144]},
     {loadUnit_maskInput_lo[14143:14128]},
     {loadUnit_maskInput_lo[14127:14112]},
     {loadUnit_maskInput_lo[14111:14096]},
     {loadUnit_maskInput_lo[14095:14080]},
     {loadUnit_maskInput_lo[14079:14064]},
     {loadUnit_maskInput_lo[14063:14048]},
     {loadUnit_maskInput_lo[14047:14032]},
     {loadUnit_maskInput_lo[14031:14016]},
     {loadUnit_maskInput_lo[14015:14000]},
     {loadUnit_maskInput_lo[13999:13984]},
     {loadUnit_maskInput_lo[13983:13968]},
     {loadUnit_maskInput_lo[13967:13952]},
     {loadUnit_maskInput_lo[13951:13936]},
     {loadUnit_maskInput_lo[13935:13920]},
     {loadUnit_maskInput_lo[13919:13904]},
     {loadUnit_maskInput_lo[13903:13888]},
     {loadUnit_maskInput_lo[13887:13872]},
     {loadUnit_maskInput_lo[13871:13856]},
     {loadUnit_maskInput_lo[13855:13840]},
     {loadUnit_maskInput_lo[13839:13824]},
     {loadUnit_maskInput_lo[13823:13808]},
     {loadUnit_maskInput_lo[13807:13792]},
     {loadUnit_maskInput_lo[13791:13776]},
     {loadUnit_maskInput_lo[13775:13760]},
     {loadUnit_maskInput_lo[13759:13744]},
     {loadUnit_maskInput_lo[13743:13728]},
     {loadUnit_maskInput_lo[13727:13712]},
     {loadUnit_maskInput_lo[13711:13696]},
     {loadUnit_maskInput_lo[13695:13680]},
     {loadUnit_maskInput_lo[13679:13664]},
     {loadUnit_maskInput_lo[13663:13648]},
     {loadUnit_maskInput_lo[13647:13632]},
     {loadUnit_maskInput_lo[13631:13616]},
     {loadUnit_maskInput_lo[13615:13600]},
     {loadUnit_maskInput_lo[13599:13584]},
     {loadUnit_maskInput_lo[13583:13568]},
     {loadUnit_maskInput_lo[13567:13552]},
     {loadUnit_maskInput_lo[13551:13536]},
     {loadUnit_maskInput_lo[13535:13520]},
     {loadUnit_maskInput_lo[13519:13504]},
     {loadUnit_maskInput_lo[13503:13488]},
     {loadUnit_maskInput_lo[13487:13472]},
     {loadUnit_maskInput_lo[13471:13456]},
     {loadUnit_maskInput_lo[13455:13440]},
     {loadUnit_maskInput_lo[13439:13424]},
     {loadUnit_maskInput_lo[13423:13408]},
     {loadUnit_maskInput_lo[13407:13392]},
     {loadUnit_maskInput_lo[13391:13376]},
     {loadUnit_maskInput_lo[13375:13360]},
     {loadUnit_maskInput_lo[13359:13344]},
     {loadUnit_maskInput_lo[13343:13328]},
     {loadUnit_maskInput_lo[13327:13312]},
     {loadUnit_maskInput_lo[13311:13296]},
     {loadUnit_maskInput_lo[13295:13280]},
     {loadUnit_maskInput_lo[13279:13264]},
     {loadUnit_maskInput_lo[13263:13248]},
     {loadUnit_maskInput_lo[13247:13232]},
     {loadUnit_maskInput_lo[13231:13216]},
     {loadUnit_maskInput_lo[13215:13200]},
     {loadUnit_maskInput_lo[13199:13184]},
     {loadUnit_maskInput_lo[13183:13168]},
     {loadUnit_maskInput_lo[13167:13152]},
     {loadUnit_maskInput_lo[13151:13136]},
     {loadUnit_maskInput_lo[13135:13120]},
     {loadUnit_maskInput_lo[13119:13104]},
     {loadUnit_maskInput_lo[13103:13088]},
     {loadUnit_maskInput_lo[13087:13072]},
     {loadUnit_maskInput_lo[13071:13056]},
     {loadUnit_maskInput_lo[13055:13040]},
     {loadUnit_maskInput_lo[13039:13024]},
     {loadUnit_maskInput_lo[13023:13008]},
     {loadUnit_maskInput_lo[13007:12992]},
     {loadUnit_maskInput_lo[12991:12976]},
     {loadUnit_maskInput_lo[12975:12960]},
     {loadUnit_maskInput_lo[12959:12944]},
     {loadUnit_maskInput_lo[12943:12928]},
     {loadUnit_maskInput_lo[12927:12912]},
     {loadUnit_maskInput_lo[12911:12896]},
     {loadUnit_maskInput_lo[12895:12880]},
     {loadUnit_maskInput_lo[12879:12864]},
     {loadUnit_maskInput_lo[12863:12848]},
     {loadUnit_maskInput_lo[12847:12832]},
     {loadUnit_maskInput_lo[12831:12816]},
     {loadUnit_maskInput_lo[12815:12800]},
     {loadUnit_maskInput_lo[12799:12784]},
     {loadUnit_maskInput_lo[12783:12768]},
     {loadUnit_maskInput_lo[12767:12752]},
     {loadUnit_maskInput_lo[12751:12736]},
     {loadUnit_maskInput_lo[12735:12720]},
     {loadUnit_maskInput_lo[12719:12704]},
     {loadUnit_maskInput_lo[12703:12688]},
     {loadUnit_maskInput_lo[12687:12672]},
     {loadUnit_maskInput_lo[12671:12656]},
     {loadUnit_maskInput_lo[12655:12640]},
     {loadUnit_maskInput_lo[12639:12624]},
     {loadUnit_maskInput_lo[12623:12608]},
     {loadUnit_maskInput_lo[12607:12592]},
     {loadUnit_maskInput_lo[12591:12576]},
     {loadUnit_maskInput_lo[12575:12560]},
     {loadUnit_maskInput_lo[12559:12544]},
     {loadUnit_maskInput_lo[12543:12528]},
     {loadUnit_maskInput_lo[12527:12512]},
     {loadUnit_maskInput_lo[12511:12496]},
     {loadUnit_maskInput_lo[12495:12480]},
     {loadUnit_maskInput_lo[12479:12464]},
     {loadUnit_maskInput_lo[12463:12448]},
     {loadUnit_maskInput_lo[12447:12432]},
     {loadUnit_maskInput_lo[12431:12416]},
     {loadUnit_maskInput_lo[12415:12400]},
     {loadUnit_maskInput_lo[12399:12384]},
     {loadUnit_maskInput_lo[12383:12368]},
     {loadUnit_maskInput_lo[12367:12352]},
     {loadUnit_maskInput_lo[12351:12336]},
     {loadUnit_maskInput_lo[12335:12320]},
     {loadUnit_maskInput_lo[12319:12304]},
     {loadUnit_maskInput_lo[12303:12288]},
     {loadUnit_maskInput_lo[12287:12272]},
     {loadUnit_maskInput_lo[12271:12256]},
     {loadUnit_maskInput_lo[12255:12240]},
     {loadUnit_maskInput_lo[12239:12224]},
     {loadUnit_maskInput_lo[12223:12208]},
     {loadUnit_maskInput_lo[12207:12192]},
     {loadUnit_maskInput_lo[12191:12176]},
     {loadUnit_maskInput_lo[12175:12160]},
     {loadUnit_maskInput_lo[12159:12144]},
     {loadUnit_maskInput_lo[12143:12128]},
     {loadUnit_maskInput_lo[12127:12112]},
     {loadUnit_maskInput_lo[12111:12096]},
     {loadUnit_maskInput_lo[12095:12080]},
     {loadUnit_maskInput_lo[12079:12064]},
     {loadUnit_maskInput_lo[12063:12048]},
     {loadUnit_maskInput_lo[12047:12032]},
     {loadUnit_maskInput_lo[12031:12016]},
     {loadUnit_maskInput_lo[12015:12000]},
     {loadUnit_maskInput_lo[11999:11984]},
     {loadUnit_maskInput_lo[11983:11968]},
     {loadUnit_maskInput_lo[11967:11952]},
     {loadUnit_maskInput_lo[11951:11936]},
     {loadUnit_maskInput_lo[11935:11920]},
     {loadUnit_maskInput_lo[11919:11904]},
     {loadUnit_maskInput_lo[11903:11888]},
     {loadUnit_maskInput_lo[11887:11872]},
     {loadUnit_maskInput_lo[11871:11856]},
     {loadUnit_maskInput_lo[11855:11840]},
     {loadUnit_maskInput_lo[11839:11824]},
     {loadUnit_maskInput_lo[11823:11808]},
     {loadUnit_maskInput_lo[11807:11792]},
     {loadUnit_maskInput_lo[11791:11776]},
     {loadUnit_maskInput_lo[11775:11760]},
     {loadUnit_maskInput_lo[11759:11744]},
     {loadUnit_maskInput_lo[11743:11728]},
     {loadUnit_maskInput_lo[11727:11712]},
     {loadUnit_maskInput_lo[11711:11696]},
     {loadUnit_maskInput_lo[11695:11680]},
     {loadUnit_maskInput_lo[11679:11664]},
     {loadUnit_maskInput_lo[11663:11648]},
     {loadUnit_maskInput_lo[11647:11632]},
     {loadUnit_maskInput_lo[11631:11616]},
     {loadUnit_maskInput_lo[11615:11600]},
     {loadUnit_maskInput_lo[11599:11584]},
     {loadUnit_maskInput_lo[11583:11568]},
     {loadUnit_maskInput_lo[11567:11552]},
     {loadUnit_maskInput_lo[11551:11536]},
     {loadUnit_maskInput_lo[11535:11520]},
     {loadUnit_maskInput_lo[11519:11504]},
     {loadUnit_maskInput_lo[11503:11488]},
     {loadUnit_maskInput_lo[11487:11472]},
     {loadUnit_maskInput_lo[11471:11456]},
     {loadUnit_maskInput_lo[11455:11440]},
     {loadUnit_maskInput_lo[11439:11424]},
     {loadUnit_maskInput_lo[11423:11408]},
     {loadUnit_maskInput_lo[11407:11392]},
     {loadUnit_maskInput_lo[11391:11376]},
     {loadUnit_maskInput_lo[11375:11360]},
     {loadUnit_maskInput_lo[11359:11344]},
     {loadUnit_maskInput_lo[11343:11328]},
     {loadUnit_maskInput_lo[11327:11312]},
     {loadUnit_maskInput_lo[11311:11296]},
     {loadUnit_maskInput_lo[11295:11280]},
     {loadUnit_maskInput_lo[11279:11264]},
     {loadUnit_maskInput_lo[11263:11248]},
     {loadUnit_maskInput_lo[11247:11232]},
     {loadUnit_maskInput_lo[11231:11216]},
     {loadUnit_maskInput_lo[11215:11200]},
     {loadUnit_maskInput_lo[11199:11184]},
     {loadUnit_maskInput_lo[11183:11168]},
     {loadUnit_maskInput_lo[11167:11152]},
     {loadUnit_maskInput_lo[11151:11136]},
     {loadUnit_maskInput_lo[11135:11120]},
     {loadUnit_maskInput_lo[11119:11104]},
     {loadUnit_maskInput_lo[11103:11088]},
     {loadUnit_maskInput_lo[11087:11072]},
     {loadUnit_maskInput_lo[11071:11056]},
     {loadUnit_maskInput_lo[11055:11040]},
     {loadUnit_maskInput_lo[11039:11024]},
     {loadUnit_maskInput_lo[11023:11008]},
     {loadUnit_maskInput_lo[11007:10992]},
     {loadUnit_maskInput_lo[10991:10976]},
     {loadUnit_maskInput_lo[10975:10960]},
     {loadUnit_maskInput_lo[10959:10944]},
     {loadUnit_maskInput_lo[10943:10928]},
     {loadUnit_maskInput_lo[10927:10912]},
     {loadUnit_maskInput_lo[10911:10896]},
     {loadUnit_maskInput_lo[10895:10880]},
     {loadUnit_maskInput_lo[10879:10864]},
     {loadUnit_maskInput_lo[10863:10848]},
     {loadUnit_maskInput_lo[10847:10832]},
     {loadUnit_maskInput_lo[10831:10816]},
     {loadUnit_maskInput_lo[10815:10800]},
     {loadUnit_maskInput_lo[10799:10784]},
     {loadUnit_maskInput_lo[10783:10768]},
     {loadUnit_maskInput_lo[10767:10752]},
     {loadUnit_maskInput_lo[10751:10736]},
     {loadUnit_maskInput_lo[10735:10720]},
     {loadUnit_maskInput_lo[10719:10704]},
     {loadUnit_maskInput_lo[10703:10688]},
     {loadUnit_maskInput_lo[10687:10672]},
     {loadUnit_maskInput_lo[10671:10656]},
     {loadUnit_maskInput_lo[10655:10640]},
     {loadUnit_maskInput_lo[10639:10624]},
     {loadUnit_maskInput_lo[10623:10608]},
     {loadUnit_maskInput_lo[10607:10592]},
     {loadUnit_maskInput_lo[10591:10576]},
     {loadUnit_maskInput_lo[10575:10560]},
     {loadUnit_maskInput_lo[10559:10544]},
     {loadUnit_maskInput_lo[10543:10528]},
     {loadUnit_maskInput_lo[10527:10512]},
     {loadUnit_maskInput_lo[10511:10496]},
     {loadUnit_maskInput_lo[10495:10480]},
     {loadUnit_maskInput_lo[10479:10464]},
     {loadUnit_maskInput_lo[10463:10448]},
     {loadUnit_maskInput_lo[10447:10432]},
     {loadUnit_maskInput_lo[10431:10416]},
     {loadUnit_maskInput_lo[10415:10400]},
     {loadUnit_maskInput_lo[10399:10384]},
     {loadUnit_maskInput_lo[10383:10368]},
     {loadUnit_maskInput_lo[10367:10352]},
     {loadUnit_maskInput_lo[10351:10336]},
     {loadUnit_maskInput_lo[10335:10320]},
     {loadUnit_maskInput_lo[10319:10304]},
     {loadUnit_maskInput_lo[10303:10288]},
     {loadUnit_maskInput_lo[10287:10272]},
     {loadUnit_maskInput_lo[10271:10256]},
     {loadUnit_maskInput_lo[10255:10240]},
     {loadUnit_maskInput_lo[10239:10224]},
     {loadUnit_maskInput_lo[10223:10208]},
     {loadUnit_maskInput_lo[10207:10192]},
     {loadUnit_maskInput_lo[10191:10176]},
     {loadUnit_maskInput_lo[10175:10160]},
     {loadUnit_maskInput_lo[10159:10144]},
     {loadUnit_maskInput_lo[10143:10128]},
     {loadUnit_maskInput_lo[10127:10112]},
     {loadUnit_maskInput_lo[10111:10096]},
     {loadUnit_maskInput_lo[10095:10080]},
     {loadUnit_maskInput_lo[10079:10064]},
     {loadUnit_maskInput_lo[10063:10048]},
     {loadUnit_maskInput_lo[10047:10032]},
     {loadUnit_maskInput_lo[10031:10016]},
     {loadUnit_maskInput_lo[10015:10000]},
     {loadUnit_maskInput_lo[9999:9984]},
     {loadUnit_maskInput_lo[9983:9968]},
     {loadUnit_maskInput_lo[9967:9952]},
     {loadUnit_maskInput_lo[9951:9936]},
     {loadUnit_maskInput_lo[9935:9920]},
     {loadUnit_maskInput_lo[9919:9904]},
     {loadUnit_maskInput_lo[9903:9888]},
     {loadUnit_maskInput_lo[9887:9872]},
     {loadUnit_maskInput_lo[9871:9856]},
     {loadUnit_maskInput_lo[9855:9840]},
     {loadUnit_maskInput_lo[9839:9824]},
     {loadUnit_maskInput_lo[9823:9808]},
     {loadUnit_maskInput_lo[9807:9792]},
     {loadUnit_maskInput_lo[9791:9776]},
     {loadUnit_maskInput_lo[9775:9760]},
     {loadUnit_maskInput_lo[9759:9744]},
     {loadUnit_maskInput_lo[9743:9728]},
     {loadUnit_maskInput_lo[9727:9712]},
     {loadUnit_maskInput_lo[9711:9696]},
     {loadUnit_maskInput_lo[9695:9680]},
     {loadUnit_maskInput_lo[9679:9664]},
     {loadUnit_maskInput_lo[9663:9648]},
     {loadUnit_maskInput_lo[9647:9632]},
     {loadUnit_maskInput_lo[9631:9616]},
     {loadUnit_maskInput_lo[9615:9600]},
     {loadUnit_maskInput_lo[9599:9584]},
     {loadUnit_maskInput_lo[9583:9568]},
     {loadUnit_maskInput_lo[9567:9552]},
     {loadUnit_maskInput_lo[9551:9536]},
     {loadUnit_maskInput_lo[9535:9520]},
     {loadUnit_maskInput_lo[9519:9504]},
     {loadUnit_maskInput_lo[9503:9488]},
     {loadUnit_maskInput_lo[9487:9472]},
     {loadUnit_maskInput_lo[9471:9456]},
     {loadUnit_maskInput_lo[9455:9440]},
     {loadUnit_maskInput_lo[9439:9424]},
     {loadUnit_maskInput_lo[9423:9408]},
     {loadUnit_maskInput_lo[9407:9392]},
     {loadUnit_maskInput_lo[9391:9376]},
     {loadUnit_maskInput_lo[9375:9360]},
     {loadUnit_maskInput_lo[9359:9344]},
     {loadUnit_maskInput_lo[9343:9328]},
     {loadUnit_maskInput_lo[9327:9312]},
     {loadUnit_maskInput_lo[9311:9296]},
     {loadUnit_maskInput_lo[9295:9280]},
     {loadUnit_maskInput_lo[9279:9264]},
     {loadUnit_maskInput_lo[9263:9248]},
     {loadUnit_maskInput_lo[9247:9232]},
     {loadUnit_maskInput_lo[9231:9216]},
     {loadUnit_maskInput_lo[9215:9200]},
     {loadUnit_maskInput_lo[9199:9184]},
     {loadUnit_maskInput_lo[9183:9168]},
     {loadUnit_maskInput_lo[9167:9152]},
     {loadUnit_maskInput_lo[9151:9136]},
     {loadUnit_maskInput_lo[9135:9120]},
     {loadUnit_maskInput_lo[9119:9104]},
     {loadUnit_maskInput_lo[9103:9088]},
     {loadUnit_maskInput_lo[9087:9072]},
     {loadUnit_maskInput_lo[9071:9056]},
     {loadUnit_maskInput_lo[9055:9040]},
     {loadUnit_maskInput_lo[9039:9024]},
     {loadUnit_maskInput_lo[9023:9008]},
     {loadUnit_maskInput_lo[9007:8992]},
     {loadUnit_maskInput_lo[8991:8976]},
     {loadUnit_maskInput_lo[8975:8960]},
     {loadUnit_maskInput_lo[8959:8944]},
     {loadUnit_maskInput_lo[8943:8928]},
     {loadUnit_maskInput_lo[8927:8912]},
     {loadUnit_maskInput_lo[8911:8896]},
     {loadUnit_maskInput_lo[8895:8880]},
     {loadUnit_maskInput_lo[8879:8864]},
     {loadUnit_maskInput_lo[8863:8848]},
     {loadUnit_maskInput_lo[8847:8832]},
     {loadUnit_maskInput_lo[8831:8816]},
     {loadUnit_maskInput_lo[8815:8800]},
     {loadUnit_maskInput_lo[8799:8784]},
     {loadUnit_maskInput_lo[8783:8768]},
     {loadUnit_maskInput_lo[8767:8752]},
     {loadUnit_maskInput_lo[8751:8736]},
     {loadUnit_maskInput_lo[8735:8720]},
     {loadUnit_maskInput_lo[8719:8704]},
     {loadUnit_maskInput_lo[8703:8688]},
     {loadUnit_maskInput_lo[8687:8672]},
     {loadUnit_maskInput_lo[8671:8656]},
     {loadUnit_maskInput_lo[8655:8640]},
     {loadUnit_maskInput_lo[8639:8624]},
     {loadUnit_maskInput_lo[8623:8608]},
     {loadUnit_maskInput_lo[8607:8592]},
     {loadUnit_maskInput_lo[8591:8576]},
     {loadUnit_maskInput_lo[8575:8560]},
     {loadUnit_maskInput_lo[8559:8544]},
     {loadUnit_maskInput_lo[8543:8528]},
     {loadUnit_maskInput_lo[8527:8512]},
     {loadUnit_maskInput_lo[8511:8496]},
     {loadUnit_maskInput_lo[8495:8480]},
     {loadUnit_maskInput_lo[8479:8464]},
     {loadUnit_maskInput_lo[8463:8448]},
     {loadUnit_maskInput_lo[8447:8432]},
     {loadUnit_maskInput_lo[8431:8416]},
     {loadUnit_maskInput_lo[8415:8400]},
     {loadUnit_maskInput_lo[8399:8384]},
     {loadUnit_maskInput_lo[8383:8368]},
     {loadUnit_maskInput_lo[8367:8352]},
     {loadUnit_maskInput_lo[8351:8336]},
     {loadUnit_maskInput_lo[8335:8320]},
     {loadUnit_maskInput_lo[8319:8304]},
     {loadUnit_maskInput_lo[8303:8288]},
     {loadUnit_maskInput_lo[8287:8272]},
     {loadUnit_maskInput_lo[8271:8256]},
     {loadUnit_maskInput_lo[8255:8240]},
     {loadUnit_maskInput_lo[8239:8224]},
     {loadUnit_maskInput_lo[8223:8208]},
     {loadUnit_maskInput_lo[8207:8192]},
     {loadUnit_maskInput_lo[8191:8176]},
     {loadUnit_maskInput_lo[8175:8160]},
     {loadUnit_maskInput_lo[8159:8144]},
     {loadUnit_maskInput_lo[8143:8128]},
     {loadUnit_maskInput_lo[8127:8112]},
     {loadUnit_maskInput_lo[8111:8096]},
     {loadUnit_maskInput_lo[8095:8080]},
     {loadUnit_maskInput_lo[8079:8064]},
     {loadUnit_maskInput_lo[8063:8048]},
     {loadUnit_maskInput_lo[8047:8032]},
     {loadUnit_maskInput_lo[8031:8016]},
     {loadUnit_maskInput_lo[8015:8000]},
     {loadUnit_maskInput_lo[7999:7984]},
     {loadUnit_maskInput_lo[7983:7968]},
     {loadUnit_maskInput_lo[7967:7952]},
     {loadUnit_maskInput_lo[7951:7936]},
     {loadUnit_maskInput_lo[7935:7920]},
     {loadUnit_maskInput_lo[7919:7904]},
     {loadUnit_maskInput_lo[7903:7888]},
     {loadUnit_maskInput_lo[7887:7872]},
     {loadUnit_maskInput_lo[7871:7856]},
     {loadUnit_maskInput_lo[7855:7840]},
     {loadUnit_maskInput_lo[7839:7824]},
     {loadUnit_maskInput_lo[7823:7808]},
     {loadUnit_maskInput_lo[7807:7792]},
     {loadUnit_maskInput_lo[7791:7776]},
     {loadUnit_maskInput_lo[7775:7760]},
     {loadUnit_maskInput_lo[7759:7744]},
     {loadUnit_maskInput_lo[7743:7728]},
     {loadUnit_maskInput_lo[7727:7712]},
     {loadUnit_maskInput_lo[7711:7696]},
     {loadUnit_maskInput_lo[7695:7680]},
     {loadUnit_maskInput_lo[7679:7664]},
     {loadUnit_maskInput_lo[7663:7648]},
     {loadUnit_maskInput_lo[7647:7632]},
     {loadUnit_maskInput_lo[7631:7616]},
     {loadUnit_maskInput_lo[7615:7600]},
     {loadUnit_maskInput_lo[7599:7584]},
     {loadUnit_maskInput_lo[7583:7568]},
     {loadUnit_maskInput_lo[7567:7552]},
     {loadUnit_maskInput_lo[7551:7536]},
     {loadUnit_maskInput_lo[7535:7520]},
     {loadUnit_maskInput_lo[7519:7504]},
     {loadUnit_maskInput_lo[7503:7488]},
     {loadUnit_maskInput_lo[7487:7472]},
     {loadUnit_maskInput_lo[7471:7456]},
     {loadUnit_maskInput_lo[7455:7440]},
     {loadUnit_maskInput_lo[7439:7424]},
     {loadUnit_maskInput_lo[7423:7408]},
     {loadUnit_maskInput_lo[7407:7392]},
     {loadUnit_maskInput_lo[7391:7376]},
     {loadUnit_maskInput_lo[7375:7360]},
     {loadUnit_maskInput_lo[7359:7344]},
     {loadUnit_maskInput_lo[7343:7328]},
     {loadUnit_maskInput_lo[7327:7312]},
     {loadUnit_maskInput_lo[7311:7296]},
     {loadUnit_maskInput_lo[7295:7280]},
     {loadUnit_maskInput_lo[7279:7264]},
     {loadUnit_maskInput_lo[7263:7248]},
     {loadUnit_maskInput_lo[7247:7232]},
     {loadUnit_maskInput_lo[7231:7216]},
     {loadUnit_maskInput_lo[7215:7200]},
     {loadUnit_maskInput_lo[7199:7184]},
     {loadUnit_maskInput_lo[7183:7168]},
     {loadUnit_maskInput_lo[7167:7152]},
     {loadUnit_maskInput_lo[7151:7136]},
     {loadUnit_maskInput_lo[7135:7120]},
     {loadUnit_maskInput_lo[7119:7104]},
     {loadUnit_maskInput_lo[7103:7088]},
     {loadUnit_maskInput_lo[7087:7072]},
     {loadUnit_maskInput_lo[7071:7056]},
     {loadUnit_maskInput_lo[7055:7040]},
     {loadUnit_maskInput_lo[7039:7024]},
     {loadUnit_maskInput_lo[7023:7008]},
     {loadUnit_maskInput_lo[7007:6992]},
     {loadUnit_maskInput_lo[6991:6976]},
     {loadUnit_maskInput_lo[6975:6960]},
     {loadUnit_maskInput_lo[6959:6944]},
     {loadUnit_maskInput_lo[6943:6928]},
     {loadUnit_maskInput_lo[6927:6912]},
     {loadUnit_maskInput_lo[6911:6896]},
     {loadUnit_maskInput_lo[6895:6880]},
     {loadUnit_maskInput_lo[6879:6864]},
     {loadUnit_maskInput_lo[6863:6848]},
     {loadUnit_maskInput_lo[6847:6832]},
     {loadUnit_maskInput_lo[6831:6816]},
     {loadUnit_maskInput_lo[6815:6800]},
     {loadUnit_maskInput_lo[6799:6784]},
     {loadUnit_maskInput_lo[6783:6768]},
     {loadUnit_maskInput_lo[6767:6752]},
     {loadUnit_maskInput_lo[6751:6736]},
     {loadUnit_maskInput_lo[6735:6720]},
     {loadUnit_maskInput_lo[6719:6704]},
     {loadUnit_maskInput_lo[6703:6688]},
     {loadUnit_maskInput_lo[6687:6672]},
     {loadUnit_maskInput_lo[6671:6656]},
     {loadUnit_maskInput_lo[6655:6640]},
     {loadUnit_maskInput_lo[6639:6624]},
     {loadUnit_maskInput_lo[6623:6608]},
     {loadUnit_maskInput_lo[6607:6592]},
     {loadUnit_maskInput_lo[6591:6576]},
     {loadUnit_maskInput_lo[6575:6560]},
     {loadUnit_maskInput_lo[6559:6544]},
     {loadUnit_maskInput_lo[6543:6528]},
     {loadUnit_maskInput_lo[6527:6512]},
     {loadUnit_maskInput_lo[6511:6496]},
     {loadUnit_maskInput_lo[6495:6480]},
     {loadUnit_maskInput_lo[6479:6464]},
     {loadUnit_maskInput_lo[6463:6448]},
     {loadUnit_maskInput_lo[6447:6432]},
     {loadUnit_maskInput_lo[6431:6416]},
     {loadUnit_maskInput_lo[6415:6400]},
     {loadUnit_maskInput_lo[6399:6384]},
     {loadUnit_maskInput_lo[6383:6368]},
     {loadUnit_maskInput_lo[6367:6352]},
     {loadUnit_maskInput_lo[6351:6336]},
     {loadUnit_maskInput_lo[6335:6320]},
     {loadUnit_maskInput_lo[6319:6304]},
     {loadUnit_maskInput_lo[6303:6288]},
     {loadUnit_maskInput_lo[6287:6272]},
     {loadUnit_maskInput_lo[6271:6256]},
     {loadUnit_maskInput_lo[6255:6240]},
     {loadUnit_maskInput_lo[6239:6224]},
     {loadUnit_maskInput_lo[6223:6208]},
     {loadUnit_maskInput_lo[6207:6192]},
     {loadUnit_maskInput_lo[6191:6176]},
     {loadUnit_maskInput_lo[6175:6160]},
     {loadUnit_maskInput_lo[6159:6144]},
     {loadUnit_maskInput_lo[6143:6128]},
     {loadUnit_maskInput_lo[6127:6112]},
     {loadUnit_maskInput_lo[6111:6096]},
     {loadUnit_maskInput_lo[6095:6080]},
     {loadUnit_maskInput_lo[6079:6064]},
     {loadUnit_maskInput_lo[6063:6048]},
     {loadUnit_maskInput_lo[6047:6032]},
     {loadUnit_maskInput_lo[6031:6016]},
     {loadUnit_maskInput_lo[6015:6000]},
     {loadUnit_maskInput_lo[5999:5984]},
     {loadUnit_maskInput_lo[5983:5968]},
     {loadUnit_maskInput_lo[5967:5952]},
     {loadUnit_maskInput_lo[5951:5936]},
     {loadUnit_maskInput_lo[5935:5920]},
     {loadUnit_maskInput_lo[5919:5904]},
     {loadUnit_maskInput_lo[5903:5888]},
     {loadUnit_maskInput_lo[5887:5872]},
     {loadUnit_maskInput_lo[5871:5856]},
     {loadUnit_maskInput_lo[5855:5840]},
     {loadUnit_maskInput_lo[5839:5824]},
     {loadUnit_maskInput_lo[5823:5808]},
     {loadUnit_maskInput_lo[5807:5792]},
     {loadUnit_maskInput_lo[5791:5776]},
     {loadUnit_maskInput_lo[5775:5760]},
     {loadUnit_maskInput_lo[5759:5744]},
     {loadUnit_maskInput_lo[5743:5728]},
     {loadUnit_maskInput_lo[5727:5712]},
     {loadUnit_maskInput_lo[5711:5696]},
     {loadUnit_maskInput_lo[5695:5680]},
     {loadUnit_maskInput_lo[5679:5664]},
     {loadUnit_maskInput_lo[5663:5648]},
     {loadUnit_maskInput_lo[5647:5632]},
     {loadUnit_maskInput_lo[5631:5616]},
     {loadUnit_maskInput_lo[5615:5600]},
     {loadUnit_maskInput_lo[5599:5584]},
     {loadUnit_maskInput_lo[5583:5568]},
     {loadUnit_maskInput_lo[5567:5552]},
     {loadUnit_maskInput_lo[5551:5536]},
     {loadUnit_maskInput_lo[5535:5520]},
     {loadUnit_maskInput_lo[5519:5504]},
     {loadUnit_maskInput_lo[5503:5488]},
     {loadUnit_maskInput_lo[5487:5472]},
     {loadUnit_maskInput_lo[5471:5456]},
     {loadUnit_maskInput_lo[5455:5440]},
     {loadUnit_maskInput_lo[5439:5424]},
     {loadUnit_maskInput_lo[5423:5408]},
     {loadUnit_maskInput_lo[5407:5392]},
     {loadUnit_maskInput_lo[5391:5376]},
     {loadUnit_maskInput_lo[5375:5360]},
     {loadUnit_maskInput_lo[5359:5344]},
     {loadUnit_maskInput_lo[5343:5328]},
     {loadUnit_maskInput_lo[5327:5312]},
     {loadUnit_maskInput_lo[5311:5296]},
     {loadUnit_maskInput_lo[5295:5280]},
     {loadUnit_maskInput_lo[5279:5264]},
     {loadUnit_maskInput_lo[5263:5248]},
     {loadUnit_maskInput_lo[5247:5232]},
     {loadUnit_maskInput_lo[5231:5216]},
     {loadUnit_maskInput_lo[5215:5200]},
     {loadUnit_maskInput_lo[5199:5184]},
     {loadUnit_maskInput_lo[5183:5168]},
     {loadUnit_maskInput_lo[5167:5152]},
     {loadUnit_maskInput_lo[5151:5136]},
     {loadUnit_maskInput_lo[5135:5120]},
     {loadUnit_maskInput_lo[5119:5104]},
     {loadUnit_maskInput_lo[5103:5088]},
     {loadUnit_maskInput_lo[5087:5072]},
     {loadUnit_maskInput_lo[5071:5056]},
     {loadUnit_maskInput_lo[5055:5040]},
     {loadUnit_maskInput_lo[5039:5024]},
     {loadUnit_maskInput_lo[5023:5008]},
     {loadUnit_maskInput_lo[5007:4992]},
     {loadUnit_maskInput_lo[4991:4976]},
     {loadUnit_maskInput_lo[4975:4960]},
     {loadUnit_maskInput_lo[4959:4944]},
     {loadUnit_maskInput_lo[4943:4928]},
     {loadUnit_maskInput_lo[4927:4912]},
     {loadUnit_maskInput_lo[4911:4896]},
     {loadUnit_maskInput_lo[4895:4880]},
     {loadUnit_maskInput_lo[4879:4864]},
     {loadUnit_maskInput_lo[4863:4848]},
     {loadUnit_maskInput_lo[4847:4832]},
     {loadUnit_maskInput_lo[4831:4816]},
     {loadUnit_maskInput_lo[4815:4800]},
     {loadUnit_maskInput_lo[4799:4784]},
     {loadUnit_maskInput_lo[4783:4768]},
     {loadUnit_maskInput_lo[4767:4752]},
     {loadUnit_maskInput_lo[4751:4736]},
     {loadUnit_maskInput_lo[4735:4720]},
     {loadUnit_maskInput_lo[4719:4704]},
     {loadUnit_maskInput_lo[4703:4688]},
     {loadUnit_maskInput_lo[4687:4672]},
     {loadUnit_maskInput_lo[4671:4656]},
     {loadUnit_maskInput_lo[4655:4640]},
     {loadUnit_maskInput_lo[4639:4624]},
     {loadUnit_maskInput_lo[4623:4608]},
     {loadUnit_maskInput_lo[4607:4592]},
     {loadUnit_maskInput_lo[4591:4576]},
     {loadUnit_maskInput_lo[4575:4560]},
     {loadUnit_maskInput_lo[4559:4544]},
     {loadUnit_maskInput_lo[4543:4528]},
     {loadUnit_maskInput_lo[4527:4512]},
     {loadUnit_maskInput_lo[4511:4496]},
     {loadUnit_maskInput_lo[4495:4480]},
     {loadUnit_maskInput_lo[4479:4464]},
     {loadUnit_maskInput_lo[4463:4448]},
     {loadUnit_maskInput_lo[4447:4432]},
     {loadUnit_maskInput_lo[4431:4416]},
     {loadUnit_maskInput_lo[4415:4400]},
     {loadUnit_maskInput_lo[4399:4384]},
     {loadUnit_maskInput_lo[4383:4368]},
     {loadUnit_maskInput_lo[4367:4352]},
     {loadUnit_maskInput_lo[4351:4336]},
     {loadUnit_maskInput_lo[4335:4320]},
     {loadUnit_maskInput_lo[4319:4304]},
     {loadUnit_maskInput_lo[4303:4288]},
     {loadUnit_maskInput_lo[4287:4272]},
     {loadUnit_maskInput_lo[4271:4256]},
     {loadUnit_maskInput_lo[4255:4240]},
     {loadUnit_maskInput_lo[4239:4224]},
     {loadUnit_maskInput_lo[4223:4208]},
     {loadUnit_maskInput_lo[4207:4192]},
     {loadUnit_maskInput_lo[4191:4176]},
     {loadUnit_maskInput_lo[4175:4160]},
     {loadUnit_maskInput_lo[4159:4144]},
     {loadUnit_maskInput_lo[4143:4128]},
     {loadUnit_maskInput_lo[4127:4112]},
     {loadUnit_maskInput_lo[4111:4096]},
     {loadUnit_maskInput_lo[4095:4080]},
     {loadUnit_maskInput_lo[4079:4064]},
     {loadUnit_maskInput_lo[4063:4048]},
     {loadUnit_maskInput_lo[4047:4032]},
     {loadUnit_maskInput_lo[4031:4016]},
     {loadUnit_maskInput_lo[4015:4000]},
     {loadUnit_maskInput_lo[3999:3984]},
     {loadUnit_maskInput_lo[3983:3968]},
     {loadUnit_maskInput_lo[3967:3952]},
     {loadUnit_maskInput_lo[3951:3936]},
     {loadUnit_maskInput_lo[3935:3920]},
     {loadUnit_maskInput_lo[3919:3904]},
     {loadUnit_maskInput_lo[3903:3888]},
     {loadUnit_maskInput_lo[3887:3872]},
     {loadUnit_maskInput_lo[3871:3856]},
     {loadUnit_maskInput_lo[3855:3840]},
     {loadUnit_maskInput_lo[3839:3824]},
     {loadUnit_maskInput_lo[3823:3808]},
     {loadUnit_maskInput_lo[3807:3792]},
     {loadUnit_maskInput_lo[3791:3776]},
     {loadUnit_maskInput_lo[3775:3760]},
     {loadUnit_maskInput_lo[3759:3744]},
     {loadUnit_maskInput_lo[3743:3728]},
     {loadUnit_maskInput_lo[3727:3712]},
     {loadUnit_maskInput_lo[3711:3696]},
     {loadUnit_maskInput_lo[3695:3680]},
     {loadUnit_maskInput_lo[3679:3664]},
     {loadUnit_maskInput_lo[3663:3648]},
     {loadUnit_maskInput_lo[3647:3632]},
     {loadUnit_maskInput_lo[3631:3616]},
     {loadUnit_maskInput_lo[3615:3600]},
     {loadUnit_maskInput_lo[3599:3584]},
     {loadUnit_maskInput_lo[3583:3568]},
     {loadUnit_maskInput_lo[3567:3552]},
     {loadUnit_maskInput_lo[3551:3536]},
     {loadUnit_maskInput_lo[3535:3520]},
     {loadUnit_maskInput_lo[3519:3504]},
     {loadUnit_maskInput_lo[3503:3488]},
     {loadUnit_maskInput_lo[3487:3472]},
     {loadUnit_maskInput_lo[3471:3456]},
     {loadUnit_maskInput_lo[3455:3440]},
     {loadUnit_maskInput_lo[3439:3424]},
     {loadUnit_maskInput_lo[3423:3408]},
     {loadUnit_maskInput_lo[3407:3392]},
     {loadUnit_maskInput_lo[3391:3376]},
     {loadUnit_maskInput_lo[3375:3360]},
     {loadUnit_maskInput_lo[3359:3344]},
     {loadUnit_maskInput_lo[3343:3328]},
     {loadUnit_maskInput_lo[3327:3312]},
     {loadUnit_maskInput_lo[3311:3296]},
     {loadUnit_maskInput_lo[3295:3280]},
     {loadUnit_maskInput_lo[3279:3264]},
     {loadUnit_maskInput_lo[3263:3248]},
     {loadUnit_maskInput_lo[3247:3232]},
     {loadUnit_maskInput_lo[3231:3216]},
     {loadUnit_maskInput_lo[3215:3200]},
     {loadUnit_maskInput_lo[3199:3184]},
     {loadUnit_maskInput_lo[3183:3168]},
     {loadUnit_maskInput_lo[3167:3152]},
     {loadUnit_maskInput_lo[3151:3136]},
     {loadUnit_maskInput_lo[3135:3120]},
     {loadUnit_maskInput_lo[3119:3104]},
     {loadUnit_maskInput_lo[3103:3088]},
     {loadUnit_maskInput_lo[3087:3072]},
     {loadUnit_maskInput_lo[3071:3056]},
     {loadUnit_maskInput_lo[3055:3040]},
     {loadUnit_maskInput_lo[3039:3024]},
     {loadUnit_maskInput_lo[3023:3008]},
     {loadUnit_maskInput_lo[3007:2992]},
     {loadUnit_maskInput_lo[2991:2976]},
     {loadUnit_maskInput_lo[2975:2960]},
     {loadUnit_maskInput_lo[2959:2944]},
     {loadUnit_maskInput_lo[2943:2928]},
     {loadUnit_maskInput_lo[2927:2912]},
     {loadUnit_maskInput_lo[2911:2896]},
     {loadUnit_maskInput_lo[2895:2880]},
     {loadUnit_maskInput_lo[2879:2864]},
     {loadUnit_maskInput_lo[2863:2848]},
     {loadUnit_maskInput_lo[2847:2832]},
     {loadUnit_maskInput_lo[2831:2816]},
     {loadUnit_maskInput_lo[2815:2800]},
     {loadUnit_maskInput_lo[2799:2784]},
     {loadUnit_maskInput_lo[2783:2768]},
     {loadUnit_maskInput_lo[2767:2752]},
     {loadUnit_maskInput_lo[2751:2736]},
     {loadUnit_maskInput_lo[2735:2720]},
     {loadUnit_maskInput_lo[2719:2704]},
     {loadUnit_maskInput_lo[2703:2688]},
     {loadUnit_maskInput_lo[2687:2672]},
     {loadUnit_maskInput_lo[2671:2656]},
     {loadUnit_maskInput_lo[2655:2640]},
     {loadUnit_maskInput_lo[2639:2624]},
     {loadUnit_maskInput_lo[2623:2608]},
     {loadUnit_maskInput_lo[2607:2592]},
     {loadUnit_maskInput_lo[2591:2576]},
     {loadUnit_maskInput_lo[2575:2560]},
     {loadUnit_maskInput_lo[2559:2544]},
     {loadUnit_maskInput_lo[2543:2528]},
     {loadUnit_maskInput_lo[2527:2512]},
     {loadUnit_maskInput_lo[2511:2496]},
     {loadUnit_maskInput_lo[2495:2480]},
     {loadUnit_maskInput_lo[2479:2464]},
     {loadUnit_maskInput_lo[2463:2448]},
     {loadUnit_maskInput_lo[2447:2432]},
     {loadUnit_maskInput_lo[2431:2416]},
     {loadUnit_maskInput_lo[2415:2400]},
     {loadUnit_maskInput_lo[2399:2384]},
     {loadUnit_maskInput_lo[2383:2368]},
     {loadUnit_maskInput_lo[2367:2352]},
     {loadUnit_maskInput_lo[2351:2336]},
     {loadUnit_maskInput_lo[2335:2320]},
     {loadUnit_maskInput_lo[2319:2304]},
     {loadUnit_maskInput_lo[2303:2288]},
     {loadUnit_maskInput_lo[2287:2272]},
     {loadUnit_maskInput_lo[2271:2256]},
     {loadUnit_maskInput_lo[2255:2240]},
     {loadUnit_maskInput_lo[2239:2224]},
     {loadUnit_maskInput_lo[2223:2208]},
     {loadUnit_maskInput_lo[2207:2192]},
     {loadUnit_maskInput_lo[2191:2176]},
     {loadUnit_maskInput_lo[2175:2160]},
     {loadUnit_maskInput_lo[2159:2144]},
     {loadUnit_maskInput_lo[2143:2128]},
     {loadUnit_maskInput_lo[2127:2112]},
     {loadUnit_maskInput_lo[2111:2096]},
     {loadUnit_maskInput_lo[2095:2080]},
     {loadUnit_maskInput_lo[2079:2064]},
     {loadUnit_maskInput_lo[2063:2048]},
     {loadUnit_maskInput_lo[2047:2032]},
     {loadUnit_maskInput_lo[2031:2016]},
     {loadUnit_maskInput_lo[2015:2000]},
     {loadUnit_maskInput_lo[1999:1984]},
     {loadUnit_maskInput_lo[1983:1968]},
     {loadUnit_maskInput_lo[1967:1952]},
     {loadUnit_maskInput_lo[1951:1936]},
     {loadUnit_maskInput_lo[1935:1920]},
     {loadUnit_maskInput_lo[1919:1904]},
     {loadUnit_maskInput_lo[1903:1888]},
     {loadUnit_maskInput_lo[1887:1872]},
     {loadUnit_maskInput_lo[1871:1856]},
     {loadUnit_maskInput_lo[1855:1840]},
     {loadUnit_maskInput_lo[1839:1824]},
     {loadUnit_maskInput_lo[1823:1808]},
     {loadUnit_maskInput_lo[1807:1792]},
     {loadUnit_maskInput_lo[1791:1776]},
     {loadUnit_maskInput_lo[1775:1760]},
     {loadUnit_maskInput_lo[1759:1744]},
     {loadUnit_maskInput_lo[1743:1728]},
     {loadUnit_maskInput_lo[1727:1712]},
     {loadUnit_maskInput_lo[1711:1696]},
     {loadUnit_maskInput_lo[1695:1680]},
     {loadUnit_maskInput_lo[1679:1664]},
     {loadUnit_maskInput_lo[1663:1648]},
     {loadUnit_maskInput_lo[1647:1632]},
     {loadUnit_maskInput_lo[1631:1616]},
     {loadUnit_maskInput_lo[1615:1600]},
     {loadUnit_maskInput_lo[1599:1584]},
     {loadUnit_maskInput_lo[1583:1568]},
     {loadUnit_maskInput_lo[1567:1552]},
     {loadUnit_maskInput_lo[1551:1536]},
     {loadUnit_maskInput_lo[1535:1520]},
     {loadUnit_maskInput_lo[1519:1504]},
     {loadUnit_maskInput_lo[1503:1488]},
     {loadUnit_maskInput_lo[1487:1472]},
     {loadUnit_maskInput_lo[1471:1456]},
     {loadUnit_maskInput_lo[1455:1440]},
     {loadUnit_maskInput_lo[1439:1424]},
     {loadUnit_maskInput_lo[1423:1408]},
     {loadUnit_maskInput_lo[1407:1392]},
     {loadUnit_maskInput_lo[1391:1376]},
     {loadUnit_maskInput_lo[1375:1360]},
     {loadUnit_maskInput_lo[1359:1344]},
     {loadUnit_maskInput_lo[1343:1328]},
     {loadUnit_maskInput_lo[1327:1312]},
     {loadUnit_maskInput_lo[1311:1296]},
     {loadUnit_maskInput_lo[1295:1280]},
     {loadUnit_maskInput_lo[1279:1264]},
     {loadUnit_maskInput_lo[1263:1248]},
     {loadUnit_maskInput_lo[1247:1232]},
     {loadUnit_maskInput_lo[1231:1216]},
     {loadUnit_maskInput_lo[1215:1200]},
     {loadUnit_maskInput_lo[1199:1184]},
     {loadUnit_maskInput_lo[1183:1168]},
     {loadUnit_maskInput_lo[1167:1152]},
     {loadUnit_maskInput_lo[1151:1136]},
     {loadUnit_maskInput_lo[1135:1120]},
     {loadUnit_maskInput_lo[1119:1104]},
     {loadUnit_maskInput_lo[1103:1088]},
     {loadUnit_maskInput_lo[1087:1072]},
     {loadUnit_maskInput_lo[1071:1056]},
     {loadUnit_maskInput_lo[1055:1040]},
     {loadUnit_maskInput_lo[1039:1024]},
     {loadUnit_maskInput_lo[1023:1008]},
     {loadUnit_maskInput_lo[1007:992]},
     {loadUnit_maskInput_lo[991:976]},
     {loadUnit_maskInput_lo[975:960]},
     {loadUnit_maskInput_lo[959:944]},
     {loadUnit_maskInput_lo[943:928]},
     {loadUnit_maskInput_lo[927:912]},
     {loadUnit_maskInput_lo[911:896]},
     {loadUnit_maskInput_lo[895:880]},
     {loadUnit_maskInput_lo[879:864]},
     {loadUnit_maskInput_lo[863:848]},
     {loadUnit_maskInput_lo[847:832]},
     {loadUnit_maskInput_lo[831:816]},
     {loadUnit_maskInput_lo[815:800]},
     {loadUnit_maskInput_lo[799:784]},
     {loadUnit_maskInput_lo[783:768]},
     {loadUnit_maskInput_lo[767:752]},
     {loadUnit_maskInput_lo[751:736]},
     {loadUnit_maskInput_lo[735:720]},
     {loadUnit_maskInput_lo[719:704]},
     {loadUnit_maskInput_lo[703:688]},
     {loadUnit_maskInput_lo[687:672]},
     {loadUnit_maskInput_lo[671:656]},
     {loadUnit_maskInput_lo[655:640]},
     {loadUnit_maskInput_lo[639:624]},
     {loadUnit_maskInput_lo[623:608]},
     {loadUnit_maskInput_lo[607:592]},
     {loadUnit_maskInput_lo[591:576]},
     {loadUnit_maskInput_lo[575:560]},
     {loadUnit_maskInput_lo[559:544]},
     {loadUnit_maskInput_lo[543:528]},
     {loadUnit_maskInput_lo[527:512]},
     {loadUnit_maskInput_lo[511:496]},
     {loadUnit_maskInput_lo[495:480]},
     {loadUnit_maskInput_lo[479:464]},
     {loadUnit_maskInput_lo[463:448]},
     {loadUnit_maskInput_lo[447:432]},
     {loadUnit_maskInput_lo[431:416]},
     {loadUnit_maskInput_lo[415:400]},
     {loadUnit_maskInput_lo[399:384]},
     {loadUnit_maskInput_lo[383:368]},
     {loadUnit_maskInput_lo[367:352]},
     {loadUnit_maskInput_lo[351:336]},
     {loadUnit_maskInput_lo[335:320]},
     {loadUnit_maskInput_lo[319:304]},
     {loadUnit_maskInput_lo[303:288]},
     {loadUnit_maskInput_lo[287:272]},
     {loadUnit_maskInput_lo[271:256]},
     {loadUnit_maskInput_lo[255:240]},
     {loadUnit_maskInput_lo[239:224]},
     {loadUnit_maskInput_lo[223:208]},
     {loadUnit_maskInput_lo[207:192]},
     {loadUnit_maskInput_lo[191:176]},
     {loadUnit_maskInput_lo[175:160]},
     {loadUnit_maskInput_lo[159:144]},
     {loadUnit_maskInput_lo[143:128]},
     {loadUnit_maskInput_lo[127:112]},
     {loadUnit_maskInput_lo[111:96]},
     {loadUnit_maskInput_lo[95:80]},
     {loadUnit_maskInput_lo[79:64]},
     {loadUnit_maskInput_lo[63:48]},
     {loadUnit_maskInput_lo[47:32]},
     {loadUnit_maskInput_lo[31:16]},
     {loadUnit_maskInput_lo[15:0]}};
  wire [11:0]         maskSelect_1 = _storeUnit_maskSelect_valid ? _storeUnit_maskSelect_bits : 12'h0;
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi = {storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo = {storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi = {storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi = {storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo = {storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi = {storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo = {storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo = {storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi = {storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi = {storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi = {storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_lo_lo_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi = {storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo = {storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo = {storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi = {storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi = {storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo = {storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo = {storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi = {storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo = {storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo = {storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi = {storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi = {storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi = {storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_lo_lo_lo_lo_hi = {storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo};
  wire [2047:0]       storeUnit_maskInput_lo_lo_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi = {storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo = {storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi = {storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi = {storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo = {storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo = {storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi = {storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo = {storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo = {storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi = {storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi = {storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi = {storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_lo_lo_lo_hi_lo = {storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi = {storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo = {storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo = {storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi = {storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi = {storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo = {storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo = {storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi = {storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo = {storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo = {storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi = {storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi = {storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi = {storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_lo_lo_lo_hi_hi = {storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo};
  wire [2047:0]       storeUnit_maskInput_lo_lo_lo_lo_hi = {storeUnit_maskInput_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_lo};
  wire [4095:0]       storeUnit_maskInput_lo_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi = {storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo = {storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi = {storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi = {storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo = {storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi = {storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo = {storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo = {storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi = {storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi = {storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi = {storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_lo_lo_hi_lo_lo = {storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi = {storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo = {storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo = {storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi = {storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi = {storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo = {storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo = {storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi = {storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo = {storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo = {storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi = {storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi = {storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi = {storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_lo_lo_hi_lo_hi = {storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo};
  wire [2047:0]       storeUnit_maskInput_lo_lo_lo_hi_lo = {storeUnit_maskInput_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi = {storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo = {storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi = {storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi = {storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo = {storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo = {storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi = {storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo = {storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo = {storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi = {storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi = {storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi = {storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_lo_lo_hi_hi_lo = {storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi = {storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo = {storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo = {storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi = {storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi = {storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo = {storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo = {storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi = {storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo = {storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo = {storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi = {storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi = {storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi = {storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_lo_lo_hi_hi_hi = {storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo};
  wire [2047:0]       storeUnit_maskInput_lo_lo_lo_hi_hi = {storeUnit_maskInput_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_lo};
  wire [4095:0]       storeUnit_maskInput_lo_lo_lo_hi = {storeUnit_maskInput_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_lo};
  wire [8191:0]       storeUnit_maskInput_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo = {storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi = {storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo = {storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo = {storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi = {storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi = {storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo = {storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo = {storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi = {storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo = {storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo = {storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi = {storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi = {storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi = {storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_lo_hi_lo_lo_lo = {storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo = {storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi = {storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo = {storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo = {storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi = {storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi = {storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo = {storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo = {storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi = {storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo = {storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo = {storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi = {storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi = {storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi = {storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_lo_hi_lo_lo_hi = {storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo};
  wire [2047:0]       storeUnit_maskInput_lo_lo_hi_lo_lo = {storeUnit_maskInput_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo = {storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi = {storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo = {storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo = {storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi = {storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi = {storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo = {storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo = {storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi = {storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo = {storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo = {storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi = {storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi = {storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi = {storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_lo_hi_lo_hi_lo = {storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo = {storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi = {storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo = {storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo = {storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi = {storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi = {storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo = {storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo = {storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi = {storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo = {storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo = {storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi = {storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi = {storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi = {storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_lo_hi_lo_hi_hi = {storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo};
  wire [2047:0]       storeUnit_maskInput_lo_lo_hi_lo_hi = {storeUnit_maskInput_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_lo};
  wire [4095:0]       storeUnit_maskInput_lo_lo_hi_lo = {storeUnit_maskInput_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo = {storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi = {storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo = {storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo = {storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi = {storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi = {storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo = {storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo = {storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi = {storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo = {storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo = {storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi = {storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi = {storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi = {storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_lo_hi_hi_lo_lo = {storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo = {storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi = {storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo = {storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo = {storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi = {storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi = {storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo = {storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo = {storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi = {storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo = {storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo = {storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi = {storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi = {storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi = {storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_lo_hi_hi_lo_hi = {storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo};
  wire [2047:0]       storeUnit_maskInput_lo_lo_hi_hi_lo = {storeUnit_maskInput_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo = {storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi = {storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo = {storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo = {storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi = {storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi = {storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo = {storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo = {storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi = {storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo = {storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo = {storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi = {storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi = {storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi = {storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_lo_hi_hi_hi_lo = {storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo = {storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi = {storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo = {storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo = {storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi = {storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi = {storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo = {storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo = {storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi = {storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo = {storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo = {storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi = {storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi = {storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi = {storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_lo_hi_hi_hi_hi = {storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo};
  wire [2047:0]       storeUnit_maskInput_lo_lo_hi_hi_hi = {storeUnit_maskInput_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_lo};
  wire [4095:0]       storeUnit_maskInput_lo_lo_hi_hi = {storeUnit_maskInput_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_lo};
  wire [8191:0]       storeUnit_maskInput_lo_lo_hi = {storeUnit_maskInput_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo};
  wire [16383:0]      storeUnit_maskInput_lo_lo = {storeUnit_maskInput_lo_lo_hi, storeUnit_maskInput_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo = {storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi = {storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo = {storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi = {storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi = {storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo = {storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo = {storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi = {storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo = {storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi = {storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi = {storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi = {storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_hi_lo_lo_lo_lo = {storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo = {storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi = {storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo = {storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi = {storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi = {storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo = {storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi = {storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo = {storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo = {storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi = {storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi = {storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi = {storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_hi_lo_lo_lo_hi = {storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo};
  wire [2047:0]       storeUnit_maskInput_lo_hi_lo_lo_lo = {storeUnit_maskInput_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo = {storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi = {storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo = {storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi = {storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi = {storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo = {storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo = {storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi = {storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo = {storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi = {storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi = {storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi = {storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_hi_lo_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo = {storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi = {storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo = {storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi = {storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi = {storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo = {storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo = {storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi = {storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo = {storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo = {storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi = {storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi = {storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi = {storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_hi_lo_lo_hi_hi = {storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo};
  wire [2047:0]       storeUnit_maskInput_lo_hi_lo_lo_hi = {storeUnit_maskInput_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_lo};
  wire [4095:0]       storeUnit_maskInput_lo_hi_lo_lo = {storeUnit_maskInput_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo = {storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi = {storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo = {storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi = {storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi = {storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo = {storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo = {storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi = {storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi = {storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi = {storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi = {storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_hi_lo_hi_lo_lo = {storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo = {storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi = {storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo = {storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi = {storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi = {storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo = {storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi = {storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi = {storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi = {storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi = {storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_hi_lo_hi_lo_hi = {storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo};
  wire [2047:0]       storeUnit_maskInput_lo_hi_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo = {storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi = {storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo = {storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi = {storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi = {storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo = {storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo = {storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi = {storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi = {storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi = {storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi = {storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_hi_lo_hi_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo = {storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi = {storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo = {storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi = {storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi = {storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo = {storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi = {storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi = {storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi = {storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi = {storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_hi_lo_hi_hi_hi = {storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo};
  wire [2047:0]       storeUnit_maskInput_lo_hi_lo_hi_hi = {storeUnit_maskInput_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_lo};
  wire [4095:0]       storeUnit_maskInput_lo_hi_lo_hi = {storeUnit_maskInput_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_lo};
  wire [8191:0]       storeUnit_maskInput_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo = {storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi = {storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo = {storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo = {storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi = {storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi = {storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo = {storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo = {storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi = {storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo = {storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo = {storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi = {storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi = {storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi = {storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_hi_hi_lo_lo_lo = {storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo = {storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi = {storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo = {storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo = {storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi = {storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi = {storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo = {storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo = {storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi = {storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo = {storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo = {storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi = {storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi = {storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi = {storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_hi_hi_lo_lo_hi = {storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo};
  wire [2047:0]       storeUnit_maskInput_lo_hi_hi_lo_lo = {storeUnit_maskInput_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo = {storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi = {storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo = {storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo = {storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi = {storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi = {storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo = {storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo = {storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi = {storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo = {storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo = {storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi = {storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi = {storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi = {storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_hi_hi_lo_hi_lo = {storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo = {storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi = {storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo = {storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo = {storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi = {storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi = {storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo = {storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo = {storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi = {storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo = {storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo = {storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi = {storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi = {storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi = {storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_hi_hi_lo_hi_hi = {storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo};
  wire [2047:0]       storeUnit_maskInput_lo_hi_hi_lo_hi = {storeUnit_maskInput_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_lo};
  wire [4095:0]       storeUnit_maskInput_lo_hi_hi_lo = {storeUnit_maskInput_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo = {storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi = {storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo = {storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo = {storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi = {storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo = {storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo = {storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi = {storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo = {storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo = {storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi = {storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_hi_hi_hi_lo_lo = {storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo = {storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi = {storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo = {storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo = {storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi = {storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo = {storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo = {storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi = {storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo = {storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo = {storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_hi_hi_hi_lo_hi = {storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo};
  wire [2047:0]       storeUnit_maskInput_lo_hi_hi_hi_lo = {storeUnit_maskInput_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo = {storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi = {storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo = {storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo = {storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi = {storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo = {storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo = {storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi = {storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo = {storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo = {storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi = {storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_hi_hi_hi_hi_lo = {storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo = {storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi = {storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo = {storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo = {storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi = {storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo = {storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo = {storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi = {storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo = {storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo = {storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_hi_hi_hi_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo};
  wire [2047:0]       storeUnit_maskInput_lo_hi_hi_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_lo};
  wire [4095:0]       storeUnit_maskInput_lo_hi_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_lo};
  wire [8191:0]       storeUnit_maskInput_lo_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_lo};
  wire [16383:0]      storeUnit_maskInput_lo_hi = {storeUnit_maskInput_lo_hi_hi, storeUnit_maskInput_lo_hi_lo};
  wire [32767:0]      storeUnit_maskInput_lo = {storeUnit_maskInput_lo_hi, storeUnit_maskInput_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo = {storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi = {storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo = {storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo = {storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi = {storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi = {storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo = {storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo = {storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi = {storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo = {storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo = {storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi = {storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi = {storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi = {storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_lo_lo_lo_lo_lo = {storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo = {storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi = {storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo = {storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo = {storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi = {storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi = {storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo = {storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo = {storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi = {storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo = {storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo = {storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi = {storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi = {storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi = {storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_lo_lo_lo_lo_hi = {storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo};
  wire [2047:0]       storeUnit_maskInput_hi_lo_lo_lo_lo = {storeUnit_maskInput_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo = {storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi = {storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo = {storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo = {storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi = {storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi = {storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo = {storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo = {storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi = {storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo = {storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo = {storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi = {storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi = {storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi = {storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_lo_lo_lo_hi_lo = {storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo = {storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi = {storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo = {storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo = {storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi = {storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi = {storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo = {storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo = {storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi = {storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo = {storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo = {storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi = {storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi = {storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi = {storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_lo_lo_lo_hi_hi = {storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo};
  wire [2047:0]       storeUnit_maskInput_hi_lo_lo_lo_hi = {storeUnit_maskInput_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_lo};
  wire [4095:0]       storeUnit_maskInput_hi_lo_lo_lo = {storeUnit_maskInput_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo = {storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi = {storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo = {storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo = {storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi = {storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi = {storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo = {storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo = {storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi = {storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo = {storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo = {storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi = {storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi = {storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi = {storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_lo_lo_hi_lo_lo = {storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo = {storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi = {storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo = {storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo = {storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi = {storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi = {storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo = {storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo = {storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi = {storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo = {storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo = {storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi = {storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi = {storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi = {storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_lo_lo_hi_lo_hi = {storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo};
  wire [2047:0]       storeUnit_maskInput_hi_lo_lo_hi_lo = {storeUnit_maskInput_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo = {storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi = {storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo = {storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo = {storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi = {storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi = {storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo = {storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo = {storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi = {storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo = {storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo = {storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi = {storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi = {storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi = {storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_lo_lo_hi_hi_lo = {storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo = {storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi = {storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo = {storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo = {storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi = {storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi = {storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo = {storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo = {storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi = {storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo = {storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo = {storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi = {storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi = {storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi = {storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_lo_lo_hi_hi_hi = {storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo};
  wire [2047:0]       storeUnit_maskInput_hi_lo_lo_hi_hi = {storeUnit_maskInput_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_lo};
  wire [4095:0]       storeUnit_maskInput_hi_lo_lo_hi = {storeUnit_maskInput_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_lo};
  wire [8191:0]       storeUnit_maskInput_hi_lo_lo = {storeUnit_maskInput_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo = {storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi = {storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo = {storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo = {storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi = {storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi = {storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo = {storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo = {storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo = {storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo = {storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi = {storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi = {storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi = {storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_lo_hi_lo_lo_lo = {storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo = {storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi = {storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo = {storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo = {storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi = {storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo = {storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo = {storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo = {storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo = {storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi = {storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi = {storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi = {storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_lo_hi_lo_lo_hi = {storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo};
  wire [2047:0]       storeUnit_maskInput_hi_lo_hi_lo_lo = {storeUnit_maskInput_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo = {storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi = {storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo = {storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo = {storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi = {storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi = {storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo = {storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo = {storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo = {storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo = {storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi = {storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi = {storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_lo_hi_lo_hi_lo = {storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo = {storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi = {storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo = {storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo = {storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi = {storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo = {storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo = {storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo = {storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo = {storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi = {storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi = {storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi = {storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_lo_hi_lo_hi_hi = {storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo};
  wire [2047:0]       storeUnit_maskInput_hi_lo_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_lo};
  wire [4095:0]       storeUnit_maskInput_hi_lo_hi_lo = {storeUnit_maskInput_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo = {storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi = {storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo = {storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo = {storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi = {storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi = {storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo = {storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo = {storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo = {storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo = {storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi = {storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi = {storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi = {storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_lo_hi_hi_lo_lo = {storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo = {storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi = {storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo = {storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo = {storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi = {storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo = {storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo = {storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo = {storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo = {storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi = {storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi = {storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi = {storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_lo_hi_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo};
  wire [2047:0]       storeUnit_maskInput_hi_lo_hi_hi_lo = {storeUnit_maskInput_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo = {storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi = {storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo = {storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo = {storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi = {storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi = {storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo = {storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo = {storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo = {storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo = {storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi = {storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi = {storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_lo_hi_hi_hi_lo = {storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo = {storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi = {storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo = {storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo = {storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi = {storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo = {storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo = {storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo = {storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo = {storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi = {storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi = {storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi = {storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_lo_hi_hi_hi_hi = {storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo};
  wire [2047:0]       storeUnit_maskInput_hi_lo_hi_hi_hi = {storeUnit_maskInput_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_lo};
  wire [4095:0]       storeUnit_maskInput_hi_lo_hi_hi = {storeUnit_maskInput_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_lo};
  wire [8191:0]       storeUnit_maskInput_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo};
  wire [16383:0]      storeUnit_maskInput_hi_lo = {storeUnit_maskInput_hi_lo_hi, storeUnit_maskInput_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo = {storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi = {storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo = {storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo = {storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi = {storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi = {storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo = {storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo = {storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi = {storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo = {storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo = {storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi = {storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi = {storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi = {storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_hi_lo_lo_lo_lo = {storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo = {storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi = {storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo = {storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo = {storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi = {storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi = {storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo = {storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo = {storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi = {storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo = {storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo = {storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi = {storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi = {storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi = {storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_hi_lo_lo_lo_hi = {storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo};
  wire [2047:0]       storeUnit_maskInput_hi_hi_lo_lo_lo = {storeUnit_maskInput_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo = {storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi = {storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo = {storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo = {storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi = {storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi = {storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo = {storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo = {storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi = {storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo = {storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo = {storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi = {storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi = {storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi = {storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_hi_lo_lo_hi_lo = {storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo = {storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi = {storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo = {storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo = {storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi = {storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi = {storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo = {storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo = {storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi = {storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo = {storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo = {storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi = {storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi = {storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi = {storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_hi_lo_lo_hi_hi = {storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo};
  wire [2047:0]       storeUnit_maskInput_hi_hi_lo_lo_hi = {storeUnit_maskInput_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_lo};
  wire [4095:0]       storeUnit_maskInput_hi_hi_lo_lo = {storeUnit_maskInput_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo = {storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi = {storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo = {storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi = {storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi = {storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo = {storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo = {storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi = {storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi = {storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi = {storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi = {storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_hi_lo_hi_lo_lo = {storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo = {storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi = {storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo = {storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi = {storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi = {storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo = {storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi = {storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi = {storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi = {storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi = {storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_hi_lo_hi_lo_hi = {storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo};
  wire [2047:0]       storeUnit_maskInput_hi_hi_lo_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo = {storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi = {storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo = {storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi = {storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi = {storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo = {storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo = {storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi = {storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi = {storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi = {storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi = {storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_hi_lo_hi_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo = {storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi = {storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo = {storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi = {storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi = {storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo = {storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi = {storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi = {storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi = {storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi = {storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_hi_lo_hi_hi_hi = {storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo};
  wire [2047:0]       storeUnit_maskInput_hi_hi_lo_hi_hi = {storeUnit_maskInput_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_lo};
  wire [4095:0]       storeUnit_maskInput_hi_hi_lo_hi = {storeUnit_maskInput_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_lo};
  wire [8191:0]       storeUnit_maskInput_hi_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo = {storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi = {storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo = {storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo = {storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi = {storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi = {storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo = {storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo = {storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi = {storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo = {storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo = {storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi = {storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi = {storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_hi_hi_lo_lo_lo = {storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo = {storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi = {storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo = {storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo = {storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi = {storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi = {storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo = {storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo = {storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi = {storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo = {storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo = {storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi = {storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_hi_hi_lo_lo_hi = {storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo};
  wire [2047:0]       storeUnit_maskInput_hi_hi_hi_lo_lo = {storeUnit_maskInput_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo = {storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi = {storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo = {storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo = {storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi = {storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi = {storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo = {storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo = {storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi = {storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo = {storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo = {storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi = {storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi = {storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_hi_hi_lo_hi_lo = {storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo = {storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi = {storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo = {storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo = {storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi = {storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi = {storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo = {storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo = {storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi = {storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo = {storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo = {storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_hi_hi_lo_hi_hi = {storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo};
  wire [2047:0]       storeUnit_maskInput_hi_hi_hi_lo_hi = {storeUnit_maskInput_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_lo};
  wire [4095:0]       storeUnit_maskInput_hi_hi_hi_lo = {storeUnit_maskInput_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo = {storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi = {storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo = {storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo = {storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi = {storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo = {storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo = {storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi = {storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo = {storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo = {storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi = {storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_hi_hi_hi_lo_lo = {storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo = {storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi = {storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo = {storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo = {storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi = {storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo = {storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo = {storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi = {storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo = {storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo = {storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_hi_hi_hi_lo_hi = {storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo};
  wire [2047:0]       storeUnit_maskInput_hi_hi_hi_hi_lo = {storeUnit_maskInput_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo = {storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi = {storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo = {storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo = {storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi = {storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo = {storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo = {storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi = {storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo = {storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo = {storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi = {storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_hi_hi_hi_hi_lo = {storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo = {storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi = {storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo = {storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo = {storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi = {storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo = {storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo = {storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi = {storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo = {storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo = {storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_hi_hi_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo};
  wire [2047:0]       storeUnit_maskInput_hi_hi_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_lo};
  wire [4095:0]       storeUnit_maskInput_hi_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_lo};
  wire [8191:0]       storeUnit_maskInput_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_lo};
  wire [16383:0]      storeUnit_maskInput_hi_hi = {storeUnit_maskInput_hi_hi_hi, storeUnit_maskInput_hi_hi_lo};
  wire [32767:0]      storeUnit_maskInput_hi = {storeUnit_maskInput_hi_hi, storeUnit_maskInput_hi_lo};
  wire [4095:0][15:0] _GEN_1024 =
    {{storeUnit_maskInput_hi[32767:32752]},
     {storeUnit_maskInput_hi[32751:32736]},
     {storeUnit_maskInput_hi[32735:32720]},
     {storeUnit_maskInput_hi[32719:32704]},
     {storeUnit_maskInput_hi[32703:32688]},
     {storeUnit_maskInput_hi[32687:32672]},
     {storeUnit_maskInput_hi[32671:32656]},
     {storeUnit_maskInput_hi[32655:32640]},
     {storeUnit_maskInput_hi[32639:32624]},
     {storeUnit_maskInput_hi[32623:32608]},
     {storeUnit_maskInput_hi[32607:32592]},
     {storeUnit_maskInput_hi[32591:32576]},
     {storeUnit_maskInput_hi[32575:32560]},
     {storeUnit_maskInput_hi[32559:32544]},
     {storeUnit_maskInput_hi[32543:32528]},
     {storeUnit_maskInput_hi[32527:32512]},
     {storeUnit_maskInput_hi[32511:32496]},
     {storeUnit_maskInput_hi[32495:32480]},
     {storeUnit_maskInput_hi[32479:32464]},
     {storeUnit_maskInput_hi[32463:32448]},
     {storeUnit_maskInput_hi[32447:32432]},
     {storeUnit_maskInput_hi[32431:32416]},
     {storeUnit_maskInput_hi[32415:32400]},
     {storeUnit_maskInput_hi[32399:32384]},
     {storeUnit_maskInput_hi[32383:32368]},
     {storeUnit_maskInput_hi[32367:32352]},
     {storeUnit_maskInput_hi[32351:32336]},
     {storeUnit_maskInput_hi[32335:32320]},
     {storeUnit_maskInput_hi[32319:32304]},
     {storeUnit_maskInput_hi[32303:32288]},
     {storeUnit_maskInput_hi[32287:32272]},
     {storeUnit_maskInput_hi[32271:32256]},
     {storeUnit_maskInput_hi[32255:32240]},
     {storeUnit_maskInput_hi[32239:32224]},
     {storeUnit_maskInput_hi[32223:32208]},
     {storeUnit_maskInput_hi[32207:32192]},
     {storeUnit_maskInput_hi[32191:32176]},
     {storeUnit_maskInput_hi[32175:32160]},
     {storeUnit_maskInput_hi[32159:32144]},
     {storeUnit_maskInput_hi[32143:32128]},
     {storeUnit_maskInput_hi[32127:32112]},
     {storeUnit_maskInput_hi[32111:32096]},
     {storeUnit_maskInput_hi[32095:32080]},
     {storeUnit_maskInput_hi[32079:32064]},
     {storeUnit_maskInput_hi[32063:32048]},
     {storeUnit_maskInput_hi[32047:32032]},
     {storeUnit_maskInput_hi[32031:32016]},
     {storeUnit_maskInput_hi[32015:32000]},
     {storeUnit_maskInput_hi[31999:31984]},
     {storeUnit_maskInput_hi[31983:31968]},
     {storeUnit_maskInput_hi[31967:31952]},
     {storeUnit_maskInput_hi[31951:31936]},
     {storeUnit_maskInput_hi[31935:31920]},
     {storeUnit_maskInput_hi[31919:31904]},
     {storeUnit_maskInput_hi[31903:31888]},
     {storeUnit_maskInput_hi[31887:31872]},
     {storeUnit_maskInput_hi[31871:31856]},
     {storeUnit_maskInput_hi[31855:31840]},
     {storeUnit_maskInput_hi[31839:31824]},
     {storeUnit_maskInput_hi[31823:31808]},
     {storeUnit_maskInput_hi[31807:31792]},
     {storeUnit_maskInput_hi[31791:31776]},
     {storeUnit_maskInput_hi[31775:31760]},
     {storeUnit_maskInput_hi[31759:31744]},
     {storeUnit_maskInput_hi[31743:31728]},
     {storeUnit_maskInput_hi[31727:31712]},
     {storeUnit_maskInput_hi[31711:31696]},
     {storeUnit_maskInput_hi[31695:31680]},
     {storeUnit_maskInput_hi[31679:31664]},
     {storeUnit_maskInput_hi[31663:31648]},
     {storeUnit_maskInput_hi[31647:31632]},
     {storeUnit_maskInput_hi[31631:31616]},
     {storeUnit_maskInput_hi[31615:31600]},
     {storeUnit_maskInput_hi[31599:31584]},
     {storeUnit_maskInput_hi[31583:31568]},
     {storeUnit_maskInput_hi[31567:31552]},
     {storeUnit_maskInput_hi[31551:31536]},
     {storeUnit_maskInput_hi[31535:31520]},
     {storeUnit_maskInput_hi[31519:31504]},
     {storeUnit_maskInput_hi[31503:31488]},
     {storeUnit_maskInput_hi[31487:31472]},
     {storeUnit_maskInput_hi[31471:31456]},
     {storeUnit_maskInput_hi[31455:31440]},
     {storeUnit_maskInput_hi[31439:31424]},
     {storeUnit_maskInput_hi[31423:31408]},
     {storeUnit_maskInput_hi[31407:31392]},
     {storeUnit_maskInput_hi[31391:31376]},
     {storeUnit_maskInput_hi[31375:31360]},
     {storeUnit_maskInput_hi[31359:31344]},
     {storeUnit_maskInput_hi[31343:31328]},
     {storeUnit_maskInput_hi[31327:31312]},
     {storeUnit_maskInput_hi[31311:31296]},
     {storeUnit_maskInput_hi[31295:31280]},
     {storeUnit_maskInput_hi[31279:31264]},
     {storeUnit_maskInput_hi[31263:31248]},
     {storeUnit_maskInput_hi[31247:31232]},
     {storeUnit_maskInput_hi[31231:31216]},
     {storeUnit_maskInput_hi[31215:31200]},
     {storeUnit_maskInput_hi[31199:31184]},
     {storeUnit_maskInput_hi[31183:31168]},
     {storeUnit_maskInput_hi[31167:31152]},
     {storeUnit_maskInput_hi[31151:31136]},
     {storeUnit_maskInput_hi[31135:31120]},
     {storeUnit_maskInput_hi[31119:31104]},
     {storeUnit_maskInput_hi[31103:31088]},
     {storeUnit_maskInput_hi[31087:31072]},
     {storeUnit_maskInput_hi[31071:31056]},
     {storeUnit_maskInput_hi[31055:31040]},
     {storeUnit_maskInput_hi[31039:31024]},
     {storeUnit_maskInput_hi[31023:31008]},
     {storeUnit_maskInput_hi[31007:30992]},
     {storeUnit_maskInput_hi[30991:30976]},
     {storeUnit_maskInput_hi[30975:30960]},
     {storeUnit_maskInput_hi[30959:30944]},
     {storeUnit_maskInput_hi[30943:30928]},
     {storeUnit_maskInput_hi[30927:30912]},
     {storeUnit_maskInput_hi[30911:30896]},
     {storeUnit_maskInput_hi[30895:30880]},
     {storeUnit_maskInput_hi[30879:30864]},
     {storeUnit_maskInput_hi[30863:30848]},
     {storeUnit_maskInput_hi[30847:30832]},
     {storeUnit_maskInput_hi[30831:30816]},
     {storeUnit_maskInput_hi[30815:30800]},
     {storeUnit_maskInput_hi[30799:30784]},
     {storeUnit_maskInput_hi[30783:30768]},
     {storeUnit_maskInput_hi[30767:30752]},
     {storeUnit_maskInput_hi[30751:30736]},
     {storeUnit_maskInput_hi[30735:30720]},
     {storeUnit_maskInput_hi[30719:30704]},
     {storeUnit_maskInput_hi[30703:30688]},
     {storeUnit_maskInput_hi[30687:30672]},
     {storeUnit_maskInput_hi[30671:30656]},
     {storeUnit_maskInput_hi[30655:30640]},
     {storeUnit_maskInput_hi[30639:30624]},
     {storeUnit_maskInput_hi[30623:30608]},
     {storeUnit_maskInput_hi[30607:30592]},
     {storeUnit_maskInput_hi[30591:30576]},
     {storeUnit_maskInput_hi[30575:30560]},
     {storeUnit_maskInput_hi[30559:30544]},
     {storeUnit_maskInput_hi[30543:30528]},
     {storeUnit_maskInput_hi[30527:30512]},
     {storeUnit_maskInput_hi[30511:30496]},
     {storeUnit_maskInput_hi[30495:30480]},
     {storeUnit_maskInput_hi[30479:30464]},
     {storeUnit_maskInput_hi[30463:30448]},
     {storeUnit_maskInput_hi[30447:30432]},
     {storeUnit_maskInput_hi[30431:30416]},
     {storeUnit_maskInput_hi[30415:30400]},
     {storeUnit_maskInput_hi[30399:30384]},
     {storeUnit_maskInput_hi[30383:30368]},
     {storeUnit_maskInput_hi[30367:30352]},
     {storeUnit_maskInput_hi[30351:30336]},
     {storeUnit_maskInput_hi[30335:30320]},
     {storeUnit_maskInput_hi[30319:30304]},
     {storeUnit_maskInput_hi[30303:30288]},
     {storeUnit_maskInput_hi[30287:30272]},
     {storeUnit_maskInput_hi[30271:30256]},
     {storeUnit_maskInput_hi[30255:30240]},
     {storeUnit_maskInput_hi[30239:30224]},
     {storeUnit_maskInput_hi[30223:30208]},
     {storeUnit_maskInput_hi[30207:30192]},
     {storeUnit_maskInput_hi[30191:30176]},
     {storeUnit_maskInput_hi[30175:30160]},
     {storeUnit_maskInput_hi[30159:30144]},
     {storeUnit_maskInput_hi[30143:30128]},
     {storeUnit_maskInput_hi[30127:30112]},
     {storeUnit_maskInput_hi[30111:30096]},
     {storeUnit_maskInput_hi[30095:30080]},
     {storeUnit_maskInput_hi[30079:30064]},
     {storeUnit_maskInput_hi[30063:30048]},
     {storeUnit_maskInput_hi[30047:30032]},
     {storeUnit_maskInput_hi[30031:30016]},
     {storeUnit_maskInput_hi[30015:30000]},
     {storeUnit_maskInput_hi[29999:29984]},
     {storeUnit_maskInput_hi[29983:29968]},
     {storeUnit_maskInput_hi[29967:29952]},
     {storeUnit_maskInput_hi[29951:29936]},
     {storeUnit_maskInput_hi[29935:29920]},
     {storeUnit_maskInput_hi[29919:29904]},
     {storeUnit_maskInput_hi[29903:29888]},
     {storeUnit_maskInput_hi[29887:29872]},
     {storeUnit_maskInput_hi[29871:29856]},
     {storeUnit_maskInput_hi[29855:29840]},
     {storeUnit_maskInput_hi[29839:29824]},
     {storeUnit_maskInput_hi[29823:29808]},
     {storeUnit_maskInput_hi[29807:29792]},
     {storeUnit_maskInput_hi[29791:29776]},
     {storeUnit_maskInput_hi[29775:29760]},
     {storeUnit_maskInput_hi[29759:29744]},
     {storeUnit_maskInput_hi[29743:29728]},
     {storeUnit_maskInput_hi[29727:29712]},
     {storeUnit_maskInput_hi[29711:29696]},
     {storeUnit_maskInput_hi[29695:29680]},
     {storeUnit_maskInput_hi[29679:29664]},
     {storeUnit_maskInput_hi[29663:29648]},
     {storeUnit_maskInput_hi[29647:29632]},
     {storeUnit_maskInput_hi[29631:29616]},
     {storeUnit_maskInput_hi[29615:29600]},
     {storeUnit_maskInput_hi[29599:29584]},
     {storeUnit_maskInput_hi[29583:29568]},
     {storeUnit_maskInput_hi[29567:29552]},
     {storeUnit_maskInput_hi[29551:29536]},
     {storeUnit_maskInput_hi[29535:29520]},
     {storeUnit_maskInput_hi[29519:29504]},
     {storeUnit_maskInput_hi[29503:29488]},
     {storeUnit_maskInput_hi[29487:29472]},
     {storeUnit_maskInput_hi[29471:29456]},
     {storeUnit_maskInput_hi[29455:29440]},
     {storeUnit_maskInput_hi[29439:29424]},
     {storeUnit_maskInput_hi[29423:29408]},
     {storeUnit_maskInput_hi[29407:29392]},
     {storeUnit_maskInput_hi[29391:29376]},
     {storeUnit_maskInput_hi[29375:29360]},
     {storeUnit_maskInput_hi[29359:29344]},
     {storeUnit_maskInput_hi[29343:29328]},
     {storeUnit_maskInput_hi[29327:29312]},
     {storeUnit_maskInput_hi[29311:29296]},
     {storeUnit_maskInput_hi[29295:29280]},
     {storeUnit_maskInput_hi[29279:29264]},
     {storeUnit_maskInput_hi[29263:29248]},
     {storeUnit_maskInput_hi[29247:29232]},
     {storeUnit_maskInput_hi[29231:29216]},
     {storeUnit_maskInput_hi[29215:29200]},
     {storeUnit_maskInput_hi[29199:29184]},
     {storeUnit_maskInput_hi[29183:29168]},
     {storeUnit_maskInput_hi[29167:29152]},
     {storeUnit_maskInput_hi[29151:29136]},
     {storeUnit_maskInput_hi[29135:29120]},
     {storeUnit_maskInput_hi[29119:29104]},
     {storeUnit_maskInput_hi[29103:29088]},
     {storeUnit_maskInput_hi[29087:29072]},
     {storeUnit_maskInput_hi[29071:29056]},
     {storeUnit_maskInput_hi[29055:29040]},
     {storeUnit_maskInput_hi[29039:29024]},
     {storeUnit_maskInput_hi[29023:29008]},
     {storeUnit_maskInput_hi[29007:28992]},
     {storeUnit_maskInput_hi[28991:28976]},
     {storeUnit_maskInput_hi[28975:28960]},
     {storeUnit_maskInput_hi[28959:28944]},
     {storeUnit_maskInput_hi[28943:28928]},
     {storeUnit_maskInput_hi[28927:28912]},
     {storeUnit_maskInput_hi[28911:28896]},
     {storeUnit_maskInput_hi[28895:28880]},
     {storeUnit_maskInput_hi[28879:28864]},
     {storeUnit_maskInput_hi[28863:28848]},
     {storeUnit_maskInput_hi[28847:28832]},
     {storeUnit_maskInput_hi[28831:28816]},
     {storeUnit_maskInput_hi[28815:28800]},
     {storeUnit_maskInput_hi[28799:28784]},
     {storeUnit_maskInput_hi[28783:28768]},
     {storeUnit_maskInput_hi[28767:28752]},
     {storeUnit_maskInput_hi[28751:28736]},
     {storeUnit_maskInput_hi[28735:28720]},
     {storeUnit_maskInput_hi[28719:28704]},
     {storeUnit_maskInput_hi[28703:28688]},
     {storeUnit_maskInput_hi[28687:28672]},
     {storeUnit_maskInput_hi[28671:28656]},
     {storeUnit_maskInput_hi[28655:28640]},
     {storeUnit_maskInput_hi[28639:28624]},
     {storeUnit_maskInput_hi[28623:28608]},
     {storeUnit_maskInput_hi[28607:28592]},
     {storeUnit_maskInput_hi[28591:28576]},
     {storeUnit_maskInput_hi[28575:28560]},
     {storeUnit_maskInput_hi[28559:28544]},
     {storeUnit_maskInput_hi[28543:28528]},
     {storeUnit_maskInput_hi[28527:28512]},
     {storeUnit_maskInput_hi[28511:28496]},
     {storeUnit_maskInput_hi[28495:28480]},
     {storeUnit_maskInput_hi[28479:28464]},
     {storeUnit_maskInput_hi[28463:28448]},
     {storeUnit_maskInput_hi[28447:28432]},
     {storeUnit_maskInput_hi[28431:28416]},
     {storeUnit_maskInput_hi[28415:28400]},
     {storeUnit_maskInput_hi[28399:28384]},
     {storeUnit_maskInput_hi[28383:28368]},
     {storeUnit_maskInput_hi[28367:28352]},
     {storeUnit_maskInput_hi[28351:28336]},
     {storeUnit_maskInput_hi[28335:28320]},
     {storeUnit_maskInput_hi[28319:28304]},
     {storeUnit_maskInput_hi[28303:28288]},
     {storeUnit_maskInput_hi[28287:28272]},
     {storeUnit_maskInput_hi[28271:28256]},
     {storeUnit_maskInput_hi[28255:28240]},
     {storeUnit_maskInput_hi[28239:28224]},
     {storeUnit_maskInput_hi[28223:28208]},
     {storeUnit_maskInput_hi[28207:28192]},
     {storeUnit_maskInput_hi[28191:28176]},
     {storeUnit_maskInput_hi[28175:28160]},
     {storeUnit_maskInput_hi[28159:28144]},
     {storeUnit_maskInput_hi[28143:28128]},
     {storeUnit_maskInput_hi[28127:28112]},
     {storeUnit_maskInput_hi[28111:28096]},
     {storeUnit_maskInput_hi[28095:28080]},
     {storeUnit_maskInput_hi[28079:28064]},
     {storeUnit_maskInput_hi[28063:28048]},
     {storeUnit_maskInput_hi[28047:28032]},
     {storeUnit_maskInput_hi[28031:28016]},
     {storeUnit_maskInput_hi[28015:28000]},
     {storeUnit_maskInput_hi[27999:27984]},
     {storeUnit_maskInput_hi[27983:27968]},
     {storeUnit_maskInput_hi[27967:27952]},
     {storeUnit_maskInput_hi[27951:27936]},
     {storeUnit_maskInput_hi[27935:27920]},
     {storeUnit_maskInput_hi[27919:27904]},
     {storeUnit_maskInput_hi[27903:27888]},
     {storeUnit_maskInput_hi[27887:27872]},
     {storeUnit_maskInput_hi[27871:27856]},
     {storeUnit_maskInput_hi[27855:27840]},
     {storeUnit_maskInput_hi[27839:27824]},
     {storeUnit_maskInput_hi[27823:27808]},
     {storeUnit_maskInput_hi[27807:27792]},
     {storeUnit_maskInput_hi[27791:27776]},
     {storeUnit_maskInput_hi[27775:27760]},
     {storeUnit_maskInput_hi[27759:27744]},
     {storeUnit_maskInput_hi[27743:27728]},
     {storeUnit_maskInput_hi[27727:27712]},
     {storeUnit_maskInput_hi[27711:27696]},
     {storeUnit_maskInput_hi[27695:27680]},
     {storeUnit_maskInput_hi[27679:27664]},
     {storeUnit_maskInput_hi[27663:27648]},
     {storeUnit_maskInput_hi[27647:27632]},
     {storeUnit_maskInput_hi[27631:27616]},
     {storeUnit_maskInput_hi[27615:27600]},
     {storeUnit_maskInput_hi[27599:27584]},
     {storeUnit_maskInput_hi[27583:27568]},
     {storeUnit_maskInput_hi[27567:27552]},
     {storeUnit_maskInput_hi[27551:27536]},
     {storeUnit_maskInput_hi[27535:27520]},
     {storeUnit_maskInput_hi[27519:27504]},
     {storeUnit_maskInput_hi[27503:27488]},
     {storeUnit_maskInput_hi[27487:27472]},
     {storeUnit_maskInput_hi[27471:27456]},
     {storeUnit_maskInput_hi[27455:27440]},
     {storeUnit_maskInput_hi[27439:27424]},
     {storeUnit_maskInput_hi[27423:27408]},
     {storeUnit_maskInput_hi[27407:27392]},
     {storeUnit_maskInput_hi[27391:27376]},
     {storeUnit_maskInput_hi[27375:27360]},
     {storeUnit_maskInput_hi[27359:27344]},
     {storeUnit_maskInput_hi[27343:27328]},
     {storeUnit_maskInput_hi[27327:27312]},
     {storeUnit_maskInput_hi[27311:27296]},
     {storeUnit_maskInput_hi[27295:27280]},
     {storeUnit_maskInput_hi[27279:27264]},
     {storeUnit_maskInput_hi[27263:27248]},
     {storeUnit_maskInput_hi[27247:27232]},
     {storeUnit_maskInput_hi[27231:27216]},
     {storeUnit_maskInput_hi[27215:27200]},
     {storeUnit_maskInput_hi[27199:27184]},
     {storeUnit_maskInput_hi[27183:27168]},
     {storeUnit_maskInput_hi[27167:27152]},
     {storeUnit_maskInput_hi[27151:27136]},
     {storeUnit_maskInput_hi[27135:27120]},
     {storeUnit_maskInput_hi[27119:27104]},
     {storeUnit_maskInput_hi[27103:27088]},
     {storeUnit_maskInput_hi[27087:27072]},
     {storeUnit_maskInput_hi[27071:27056]},
     {storeUnit_maskInput_hi[27055:27040]},
     {storeUnit_maskInput_hi[27039:27024]},
     {storeUnit_maskInput_hi[27023:27008]},
     {storeUnit_maskInput_hi[27007:26992]},
     {storeUnit_maskInput_hi[26991:26976]},
     {storeUnit_maskInput_hi[26975:26960]},
     {storeUnit_maskInput_hi[26959:26944]},
     {storeUnit_maskInput_hi[26943:26928]},
     {storeUnit_maskInput_hi[26927:26912]},
     {storeUnit_maskInput_hi[26911:26896]},
     {storeUnit_maskInput_hi[26895:26880]},
     {storeUnit_maskInput_hi[26879:26864]},
     {storeUnit_maskInput_hi[26863:26848]},
     {storeUnit_maskInput_hi[26847:26832]},
     {storeUnit_maskInput_hi[26831:26816]},
     {storeUnit_maskInput_hi[26815:26800]},
     {storeUnit_maskInput_hi[26799:26784]},
     {storeUnit_maskInput_hi[26783:26768]},
     {storeUnit_maskInput_hi[26767:26752]},
     {storeUnit_maskInput_hi[26751:26736]},
     {storeUnit_maskInput_hi[26735:26720]},
     {storeUnit_maskInput_hi[26719:26704]},
     {storeUnit_maskInput_hi[26703:26688]},
     {storeUnit_maskInput_hi[26687:26672]},
     {storeUnit_maskInput_hi[26671:26656]},
     {storeUnit_maskInput_hi[26655:26640]},
     {storeUnit_maskInput_hi[26639:26624]},
     {storeUnit_maskInput_hi[26623:26608]},
     {storeUnit_maskInput_hi[26607:26592]},
     {storeUnit_maskInput_hi[26591:26576]},
     {storeUnit_maskInput_hi[26575:26560]},
     {storeUnit_maskInput_hi[26559:26544]},
     {storeUnit_maskInput_hi[26543:26528]},
     {storeUnit_maskInput_hi[26527:26512]},
     {storeUnit_maskInput_hi[26511:26496]},
     {storeUnit_maskInput_hi[26495:26480]},
     {storeUnit_maskInput_hi[26479:26464]},
     {storeUnit_maskInput_hi[26463:26448]},
     {storeUnit_maskInput_hi[26447:26432]},
     {storeUnit_maskInput_hi[26431:26416]},
     {storeUnit_maskInput_hi[26415:26400]},
     {storeUnit_maskInput_hi[26399:26384]},
     {storeUnit_maskInput_hi[26383:26368]},
     {storeUnit_maskInput_hi[26367:26352]},
     {storeUnit_maskInput_hi[26351:26336]},
     {storeUnit_maskInput_hi[26335:26320]},
     {storeUnit_maskInput_hi[26319:26304]},
     {storeUnit_maskInput_hi[26303:26288]},
     {storeUnit_maskInput_hi[26287:26272]},
     {storeUnit_maskInput_hi[26271:26256]},
     {storeUnit_maskInput_hi[26255:26240]},
     {storeUnit_maskInput_hi[26239:26224]},
     {storeUnit_maskInput_hi[26223:26208]},
     {storeUnit_maskInput_hi[26207:26192]},
     {storeUnit_maskInput_hi[26191:26176]},
     {storeUnit_maskInput_hi[26175:26160]},
     {storeUnit_maskInput_hi[26159:26144]},
     {storeUnit_maskInput_hi[26143:26128]},
     {storeUnit_maskInput_hi[26127:26112]},
     {storeUnit_maskInput_hi[26111:26096]},
     {storeUnit_maskInput_hi[26095:26080]},
     {storeUnit_maskInput_hi[26079:26064]},
     {storeUnit_maskInput_hi[26063:26048]},
     {storeUnit_maskInput_hi[26047:26032]},
     {storeUnit_maskInput_hi[26031:26016]},
     {storeUnit_maskInput_hi[26015:26000]},
     {storeUnit_maskInput_hi[25999:25984]},
     {storeUnit_maskInput_hi[25983:25968]},
     {storeUnit_maskInput_hi[25967:25952]},
     {storeUnit_maskInput_hi[25951:25936]},
     {storeUnit_maskInput_hi[25935:25920]},
     {storeUnit_maskInput_hi[25919:25904]},
     {storeUnit_maskInput_hi[25903:25888]},
     {storeUnit_maskInput_hi[25887:25872]},
     {storeUnit_maskInput_hi[25871:25856]},
     {storeUnit_maskInput_hi[25855:25840]},
     {storeUnit_maskInput_hi[25839:25824]},
     {storeUnit_maskInput_hi[25823:25808]},
     {storeUnit_maskInput_hi[25807:25792]},
     {storeUnit_maskInput_hi[25791:25776]},
     {storeUnit_maskInput_hi[25775:25760]},
     {storeUnit_maskInput_hi[25759:25744]},
     {storeUnit_maskInput_hi[25743:25728]},
     {storeUnit_maskInput_hi[25727:25712]},
     {storeUnit_maskInput_hi[25711:25696]},
     {storeUnit_maskInput_hi[25695:25680]},
     {storeUnit_maskInput_hi[25679:25664]},
     {storeUnit_maskInput_hi[25663:25648]},
     {storeUnit_maskInput_hi[25647:25632]},
     {storeUnit_maskInput_hi[25631:25616]},
     {storeUnit_maskInput_hi[25615:25600]},
     {storeUnit_maskInput_hi[25599:25584]},
     {storeUnit_maskInput_hi[25583:25568]},
     {storeUnit_maskInput_hi[25567:25552]},
     {storeUnit_maskInput_hi[25551:25536]},
     {storeUnit_maskInput_hi[25535:25520]},
     {storeUnit_maskInput_hi[25519:25504]},
     {storeUnit_maskInput_hi[25503:25488]},
     {storeUnit_maskInput_hi[25487:25472]},
     {storeUnit_maskInput_hi[25471:25456]},
     {storeUnit_maskInput_hi[25455:25440]},
     {storeUnit_maskInput_hi[25439:25424]},
     {storeUnit_maskInput_hi[25423:25408]},
     {storeUnit_maskInput_hi[25407:25392]},
     {storeUnit_maskInput_hi[25391:25376]},
     {storeUnit_maskInput_hi[25375:25360]},
     {storeUnit_maskInput_hi[25359:25344]},
     {storeUnit_maskInput_hi[25343:25328]},
     {storeUnit_maskInput_hi[25327:25312]},
     {storeUnit_maskInput_hi[25311:25296]},
     {storeUnit_maskInput_hi[25295:25280]},
     {storeUnit_maskInput_hi[25279:25264]},
     {storeUnit_maskInput_hi[25263:25248]},
     {storeUnit_maskInput_hi[25247:25232]},
     {storeUnit_maskInput_hi[25231:25216]},
     {storeUnit_maskInput_hi[25215:25200]},
     {storeUnit_maskInput_hi[25199:25184]},
     {storeUnit_maskInput_hi[25183:25168]},
     {storeUnit_maskInput_hi[25167:25152]},
     {storeUnit_maskInput_hi[25151:25136]},
     {storeUnit_maskInput_hi[25135:25120]},
     {storeUnit_maskInput_hi[25119:25104]},
     {storeUnit_maskInput_hi[25103:25088]},
     {storeUnit_maskInput_hi[25087:25072]},
     {storeUnit_maskInput_hi[25071:25056]},
     {storeUnit_maskInput_hi[25055:25040]},
     {storeUnit_maskInput_hi[25039:25024]},
     {storeUnit_maskInput_hi[25023:25008]},
     {storeUnit_maskInput_hi[25007:24992]},
     {storeUnit_maskInput_hi[24991:24976]},
     {storeUnit_maskInput_hi[24975:24960]},
     {storeUnit_maskInput_hi[24959:24944]},
     {storeUnit_maskInput_hi[24943:24928]},
     {storeUnit_maskInput_hi[24927:24912]},
     {storeUnit_maskInput_hi[24911:24896]},
     {storeUnit_maskInput_hi[24895:24880]},
     {storeUnit_maskInput_hi[24879:24864]},
     {storeUnit_maskInput_hi[24863:24848]},
     {storeUnit_maskInput_hi[24847:24832]},
     {storeUnit_maskInput_hi[24831:24816]},
     {storeUnit_maskInput_hi[24815:24800]},
     {storeUnit_maskInput_hi[24799:24784]},
     {storeUnit_maskInput_hi[24783:24768]},
     {storeUnit_maskInput_hi[24767:24752]},
     {storeUnit_maskInput_hi[24751:24736]},
     {storeUnit_maskInput_hi[24735:24720]},
     {storeUnit_maskInput_hi[24719:24704]},
     {storeUnit_maskInput_hi[24703:24688]},
     {storeUnit_maskInput_hi[24687:24672]},
     {storeUnit_maskInput_hi[24671:24656]},
     {storeUnit_maskInput_hi[24655:24640]},
     {storeUnit_maskInput_hi[24639:24624]},
     {storeUnit_maskInput_hi[24623:24608]},
     {storeUnit_maskInput_hi[24607:24592]},
     {storeUnit_maskInput_hi[24591:24576]},
     {storeUnit_maskInput_hi[24575:24560]},
     {storeUnit_maskInput_hi[24559:24544]},
     {storeUnit_maskInput_hi[24543:24528]},
     {storeUnit_maskInput_hi[24527:24512]},
     {storeUnit_maskInput_hi[24511:24496]},
     {storeUnit_maskInput_hi[24495:24480]},
     {storeUnit_maskInput_hi[24479:24464]},
     {storeUnit_maskInput_hi[24463:24448]},
     {storeUnit_maskInput_hi[24447:24432]},
     {storeUnit_maskInput_hi[24431:24416]},
     {storeUnit_maskInput_hi[24415:24400]},
     {storeUnit_maskInput_hi[24399:24384]},
     {storeUnit_maskInput_hi[24383:24368]},
     {storeUnit_maskInput_hi[24367:24352]},
     {storeUnit_maskInput_hi[24351:24336]},
     {storeUnit_maskInput_hi[24335:24320]},
     {storeUnit_maskInput_hi[24319:24304]},
     {storeUnit_maskInput_hi[24303:24288]},
     {storeUnit_maskInput_hi[24287:24272]},
     {storeUnit_maskInput_hi[24271:24256]},
     {storeUnit_maskInput_hi[24255:24240]},
     {storeUnit_maskInput_hi[24239:24224]},
     {storeUnit_maskInput_hi[24223:24208]},
     {storeUnit_maskInput_hi[24207:24192]},
     {storeUnit_maskInput_hi[24191:24176]},
     {storeUnit_maskInput_hi[24175:24160]},
     {storeUnit_maskInput_hi[24159:24144]},
     {storeUnit_maskInput_hi[24143:24128]},
     {storeUnit_maskInput_hi[24127:24112]},
     {storeUnit_maskInput_hi[24111:24096]},
     {storeUnit_maskInput_hi[24095:24080]},
     {storeUnit_maskInput_hi[24079:24064]},
     {storeUnit_maskInput_hi[24063:24048]},
     {storeUnit_maskInput_hi[24047:24032]},
     {storeUnit_maskInput_hi[24031:24016]},
     {storeUnit_maskInput_hi[24015:24000]},
     {storeUnit_maskInput_hi[23999:23984]},
     {storeUnit_maskInput_hi[23983:23968]},
     {storeUnit_maskInput_hi[23967:23952]},
     {storeUnit_maskInput_hi[23951:23936]},
     {storeUnit_maskInput_hi[23935:23920]},
     {storeUnit_maskInput_hi[23919:23904]},
     {storeUnit_maskInput_hi[23903:23888]},
     {storeUnit_maskInput_hi[23887:23872]},
     {storeUnit_maskInput_hi[23871:23856]},
     {storeUnit_maskInput_hi[23855:23840]},
     {storeUnit_maskInput_hi[23839:23824]},
     {storeUnit_maskInput_hi[23823:23808]},
     {storeUnit_maskInput_hi[23807:23792]},
     {storeUnit_maskInput_hi[23791:23776]},
     {storeUnit_maskInput_hi[23775:23760]},
     {storeUnit_maskInput_hi[23759:23744]},
     {storeUnit_maskInput_hi[23743:23728]},
     {storeUnit_maskInput_hi[23727:23712]},
     {storeUnit_maskInput_hi[23711:23696]},
     {storeUnit_maskInput_hi[23695:23680]},
     {storeUnit_maskInput_hi[23679:23664]},
     {storeUnit_maskInput_hi[23663:23648]},
     {storeUnit_maskInput_hi[23647:23632]},
     {storeUnit_maskInput_hi[23631:23616]},
     {storeUnit_maskInput_hi[23615:23600]},
     {storeUnit_maskInput_hi[23599:23584]},
     {storeUnit_maskInput_hi[23583:23568]},
     {storeUnit_maskInput_hi[23567:23552]},
     {storeUnit_maskInput_hi[23551:23536]},
     {storeUnit_maskInput_hi[23535:23520]},
     {storeUnit_maskInput_hi[23519:23504]},
     {storeUnit_maskInput_hi[23503:23488]},
     {storeUnit_maskInput_hi[23487:23472]},
     {storeUnit_maskInput_hi[23471:23456]},
     {storeUnit_maskInput_hi[23455:23440]},
     {storeUnit_maskInput_hi[23439:23424]},
     {storeUnit_maskInput_hi[23423:23408]},
     {storeUnit_maskInput_hi[23407:23392]},
     {storeUnit_maskInput_hi[23391:23376]},
     {storeUnit_maskInput_hi[23375:23360]},
     {storeUnit_maskInput_hi[23359:23344]},
     {storeUnit_maskInput_hi[23343:23328]},
     {storeUnit_maskInput_hi[23327:23312]},
     {storeUnit_maskInput_hi[23311:23296]},
     {storeUnit_maskInput_hi[23295:23280]},
     {storeUnit_maskInput_hi[23279:23264]},
     {storeUnit_maskInput_hi[23263:23248]},
     {storeUnit_maskInput_hi[23247:23232]},
     {storeUnit_maskInput_hi[23231:23216]},
     {storeUnit_maskInput_hi[23215:23200]},
     {storeUnit_maskInput_hi[23199:23184]},
     {storeUnit_maskInput_hi[23183:23168]},
     {storeUnit_maskInput_hi[23167:23152]},
     {storeUnit_maskInput_hi[23151:23136]},
     {storeUnit_maskInput_hi[23135:23120]},
     {storeUnit_maskInput_hi[23119:23104]},
     {storeUnit_maskInput_hi[23103:23088]},
     {storeUnit_maskInput_hi[23087:23072]},
     {storeUnit_maskInput_hi[23071:23056]},
     {storeUnit_maskInput_hi[23055:23040]},
     {storeUnit_maskInput_hi[23039:23024]},
     {storeUnit_maskInput_hi[23023:23008]},
     {storeUnit_maskInput_hi[23007:22992]},
     {storeUnit_maskInput_hi[22991:22976]},
     {storeUnit_maskInput_hi[22975:22960]},
     {storeUnit_maskInput_hi[22959:22944]},
     {storeUnit_maskInput_hi[22943:22928]},
     {storeUnit_maskInput_hi[22927:22912]},
     {storeUnit_maskInput_hi[22911:22896]},
     {storeUnit_maskInput_hi[22895:22880]},
     {storeUnit_maskInput_hi[22879:22864]},
     {storeUnit_maskInput_hi[22863:22848]},
     {storeUnit_maskInput_hi[22847:22832]},
     {storeUnit_maskInput_hi[22831:22816]},
     {storeUnit_maskInput_hi[22815:22800]},
     {storeUnit_maskInput_hi[22799:22784]},
     {storeUnit_maskInput_hi[22783:22768]},
     {storeUnit_maskInput_hi[22767:22752]},
     {storeUnit_maskInput_hi[22751:22736]},
     {storeUnit_maskInput_hi[22735:22720]},
     {storeUnit_maskInput_hi[22719:22704]},
     {storeUnit_maskInput_hi[22703:22688]},
     {storeUnit_maskInput_hi[22687:22672]},
     {storeUnit_maskInput_hi[22671:22656]},
     {storeUnit_maskInput_hi[22655:22640]},
     {storeUnit_maskInput_hi[22639:22624]},
     {storeUnit_maskInput_hi[22623:22608]},
     {storeUnit_maskInput_hi[22607:22592]},
     {storeUnit_maskInput_hi[22591:22576]},
     {storeUnit_maskInput_hi[22575:22560]},
     {storeUnit_maskInput_hi[22559:22544]},
     {storeUnit_maskInput_hi[22543:22528]},
     {storeUnit_maskInput_hi[22527:22512]},
     {storeUnit_maskInput_hi[22511:22496]},
     {storeUnit_maskInput_hi[22495:22480]},
     {storeUnit_maskInput_hi[22479:22464]},
     {storeUnit_maskInput_hi[22463:22448]},
     {storeUnit_maskInput_hi[22447:22432]},
     {storeUnit_maskInput_hi[22431:22416]},
     {storeUnit_maskInput_hi[22415:22400]},
     {storeUnit_maskInput_hi[22399:22384]},
     {storeUnit_maskInput_hi[22383:22368]},
     {storeUnit_maskInput_hi[22367:22352]},
     {storeUnit_maskInput_hi[22351:22336]},
     {storeUnit_maskInput_hi[22335:22320]},
     {storeUnit_maskInput_hi[22319:22304]},
     {storeUnit_maskInput_hi[22303:22288]},
     {storeUnit_maskInput_hi[22287:22272]},
     {storeUnit_maskInput_hi[22271:22256]},
     {storeUnit_maskInput_hi[22255:22240]},
     {storeUnit_maskInput_hi[22239:22224]},
     {storeUnit_maskInput_hi[22223:22208]},
     {storeUnit_maskInput_hi[22207:22192]},
     {storeUnit_maskInput_hi[22191:22176]},
     {storeUnit_maskInput_hi[22175:22160]},
     {storeUnit_maskInput_hi[22159:22144]},
     {storeUnit_maskInput_hi[22143:22128]},
     {storeUnit_maskInput_hi[22127:22112]},
     {storeUnit_maskInput_hi[22111:22096]},
     {storeUnit_maskInput_hi[22095:22080]},
     {storeUnit_maskInput_hi[22079:22064]},
     {storeUnit_maskInput_hi[22063:22048]},
     {storeUnit_maskInput_hi[22047:22032]},
     {storeUnit_maskInput_hi[22031:22016]},
     {storeUnit_maskInput_hi[22015:22000]},
     {storeUnit_maskInput_hi[21999:21984]},
     {storeUnit_maskInput_hi[21983:21968]},
     {storeUnit_maskInput_hi[21967:21952]},
     {storeUnit_maskInput_hi[21951:21936]},
     {storeUnit_maskInput_hi[21935:21920]},
     {storeUnit_maskInput_hi[21919:21904]},
     {storeUnit_maskInput_hi[21903:21888]},
     {storeUnit_maskInput_hi[21887:21872]},
     {storeUnit_maskInput_hi[21871:21856]},
     {storeUnit_maskInput_hi[21855:21840]},
     {storeUnit_maskInput_hi[21839:21824]},
     {storeUnit_maskInput_hi[21823:21808]},
     {storeUnit_maskInput_hi[21807:21792]},
     {storeUnit_maskInput_hi[21791:21776]},
     {storeUnit_maskInput_hi[21775:21760]},
     {storeUnit_maskInput_hi[21759:21744]},
     {storeUnit_maskInput_hi[21743:21728]},
     {storeUnit_maskInput_hi[21727:21712]},
     {storeUnit_maskInput_hi[21711:21696]},
     {storeUnit_maskInput_hi[21695:21680]},
     {storeUnit_maskInput_hi[21679:21664]},
     {storeUnit_maskInput_hi[21663:21648]},
     {storeUnit_maskInput_hi[21647:21632]},
     {storeUnit_maskInput_hi[21631:21616]},
     {storeUnit_maskInput_hi[21615:21600]},
     {storeUnit_maskInput_hi[21599:21584]},
     {storeUnit_maskInput_hi[21583:21568]},
     {storeUnit_maskInput_hi[21567:21552]},
     {storeUnit_maskInput_hi[21551:21536]},
     {storeUnit_maskInput_hi[21535:21520]},
     {storeUnit_maskInput_hi[21519:21504]},
     {storeUnit_maskInput_hi[21503:21488]},
     {storeUnit_maskInput_hi[21487:21472]},
     {storeUnit_maskInput_hi[21471:21456]},
     {storeUnit_maskInput_hi[21455:21440]},
     {storeUnit_maskInput_hi[21439:21424]},
     {storeUnit_maskInput_hi[21423:21408]},
     {storeUnit_maskInput_hi[21407:21392]},
     {storeUnit_maskInput_hi[21391:21376]},
     {storeUnit_maskInput_hi[21375:21360]},
     {storeUnit_maskInput_hi[21359:21344]},
     {storeUnit_maskInput_hi[21343:21328]},
     {storeUnit_maskInput_hi[21327:21312]},
     {storeUnit_maskInput_hi[21311:21296]},
     {storeUnit_maskInput_hi[21295:21280]},
     {storeUnit_maskInput_hi[21279:21264]},
     {storeUnit_maskInput_hi[21263:21248]},
     {storeUnit_maskInput_hi[21247:21232]},
     {storeUnit_maskInput_hi[21231:21216]},
     {storeUnit_maskInput_hi[21215:21200]},
     {storeUnit_maskInput_hi[21199:21184]},
     {storeUnit_maskInput_hi[21183:21168]},
     {storeUnit_maskInput_hi[21167:21152]},
     {storeUnit_maskInput_hi[21151:21136]},
     {storeUnit_maskInput_hi[21135:21120]},
     {storeUnit_maskInput_hi[21119:21104]},
     {storeUnit_maskInput_hi[21103:21088]},
     {storeUnit_maskInput_hi[21087:21072]},
     {storeUnit_maskInput_hi[21071:21056]},
     {storeUnit_maskInput_hi[21055:21040]},
     {storeUnit_maskInput_hi[21039:21024]},
     {storeUnit_maskInput_hi[21023:21008]},
     {storeUnit_maskInput_hi[21007:20992]},
     {storeUnit_maskInput_hi[20991:20976]},
     {storeUnit_maskInput_hi[20975:20960]},
     {storeUnit_maskInput_hi[20959:20944]},
     {storeUnit_maskInput_hi[20943:20928]},
     {storeUnit_maskInput_hi[20927:20912]},
     {storeUnit_maskInput_hi[20911:20896]},
     {storeUnit_maskInput_hi[20895:20880]},
     {storeUnit_maskInput_hi[20879:20864]},
     {storeUnit_maskInput_hi[20863:20848]},
     {storeUnit_maskInput_hi[20847:20832]},
     {storeUnit_maskInput_hi[20831:20816]},
     {storeUnit_maskInput_hi[20815:20800]},
     {storeUnit_maskInput_hi[20799:20784]},
     {storeUnit_maskInput_hi[20783:20768]},
     {storeUnit_maskInput_hi[20767:20752]},
     {storeUnit_maskInput_hi[20751:20736]},
     {storeUnit_maskInput_hi[20735:20720]},
     {storeUnit_maskInput_hi[20719:20704]},
     {storeUnit_maskInput_hi[20703:20688]},
     {storeUnit_maskInput_hi[20687:20672]},
     {storeUnit_maskInput_hi[20671:20656]},
     {storeUnit_maskInput_hi[20655:20640]},
     {storeUnit_maskInput_hi[20639:20624]},
     {storeUnit_maskInput_hi[20623:20608]},
     {storeUnit_maskInput_hi[20607:20592]},
     {storeUnit_maskInput_hi[20591:20576]},
     {storeUnit_maskInput_hi[20575:20560]},
     {storeUnit_maskInput_hi[20559:20544]},
     {storeUnit_maskInput_hi[20543:20528]},
     {storeUnit_maskInput_hi[20527:20512]},
     {storeUnit_maskInput_hi[20511:20496]},
     {storeUnit_maskInput_hi[20495:20480]},
     {storeUnit_maskInput_hi[20479:20464]},
     {storeUnit_maskInput_hi[20463:20448]},
     {storeUnit_maskInput_hi[20447:20432]},
     {storeUnit_maskInput_hi[20431:20416]},
     {storeUnit_maskInput_hi[20415:20400]},
     {storeUnit_maskInput_hi[20399:20384]},
     {storeUnit_maskInput_hi[20383:20368]},
     {storeUnit_maskInput_hi[20367:20352]},
     {storeUnit_maskInput_hi[20351:20336]},
     {storeUnit_maskInput_hi[20335:20320]},
     {storeUnit_maskInput_hi[20319:20304]},
     {storeUnit_maskInput_hi[20303:20288]},
     {storeUnit_maskInput_hi[20287:20272]},
     {storeUnit_maskInput_hi[20271:20256]},
     {storeUnit_maskInput_hi[20255:20240]},
     {storeUnit_maskInput_hi[20239:20224]},
     {storeUnit_maskInput_hi[20223:20208]},
     {storeUnit_maskInput_hi[20207:20192]},
     {storeUnit_maskInput_hi[20191:20176]},
     {storeUnit_maskInput_hi[20175:20160]},
     {storeUnit_maskInput_hi[20159:20144]},
     {storeUnit_maskInput_hi[20143:20128]},
     {storeUnit_maskInput_hi[20127:20112]},
     {storeUnit_maskInput_hi[20111:20096]},
     {storeUnit_maskInput_hi[20095:20080]},
     {storeUnit_maskInput_hi[20079:20064]},
     {storeUnit_maskInput_hi[20063:20048]},
     {storeUnit_maskInput_hi[20047:20032]},
     {storeUnit_maskInput_hi[20031:20016]},
     {storeUnit_maskInput_hi[20015:20000]},
     {storeUnit_maskInput_hi[19999:19984]},
     {storeUnit_maskInput_hi[19983:19968]},
     {storeUnit_maskInput_hi[19967:19952]},
     {storeUnit_maskInput_hi[19951:19936]},
     {storeUnit_maskInput_hi[19935:19920]},
     {storeUnit_maskInput_hi[19919:19904]},
     {storeUnit_maskInput_hi[19903:19888]},
     {storeUnit_maskInput_hi[19887:19872]},
     {storeUnit_maskInput_hi[19871:19856]},
     {storeUnit_maskInput_hi[19855:19840]},
     {storeUnit_maskInput_hi[19839:19824]},
     {storeUnit_maskInput_hi[19823:19808]},
     {storeUnit_maskInput_hi[19807:19792]},
     {storeUnit_maskInput_hi[19791:19776]},
     {storeUnit_maskInput_hi[19775:19760]},
     {storeUnit_maskInput_hi[19759:19744]},
     {storeUnit_maskInput_hi[19743:19728]},
     {storeUnit_maskInput_hi[19727:19712]},
     {storeUnit_maskInput_hi[19711:19696]},
     {storeUnit_maskInput_hi[19695:19680]},
     {storeUnit_maskInput_hi[19679:19664]},
     {storeUnit_maskInput_hi[19663:19648]},
     {storeUnit_maskInput_hi[19647:19632]},
     {storeUnit_maskInput_hi[19631:19616]},
     {storeUnit_maskInput_hi[19615:19600]},
     {storeUnit_maskInput_hi[19599:19584]},
     {storeUnit_maskInput_hi[19583:19568]},
     {storeUnit_maskInput_hi[19567:19552]},
     {storeUnit_maskInput_hi[19551:19536]},
     {storeUnit_maskInput_hi[19535:19520]},
     {storeUnit_maskInput_hi[19519:19504]},
     {storeUnit_maskInput_hi[19503:19488]},
     {storeUnit_maskInput_hi[19487:19472]},
     {storeUnit_maskInput_hi[19471:19456]},
     {storeUnit_maskInput_hi[19455:19440]},
     {storeUnit_maskInput_hi[19439:19424]},
     {storeUnit_maskInput_hi[19423:19408]},
     {storeUnit_maskInput_hi[19407:19392]},
     {storeUnit_maskInput_hi[19391:19376]},
     {storeUnit_maskInput_hi[19375:19360]},
     {storeUnit_maskInput_hi[19359:19344]},
     {storeUnit_maskInput_hi[19343:19328]},
     {storeUnit_maskInput_hi[19327:19312]},
     {storeUnit_maskInput_hi[19311:19296]},
     {storeUnit_maskInput_hi[19295:19280]},
     {storeUnit_maskInput_hi[19279:19264]},
     {storeUnit_maskInput_hi[19263:19248]},
     {storeUnit_maskInput_hi[19247:19232]},
     {storeUnit_maskInput_hi[19231:19216]},
     {storeUnit_maskInput_hi[19215:19200]},
     {storeUnit_maskInput_hi[19199:19184]},
     {storeUnit_maskInput_hi[19183:19168]},
     {storeUnit_maskInput_hi[19167:19152]},
     {storeUnit_maskInput_hi[19151:19136]},
     {storeUnit_maskInput_hi[19135:19120]},
     {storeUnit_maskInput_hi[19119:19104]},
     {storeUnit_maskInput_hi[19103:19088]},
     {storeUnit_maskInput_hi[19087:19072]},
     {storeUnit_maskInput_hi[19071:19056]},
     {storeUnit_maskInput_hi[19055:19040]},
     {storeUnit_maskInput_hi[19039:19024]},
     {storeUnit_maskInput_hi[19023:19008]},
     {storeUnit_maskInput_hi[19007:18992]},
     {storeUnit_maskInput_hi[18991:18976]},
     {storeUnit_maskInput_hi[18975:18960]},
     {storeUnit_maskInput_hi[18959:18944]},
     {storeUnit_maskInput_hi[18943:18928]},
     {storeUnit_maskInput_hi[18927:18912]},
     {storeUnit_maskInput_hi[18911:18896]},
     {storeUnit_maskInput_hi[18895:18880]},
     {storeUnit_maskInput_hi[18879:18864]},
     {storeUnit_maskInput_hi[18863:18848]},
     {storeUnit_maskInput_hi[18847:18832]},
     {storeUnit_maskInput_hi[18831:18816]},
     {storeUnit_maskInput_hi[18815:18800]},
     {storeUnit_maskInput_hi[18799:18784]},
     {storeUnit_maskInput_hi[18783:18768]},
     {storeUnit_maskInput_hi[18767:18752]},
     {storeUnit_maskInput_hi[18751:18736]},
     {storeUnit_maskInput_hi[18735:18720]},
     {storeUnit_maskInput_hi[18719:18704]},
     {storeUnit_maskInput_hi[18703:18688]},
     {storeUnit_maskInput_hi[18687:18672]},
     {storeUnit_maskInput_hi[18671:18656]},
     {storeUnit_maskInput_hi[18655:18640]},
     {storeUnit_maskInput_hi[18639:18624]},
     {storeUnit_maskInput_hi[18623:18608]},
     {storeUnit_maskInput_hi[18607:18592]},
     {storeUnit_maskInput_hi[18591:18576]},
     {storeUnit_maskInput_hi[18575:18560]},
     {storeUnit_maskInput_hi[18559:18544]},
     {storeUnit_maskInput_hi[18543:18528]},
     {storeUnit_maskInput_hi[18527:18512]},
     {storeUnit_maskInput_hi[18511:18496]},
     {storeUnit_maskInput_hi[18495:18480]},
     {storeUnit_maskInput_hi[18479:18464]},
     {storeUnit_maskInput_hi[18463:18448]},
     {storeUnit_maskInput_hi[18447:18432]},
     {storeUnit_maskInput_hi[18431:18416]},
     {storeUnit_maskInput_hi[18415:18400]},
     {storeUnit_maskInput_hi[18399:18384]},
     {storeUnit_maskInput_hi[18383:18368]},
     {storeUnit_maskInput_hi[18367:18352]},
     {storeUnit_maskInput_hi[18351:18336]},
     {storeUnit_maskInput_hi[18335:18320]},
     {storeUnit_maskInput_hi[18319:18304]},
     {storeUnit_maskInput_hi[18303:18288]},
     {storeUnit_maskInput_hi[18287:18272]},
     {storeUnit_maskInput_hi[18271:18256]},
     {storeUnit_maskInput_hi[18255:18240]},
     {storeUnit_maskInput_hi[18239:18224]},
     {storeUnit_maskInput_hi[18223:18208]},
     {storeUnit_maskInput_hi[18207:18192]},
     {storeUnit_maskInput_hi[18191:18176]},
     {storeUnit_maskInput_hi[18175:18160]},
     {storeUnit_maskInput_hi[18159:18144]},
     {storeUnit_maskInput_hi[18143:18128]},
     {storeUnit_maskInput_hi[18127:18112]},
     {storeUnit_maskInput_hi[18111:18096]},
     {storeUnit_maskInput_hi[18095:18080]},
     {storeUnit_maskInput_hi[18079:18064]},
     {storeUnit_maskInput_hi[18063:18048]},
     {storeUnit_maskInput_hi[18047:18032]},
     {storeUnit_maskInput_hi[18031:18016]},
     {storeUnit_maskInput_hi[18015:18000]},
     {storeUnit_maskInput_hi[17999:17984]},
     {storeUnit_maskInput_hi[17983:17968]},
     {storeUnit_maskInput_hi[17967:17952]},
     {storeUnit_maskInput_hi[17951:17936]},
     {storeUnit_maskInput_hi[17935:17920]},
     {storeUnit_maskInput_hi[17919:17904]},
     {storeUnit_maskInput_hi[17903:17888]},
     {storeUnit_maskInput_hi[17887:17872]},
     {storeUnit_maskInput_hi[17871:17856]},
     {storeUnit_maskInput_hi[17855:17840]},
     {storeUnit_maskInput_hi[17839:17824]},
     {storeUnit_maskInput_hi[17823:17808]},
     {storeUnit_maskInput_hi[17807:17792]},
     {storeUnit_maskInput_hi[17791:17776]},
     {storeUnit_maskInput_hi[17775:17760]},
     {storeUnit_maskInput_hi[17759:17744]},
     {storeUnit_maskInput_hi[17743:17728]},
     {storeUnit_maskInput_hi[17727:17712]},
     {storeUnit_maskInput_hi[17711:17696]},
     {storeUnit_maskInput_hi[17695:17680]},
     {storeUnit_maskInput_hi[17679:17664]},
     {storeUnit_maskInput_hi[17663:17648]},
     {storeUnit_maskInput_hi[17647:17632]},
     {storeUnit_maskInput_hi[17631:17616]},
     {storeUnit_maskInput_hi[17615:17600]},
     {storeUnit_maskInput_hi[17599:17584]},
     {storeUnit_maskInput_hi[17583:17568]},
     {storeUnit_maskInput_hi[17567:17552]},
     {storeUnit_maskInput_hi[17551:17536]},
     {storeUnit_maskInput_hi[17535:17520]},
     {storeUnit_maskInput_hi[17519:17504]},
     {storeUnit_maskInput_hi[17503:17488]},
     {storeUnit_maskInput_hi[17487:17472]},
     {storeUnit_maskInput_hi[17471:17456]},
     {storeUnit_maskInput_hi[17455:17440]},
     {storeUnit_maskInput_hi[17439:17424]},
     {storeUnit_maskInput_hi[17423:17408]},
     {storeUnit_maskInput_hi[17407:17392]},
     {storeUnit_maskInput_hi[17391:17376]},
     {storeUnit_maskInput_hi[17375:17360]},
     {storeUnit_maskInput_hi[17359:17344]},
     {storeUnit_maskInput_hi[17343:17328]},
     {storeUnit_maskInput_hi[17327:17312]},
     {storeUnit_maskInput_hi[17311:17296]},
     {storeUnit_maskInput_hi[17295:17280]},
     {storeUnit_maskInput_hi[17279:17264]},
     {storeUnit_maskInput_hi[17263:17248]},
     {storeUnit_maskInput_hi[17247:17232]},
     {storeUnit_maskInput_hi[17231:17216]},
     {storeUnit_maskInput_hi[17215:17200]},
     {storeUnit_maskInput_hi[17199:17184]},
     {storeUnit_maskInput_hi[17183:17168]},
     {storeUnit_maskInput_hi[17167:17152]},
     {storeUnit_maskInput_hi[17151:17136]},
     {storeUnit_maskInput_hi[17135:17120]},
     {storeUnit_maskInput_hi[17119:17104]},
     {storeUnit_maskInput_hi[17103:17088]},
     {storeUnit_maskInput_hi[17087:17072]},
     {storeUnit_maskInput_hi[17071:17056]},
     {storeUnit_maskInput_hi[17055:17040]},
     {storeUnit_maskInput_hi[17039:17024]},
     {storeUnit_maskInput_hi[17023:17008]},
     {storeUnit_maskInput_hi[17007:16992]},
     {storeUnit_maskInput_hi[16991:16976]},
     {storeUnit_maskInput_hi[16975:16960]},
     {storeUnit_maskInput_hi[16959:16944]},
     {storeUnit_maskInput_hi[16943:16928]},
     {storeUnit_maskInput_hi[16927:16912]},
     {storeUnit_maskInput_hi[16911:16896]},
     {storeUnit_maskInput_hi[16895:16880]},
     {storeUnit_maskInput_hi[16879:16864]},
     {storeUnit_maskInput_hi[16863:16848]},
     {storeUnit_maskInput_hi[16847:16832]},
     {storeUnit_maskInput_hi[16831:16816]},
     {storeUnit_maskInput_hi[16815:16800]},
     {storeUnit_maskInput_hi[16799:16784]},
     {storeUnit_maskInput_hi[16783:16768]},
     {storeUnit_maskInput_hi[16767:16752]},
     {storeUnit_maskInput_hi[16751:16736]},
     {storeUnit_maskInput_hi[16735:16720]},
     {storeUnit_maskInput_hi[16719:16704]},
     {storeUnit_maskInput_hi[16703:16688]},
     {storeUnit_maskInput_hi[16687:16672]},
     {storeUnit_maskInput_hi[16671:16656]},
     {storeUnit_maskInput_hi[16655:16640]},
     {storeUnit_maskInput_hi[16639:16624]},
     {storeUnit_maskInput_hi[16623:16608]},
     {storeUnit_maskInput_hi[16607:16592]},
     {storeUnit_maskInput_hi[16591:16576]},
     {storeUnit_maskInput_hi[16575:16560]},
     {storeUnit_maskInput_hi[16559:16544]},
     {storeUnit_maskInput_hi[16543:16528]},
     {storeUnit_maskInput_hi[16527:16512]},
     {storeUnit_maskInput_hi[16511:16496]},
     {storeUnit_maskInput_hi[16495:16480]},
     {storeUnit_maskInput_hi[16479:16464]},
     {storeUnit_maskInput_hi[16463:16448]},
     {storeUnit_maskInput_hi[16447:16432]},
     {storeUnit_maskInput_hi[16431:16416]},
     {storeUnit_maskInput_hi[16415:16400]},
     {storeUnit_maskInput_hi[16399:16384]},
     {storeUnit_maskInput_hi[16383:16368]},
     {storeUnit_maskInput_hi[16367:16352]},
     {storeUnit_maskInput_hi[16351:16336]},
     {storeUnit_maskInput_hi[16335:16320]},
     {storeUnit_maskInput_hi[16319:16304]},
     {storeUnit_maskInput_hi[16303:16288]},
     {storeUnit_maskInput_hi[16287:16272]},
     {storeUnit_maskInput_hi[16271:16256]},
     {storeUnit_maskInput_hi[16255:16240]},
     {storeUnit_maskInput_hi[16239:16224]},
     {storeUnit_maskInput_hi[16223:16208]},
     {storeUnit_maskInput_hi[16207:16192]},
     {storeUnit_maskInput_hi[16191:16176]},
     {storeUnit_maskInput_hi[16175:16160]},
     {storeUnit_maskInput_hi[16159:16144]},
     {storeUnit_maskInput_hi[16143:16128]},
     {storeUnit_maskInput_hi[16127:16112]},
     {storeUnit_maskInput_hi[16111:16096]},
     {storeUnit_maskInput_hi[16095:16080]},
     {storeUnit_maskInput_hi[16079:16064]},
     {storeUnit_maskInput_hi[16063:16048]},
     {storeUnit_maskInput_hi[16047:16032]},
     {storeUnit_maskInput_hi[16031:16016]},
     {storeUnit_maskInput_hi[16015:16000]},
     {storeUnit_maskInput_hi[15999:15984]},
     {storeUnit_maskInput_hi[15983:15968]},
     {storeUnit_maskInput_hi[15967:15952]},
     {storeUnit_maskInput_hi[15951:15936]},
     {storeUnit_maskInput_hi[15935:15920]},
     {storeUnit_maskInput_hi[15919:15904]},
     {storeUnit_maskInput_hi[15903:15888]},
     {storeUnit_maskInput_hi[15887:15872]},
     {storeUnit_maskInput_hi[15871:15856]},
     {storeUnit_maskInput_hi[15855:15840]},
     {storeUnit_maskInput_hi[15839:15824]},
     {storeUnit_maskInput_hi[15823:15808]},
     {storeUnit_maskInput_hi[15807:15792]},
     {storeUnit_maskInput_hi[15791:15776]},
     {storeUnit_maskInput_hi[15775:15760]},
     {storeUnit_maskInput_hi[15759:15744]},
     {storeUnit_maskInput_hi[15743:15728]},
     {storeUnit_maskInput_hi[15727:15712]},
     {storeUnit_maskInput_hi[15711:15696]},
     {storeUnit_maskInput_hi[15695:15680]},
     {storeUnit_maskInput_hi[15679:15664]},
     {storeUnit_maskInput_hi[15663:15648]},
     {storeUnit_maskInput_hi[15647:15632]},
     {storeUnit_maskInput_hi[15631:15616]},
     {storeUnit_maskInput_hi[15615:15600]},
     {storeUnit_maskInput_hi[15599:15584]},
     {storeUnit_maskInput_hi[15583:15568]},
     {storeUnit_maskInput_hi[15567:15552]},
     {storeUnit_maskInput_hi[15551:15536]},
     {storeUnit_maskInput_hi[15535:15520]},
     {storeUnit_maskInput_hi[15519:15504]},
     {storeUnit_maskInput_hi[15503:15488]},
     {storeUnit_maskInput_hi[15487:15472]},
     {storeUnit_maskInput_hi[15471:15456]},
     {storeUnit_maskInput_hi[15455:15440]},
     {storeUnit_maskInput_hi[15439:15424]},
     {storeUnit_maskInput_hi[15423:15408]},
     {storeUnit_maskInput_hi[15407:15392]},
     {storeUnit_maskInput_hi[15391:15376]},
     {storeUnit_maskInput_hi[15375:15360]},
     {storeUnit_maskInput_hi[15359:15344]},
     {storeUnit_maskInput_hi[15343:15328]},
     {storeUnit_maskInput_hi[15327:15312]},
     {storeUnit_maskInput_hi[15311:15296]},
     {storeUnit_maskInput_hi[15295:15280]},
     {storeUnit_maskInput_hi[15279:15264]},
     {storeUnit_maskInput_hi[15263:15248]},
     {storeUnit_maskInput_hi[15247:15232]},
     {storeUnit_maskInput_hi[15231:15216]},
     {storeUnit_maskInput_hi[15215:15200]},
     {storeUnit_maskInput_hi[15199:15184]},
     {storeUnit_maskInput_hi[15183:15168]},
     {storeUnit_maskInput_hi[15167:15152]},
     {storeUnit_maskInput_hi[15151:15136]},
     {storeUnit_maskInput_hi[15135:15120]},
     {storeUnit_maskInput_hi[15119:15104]},
     {storeUnit_maskInput_hi[15103:15088]},
     {storeUnit_maskInput_hi[15087:15072]},
     {storeUnit_maskInput_hi[15071:15056]},
     {storeUnit_maskInput_hi[15055:15040]},
     {storeUnit_maskInput_hi[15039:15024]},
     {storeUnit_maskInput_hi[15023:15008]},
     {storeUnit_maskInput_hi[15007:14992]},
     {storeUnit_maskInput_hi[14991:14976]},
     {storeUnit_maskInput_hi[14975:14960]},
     {storeUnit_maskInput_hi[14959:14944]},
     {storeUnit_maskInput_hi[14943:14928]},
     {storeUnit_maskInput_hi[14927:14912]},
     {storeUnit_maskInput_hi[14911:14896]},
     {storeUnit_maskInput_hi[14895:14880]},
     {storeUnit_maskInput_hi[14879:14864]},
     {storeUnit_maskInput_hi[14863:14848]},
     {storeUnit_maskInput_hi[14847:14832]},
     {storeUnit_maskInput_hi[14831:14816]},
     {storeUnit_maskInput_hi[14815:14800]},
     {storeUnit_maskInput_hi[14799:14784]},
     {storeUnit_maskInput_hi[14783:14768]},
     {storeUnit_maskInput_hi[14767:14752]},
     {storeUnit_maskInput_hi[14751:14736]},
     {storeUnit_maskInput_hi[14735:14720]},
     {storeUnit_maskInput_hi[14719:14704]},
     {storeUnit_maskInput_hi[14703:14688]},
     {storeUnit_maskInput_hi[14687:14672]},
     {storeUnit_maskInput_hi[14671:14656]},
     {storeUnit_maskInput_hi[14655:14640]},
     {storeUnit_maskInput_hi[14639:14624]},
     {storeUnit_maskInput_hi[14623:14608]},
     {storeUnit_maskInput_hi[14607:14592]},
     {storeUnit_maskInput_hi[14591:14576]},
     {storeUnit_maskInput_hi[14575:14560]},
     {storeUnit_maskInput_hi[14559:14544]},
     {storeUnit_maskInput_hi[14543:14528]},
     {storeUnit_maskInput_hi[14527:14512]},
     {storeUnit_maskInput_hi[14511:14496]},
     {storeUnit_maskInput_hi[14495:14480]},
     {storeUnit_maskInput_hi[14479:14464]},
     {storeUnit_maskInput_hi[14463:14448]},
     {storeUnit_maskInput_hi[14447:14432]},
     {storeUnit_maskInput_hi[14431:14416]},
     {storeUnit_maskInput_hi[14415:14400]},
     {storeUnit_maskInput_hi[14399:14384]},
     {storeUnit_maskInput_hi[14383:14368]},
     {storeUnit_maskInput_hi[14367:14352]},
     {storeUnit_maskInput_hi[14351:14336]},
     {storeUnit_maskInput_hi[14335:14320]},
     {storeUnit_maskInput_hi[14319:14304]},
     {storeUnit_maskInput_hi[14303:14288]},
     {storeUnit_maskInput_hi[14287:14272]},
     {storeUnit_maskInput_hi[14271:14256]},
     {storeUnit_maskInput_hi[14255:14240]},
     {storeUnit_maskInput_hi[14239:14224]},
     {storeUnit_maskInput_hi[14223:14208]},
     {storeUnit_maskInput_hi[14207:14192]},
     {storeUnit_maskInput_hi[14191:14176]},
     {storeUnit_maskInput_hi[14175:14160]},
     {storeUnit_maskInput_hi[14159:14144]},
     {storeUnit_maskInput_hi[14143:14128]},
     {storeUnit_maskInput_hi[14127:14112]},
     {storeUnit_maskInput_hi[14111:14096]},
     {storeUnit_maskInput_hi[14095:14080]},
     {storeUnit_maskInput_hi[14079:14064]},
     {storeUnit_maskInput_hi[14063:14048]},
     {storeUnit_maskInput_hi[14047:14032]},
     {storeUnit_maskInput_hi[14031:14016]},
     {storeUnit_maskInput_hi[14015:14000]},
     {storeUnit_maskInput_hi[13999:13984]},
     {storeUnit_maskInput_hi[13983:13968]},
     {storeUnit_maskInput_hi[13967:13952]},
     {storeUnit_maskInput_hi[13951:13936]},
     {storeUnit_maskInput_hi[13935:13920]},
     {storeUnit_maskInput_hi[13919:13904]},
     {storeUnit_maskInput_hi[13903:13888]},
     {storeUnit_maskInput_hi[13887:13872]},
     {storeUnit_maskInput_hi[13871:13856]},
     {storeUnit_maskInput_hi[13855:13840]},
     {storeUnit_maskInput_hi[13839:13824]},
     {storeUnit_maskInput_hi[13823:13808]},
     {storeUnit_maskInput_hi[13807:13792]},
     {storeUnit_maskInput_hi[13791:13776]},
     {storeUnit_maskInput_hi[13775:13760]},
     {storeUnit_maskInput_hi[13759:13744]},
     {storeUnit_maskInput_hi[13743:13728]},
     {storeUnit_maskInput_hi[13727:13712]},
     {storeUnit_maskInput_hi[13711:13696]},
     {storeUnit_maskInput_hi[13695:13680]},
     {storeUnit_maskInput_hi[13679:13664]},
     {storeUnit_maskInput_hi[13663:13648]},
     {storeUnit_maskInput_hi[13647:13632]},
     {storeUnit_maskInput_hi[13631:13616]},
     {storeUnit_maskInput_hi[13615:13600]},
     {storeUnit_maskInput_hi[13599:13584]},
     {storeUnit_maskInput_hi[13583:13568]},
     {storeUnit_maskInput_hi[13567:13552]},
     {storeUnit_maskInput_hi[13551:13536]},
     {storeUnit_maskInput_hi[13535:13520]},
     {storeUnit_maskInput_hi[13519:13504]},
     {storeUnit_maskInput_hi[13503:13488]},
     {storeUnit_maskInput_hi[13487:13472]},
     {storeUnit_maskInput_hi[13471:13456]},
     {storeUnit_maskInput_hi[13455:13440]},
     {storeUnit_maskInput_hi[13439:13424]},
     {storeUnit_maskInput_hi[13423:13408]},
     {storeUnit_maskInput_hi[13407:13392]},
     {storeUnit_maskInput_hi[13391:13376]},
     {storeUnit_maskInput_hi[13375:13360]},
     {storeUnit_maskInput_hi[13359:13344]},
     {storeUnit_maskInput_hi[13343:13328]},
     {storeUnit_maskInput_hi[13327:13312]},
     {storeUnit_maskInput_hi[13311:13296]},
     {storeUnit_maskInput_hi[13295:13280]},
     {storeUnit_maskInput_hi[13279:13264]},
     {storeUnit_maskInput_hi[13263:13248]},
     {storeUnit_maskInput_hi[13247:13232]},
     {storeUnit_maskInput_hi[13231:13216]},
     {storeUnit_maskInput_hi[13215:13200]},
     {storeUnit_maskInput_hi[13199:13184]},
     {storeUnit_maskInput_hi[13183:13168]},
     {storeUnit_maskInput_hi[13167:13152]},
     {storeUnit_maskInput_hi[13151:13136]},
     {storeUnit_maskInput_hi[13135:13120]},
     {storeUnit_maskInput_hi[13119:13104]},
     {storeUnit_maskInput_hi[13103:13088]},
     {storeUnit_maskInput_hi[13087:13072]},
     {storeUnit_maskInput_hi[13071:13056]},
     {storeUnit_maskInput_hi[13055:13040]},
     {storeUnit_maskInput_hi[13039:13024]},
     {storeUnit_maskInput_hi[13023:13008]},
     {storeUnit_maskInput_hi[13007:12992]},
     {storeUnit_maskInput_hi[12991:12976]},
     {storeUnit_maskInput_hi[12975:12960]},
     {storeUnit_maskInput_hi[12959:12944]},
     {storeUnit_maskInput_hi[12943:12928]},
     {storeUnit_maskInput_hi[12927:12912]},
     {storeUnit_maskInput_hi[12911:12896]},
     {storeUnit_maskInput_hi[12895:12880]},
     {storeUnit_maskInput_hi[12879:12864]},
     {storeUnit_maskInput_hi[12863:12848]},
     {storeUnit_maskInput_hi[12847:12832]},
     {storeUnit_maskInput_hi[12831:12816]},
     {storeUnit_maskInput_hi[12815:12800]},
     {storeUnit_maskInput_hi[12799:12784]},
     {storeUnit_maskInput_hi[12783:12768]},
     {storeUnit_maskInput_hi[12767:12752]},
     {storeUnit_maskInput_hi[12751:12736]},
     {storeUnit_maskInput_hi[12735:12720]},
     {storeUnit_maskInput_hi[12719:12704]},
     {storeUnit_maskInput_hi[12703:12688]},
     {storeUnit_maskInput_hi[12687:12672]},
     {storeUnit_maskInput_hi[12671:12656]},
     {storeUnit_maskInput_hi[12655:12640]},
     {storeUnit_maskInput_hi[12639:12624]},
     {storeUnit_maskInput_hi[12623:12608]},
     {storeUnit_maskInput_hi[12607:12592]},
     {storeUnit_maskInput_hi[12591:12576]},
     {storeUnit_maskInput_hi[12575:12560]},
     {storeUnit_maskInput_hi[12559:12544]},
     {storeUnit_maskInput_hi[12543:12528]},
     {storeUnit_maskInput_hi[12527:12512]},
     {storeUnit_maskInput_hi[12511:12496]},
     {storeUnit_maskInput_hi[12495:12480]},
     {storeUnit_maskInput_hi[12479:12464]},
     {storeUnit_maskInput_hi[12463:12448]},
     {storeUnit_maskInput_hi[12447:12432]},
     {storeUnit_maskInput_hi[12431:12416]},
     {storeUnit_maskInput_hi[12415:12400]},
     {storeUnit_maskInput_hi[12399:12384]},
     {storeUnit_maskInput_hi[12383:12368]},
     {storeUnit_maskInput_hi[12367:12352]},
     {storeUnit_maskInput_hi[12351:12336]},
     {storeUnit_maskInput_hi[12335:12320]},
     {storeUnit_maskInput_hi[12319:12304]},
     {storeUnit_maskInput_hi[12303:12288]},
     {storeUnit_maskInput_hi[12287:12272]},
     {storeUnit_maskInput_hi[12271:12256]},
     {storeUnit_maskInput_hi[12255:12240]},
     {storeUnit_maskInput_hi[12239:12224]},
     {storeUnit_maskInput_hi[12223:12208]},
     {storeUnit_maskInput_hi[12207:12192]},
     {storeUnit_maskInput_hi[12191:12176]},
     {storeUnit_maskInput_hi[12175:12160]},
     {storeUnit_maskInput_hi[12159:12144]},
     {storeUnit_maskInput_hi[12143:12128]},
     {storeUnit_maskInput_hi[12127:12112]},
     {storeUnit_maskInput_hi[12111:12096]},
     {storeUnit_maskInput_hi[12095:12080]},
     {storeUnit_maskInput_hi[12079:12064]},
     {storeUnit_maskInput_hi[12063:12048]},
     {storeUnit_maskInput_hi[12047:12032]},
     {storeUnit_maskInput_hi[12031:12016]},
     {storeUnit_maskInput_hi[12015:12000]},
     {storeUnit_maskInput_hi[11999:11984]},
     {storeUnit_maskInput_hi[11983:11968]},
     {storeUnit_maskInput_hi[11967:11952]},
     {storeUnit_maskInput_hi[11951:11936]},
     {storeUnit_maskInput_hi[11935:11920]},
     {storeUnit_maskInput_hi[11919:11904]},
     {storeUnit_maskInput_hi[11903:11888]},
     {storeUnit_maskInput_hi[11887:11872]},
     {storeUnit_maskInput_hi[11871:11856]},
     {storeUnit_maskInput_hi[11855:11840]},
     {storeUnit_maskInput_hi[11839:11824]},
     {storeUnit_maskInput_hi[11823:11808]},
     {storeUnit_maskInput_hi[11807:11792]},
     {storeUnit_maskInput_hi[11791:11776]},
     {storeUnit_maskInput_hi[11775:11760]},
     {storeUnit_maskInput_hi[11759:11744]},
     {storeUnit_maskInput_hi[11743:11728]},
     {storeUnit_maskInput_hi[11727:11712]},
     {storeUnit_maskInput_hi[11711:11696]},
     {storeUnit_maskInput_hi[11695:11680]},
     {storeUnit_maskInput_hi[11679:11664]},
     {storeUnit_maskInput_hi[11663:11648]},
     {storeUnit_maskInput_hi[11647:11632]},
     {storeUnit_maskInput_hi[11631:11616]},
     {storeUnit_maskInput_hi[11615:11600]},
     {storeUnit_maskInput_hi[11599:11584]},
     {storeUnit_maskInput_hi[11583:11568]},
     {storeUnit_maskInput_hi[11567:11552]},
     {storeUnit_maskInput_hi[11551:11536]},
     {storeUnit_maskInput_hi[11535:11520]},
     {storeUnit_maskInput_hi[11519:11504]},
     {storeUnit_maskInput_hi[11503:11488]},
     {storeUnit_maskInput_hi[11487:11472]},
     {storeUnit_maskInput_hi[11471:11456]},
     {storeUnit_maskInput_hi[11455:11440]},
     {storeUnit_maskInput_hi[11439:11424]},
     {storeUnit_maskInput_hi[11423:11408]},
     {storeUnit_maskInput_hi[11407:11392]},
     {storeUnit_maskInput_hi[11391:11376]},
     {storeUnit_maskInput_hi[11375:11360]},
     {storeUnit_maskInput_hi[11359:11344]},
     {storeUnit_maskInput_hi[11343:11328]},
     {storeUnit_maskInput_hi[11327:11312]},
     {storeUnit_maskInput_hi[11311:11296]},
     {storeUnit_maskInput_hi[11295:11280]},
     {storeUnit_maskInput_hi[11279:11264]},
     {storeUnit_maskInput_hi[11263:11248]},
     {storeUnit_maskInput_hi[11247:11232]},
     {storeUnit_maskInput_hi[11231:11216]},
     {storeUnit_maskInput_hi[11215:11200]},
     {storeUnit_maskInput_hi[11199:11184]},
     {storeUnit_maskInput_hi[11183:11168]},
     {storeUnit_maskInput_hi[11167:11152]},
     {storeUnit_maskInput_hi[11151:11136]},
     {storeUnit_maskInput_hi[11135:11120]},
     {storeUnit_maskInput_hi[11119:11104]},
     {storeUnit_maskInput_hi[11103:11088]},
     {storeUnit_maskInput_hi[11087:11072]},
     {storeUnit_maskInput_hi[11071:11056]},
     {storeUnit_maskInput_hi[11055:11040]},
     {storeUnit_maskInput_hi[11039:11024]},
     {storeUnit_maskInput_hi[11023:11008]},
     {storeUnit_maskInput_hi[11007:10992]},
     {storeUnit_maskInput_hi[10991:10976]},
     {storeUnit_maskInput_hi[10975:10960]},
     {storeUnit_maskInput_hi[10959:10944]},
     {storeUnit_maskInput_hi[10943:10928]},
     {storeUnit_maskInput_hi[10927:10912]},
     {storeUnit_maskInput_hi[10911:10896]},
     {storeUnit_maskInput_hi[10895:10880]},
     {storeUnit_maskInput_hi[10879:10864]},
     {storeUnit_maskInput_hi[10863:10848]},
     {storeUnit_maskInput_hi[10847:10832]},
     {storeUnit_maskInput_hi[10831:10816]},
     {storeUnit_maskInput_hi[10815:10800]},
     {storeUnit_maskInput_hi[10799:10784]},
     {storeUnit_maskInput_hi[10783:10768]},
     {storeUnit_maskInput_hi[10767:10752]},
     {storeUnit_maskInput_hi[10751:10736]},
     {storeUnit_maskInput_hi[10735:10720]},
     {storeUnit_maskInput_hi[10719:10704]},
     {storeUnit_maskInput_hi[10703:10688]},
     {storeUnit_maskInput_hi[10687:10672]},
     {storeUnit_maskInput_hi[10671:10656]},
     {storeUnit_maskInput_hi[10655:10640]},
     {storeUnit_maskInput_hi[10639:10624]},
     {storeUnit_maskInput_hi[10623:10608]},
     {storeUnit_maskInput_hi[10607:10592]},
     {storeUnit_maskInput_hi[10591:10576]},
     {storeUnit_maskInput_hi[10575:10560]},
     {storeUnit_maskInput_hi[10559:10544]},
     {storeUnit_maskInput_hi[10543:10528]},
     {storeUnit_maskInput_hi[10527:10512]},
     {storeUnit_maskInput_hi[10511:10496]},
     {storeUnit_maskInput_hi[10495:10480]},
     {storeUnit_maskInput_hi[10479:10464]},
     {storeUnit_maskInput_hi[10463:10448]},
     {storeUnit_maskInput_hi[10447:10432]},
     {storeUnit_maskInput_hi[10431:10416]},
     {storeUnit_maskInput_hi[10415:10400]},
     {storeUnit_maskInput_hi[10399:10384]},
     {storeUnit_maskInput_hi[10383:10368]},
     {storeUnit_maskInput_hi[10367:10352]},
     {storeUnit_maskInput_hi[10351:10336]},
     {storeUnit_maskInput_hi[10335:10320]},
     {storeUnit_maskInput_hi[10319:10304]},
     {storeUnit_maskInput_hi[10303:10288]},
     {storeUnit_maskInput_hi[10287:10272]},
     {storeUnit_maskInput_hi[10271:10256]},
     {storeUnit_maskInput_hi[10255:10240]},
     {storeUnit_maskInput_hi[10239:10224]},
     {storeUnit_maskInput_hi[10223:10208]},
     {storeUnit_maskInput_hi[10207:10192]},
     {storeUnit_maskInput_hi[10191:10176]},
     {storeUnit_maskInput_hi[10175:10160]},
     {storeUnit_maskInput_hi[10159:10144]},
     {storeUnit_maskInput_hi[10143:10128]},
     {storeUnit_maskInput_hi[10127:10112]},
     {storeUnit_maskInput_hi[10111:10096]},
     {storeUnit_maskInput_hi[10095:10080]},
     {storeUnit_maskInput_hi[10079:10064]},
     {storeUnit_maskInput_hi[10063:10048]},
     {storeUnit_maskInput_hi[10047:10032]},
     {storeUnit_maskInput_hi[10031:10016]},
     {storeUnit_maskInput_hi[10015:10000]},
     {storeUnit_maskInput_hi[9999:9984]},
     {storeUnit_maskInput_hi[9983:9968]},
     {storeUnit_maskInput_hi[9967:9952]},
     {storeUnit_maskInput_hi[9951:9936]},
     {storeUnit_maskInput_hi[9935:9920]},
     {storeUnit_maskInput_hi[9919:9904]},
     {storeUnit_maskInput_hi[9903:9888]},
     {storeUnit_maskInput_hi[9887:9872]},
     {storeUnit_maskInput_hi[9871:9856]},
     {storeUnit_maskInput_hi[9855:9840]},
     {storeUnit_maskInput_hi[9839:9824]},
     {storeUnit_maskInput_hi[9823:9808]},
     {storeUnit_maskInput_hi[9807:9792]},
     {storeUnit_maskInput_hi[9791:9776]},
     {storeUnit_maskInput_hi[9775:9760]},
     {storeUnit_maskInput_hi[9759:9744]},
     {storeUnit_maskInput_hi[9743:9728]},
     {storeUnit_maskInput_hi[9727:9712]},
     {storeUnit_maskInput_hi[9711:9696]},
     {storeUnit_maskInput_hi[9695:9680]},
     {storeUnit_maskInput_hi[9679:9664]},
     {storeUnit_maskInput_hi[9663:9648]},
     {storeUnit_maskInput_hi[9647:9632]},
     {storeUnit_maskInput_hi[9631:9616]},
     {storeUnit_maskInput_hi[9615:9600]},
     {storeUnit_maskInput_hi[9599:9584]},
     {storeUnit_maskInput_hi[9583:9568]},
     {storeUnit_maskInput_hi[9567:9552]},
     {storeUnit_maskInput_hi[9551:9536]},
     {storeUnit_maskInput_hi[9535:9520]},
     {storeUnit_maskInput_hi[9519:9504]},
     {storeUnit_maskInput_hi[9503:9488]},
     {storeUnit_maskInput_hi[9487:9472]},
     {storeUnit_maskInput_hi[9471:9456]},
     {storeUnit_maskInput_hi[9455:9440]},
     {storeUnit_maskInput_hi[9439:9424]},
     {storeUnit_maskInput_hi[9423:9408]},
     {storeUnit_maskInput_hi[9407:9392]},
     {storeUnit_maskInput_hi[9391:9376]},
     {storeUnit_maskInput_hi[9375:9360]},
     {storeUnit_maskInput_hi[9359:9344]},
     {storeUnit_maskInput_hi[9343:9328]},
     {storeUnit_maskInput_hi[9327:9312]},
     {storeUnit_maskInput_hi[9311:9296]},
     {storeUnit_maskInput_hi[9295:9280]},
     {storeUnit_maskInput_hi[9279:9264]},
     {storeUnit_maskInput_hi[9263:9248]},
     {storeUnit_maskInput_hi[9247:9232]},
     {storeUnit_maskInput_hi[9231:9216]},
     {storeUnit_maskInput_hi[9215:9200]},
     {storeUnit_maskInput_hi[9199:9184]},
     {storeUnit_maskInput_hi[9183:9168]},
     {storeUnit_maskInput_hi[9167:9152]},
     {storeUnit_maskInput_hi[9151:9136]},
     {storeUnit_maskInput_hi[9135:9120]},
     {storeUnit_maskInput_hi[9119:9104]},
     {storeUnit_maskInput_hi[9103:9088]},
     {storeUnit_maskInput_hi[9087:9072]},
     {storeUnit_maskInput_hi[9071:9056]},
     {storeUnit_maskInput_hi[9055:9040]},
     {storeUnit_maskInput_hi[9039:9024]},
     {storeUnit_maskInput_hi[9023:9008]},
     {storeUnit_maskInput_hi[9007:8992]},
     {storeUnit_maskInput_hi[8991:8976]},
     {storeUnit_maskInput_hi[8975:8960]},
     {storeUnit_maskInput_hi[8959:8944]},
     {storeUnit_maskInput_hi[8943:8928]},
     {storeUnit_maskInput_hi[8927:8912]},
     {storeUnit_maskInput_hi[8911:8896]},
     {storeUnit_maskInput_hi[8895:8880]},
     {storeUnit_maskInput_hi[8879:8864]},
     {storeUnit_maskInput_hi[8863:8848]},
     {storeUnit_maskInput_hi[8847:8832]},
     {storeUnit_maskInput_hi[8831:8816]},
     {storeUnit_maskInput_hi[8815:8800]},
     {storeUnit_maskInput_hi[8799:8784]},
     {storeUnit_maskInput_hi[8783:8768]},
     {storeUnit_maskInput_hi[8767:8752]},
     {storeUnit_maskInput_hi[8751:8736]},
     {storeUnit_maskInput_hi[8735:8720]},
     {storeUnit_maskInput_hi[8719:8704]},
     {storeUnit_maskInput_hi[8703:8688]},
     {storeUnit_maskInput_hi[8687:8672]},
     {storeUnit_maskInput_hi[8671:8656]},
     {storeUnit_maskInput_hi[8655:8640]},
     {storeUnit_maskInput_hi[8639:8624]},
     {storeUnit_maskInput_hi[8623:8608]},
     {storeUnit_maskInput_hi[8607:8592]},
     {storeUnit_maskInput_hi[8591:8576]},
     {storeUnit_maskInput_hi[8575:8560]},
     {storeUnit_maskInput_hi[8559:8544]},
     {storeUnit_maskInput_hi[8543:8528]},
     {storeUnit_maskInput_hi[8527:8512]},
     {storeUnit_maskInput_hi[8511:8496]},
     {storeUnit_maskInput_hi[8495:8480]},
     {storeUnit_maskInput_hi[8479:8464]},
     {storeUnit_maskInput_hi[8463:8448]},
     {storeUnit_maskInput_hi[8447:8432]},
     {storeUnit_maskInput_hi[8431:8416]},
     {storeUnit_maskInput_hi[8415:8400]},
     {storeUnit_maskInput_hi[8399:8384]},
     {storeUnit_maskInput_hi[8383:8368]},
     {storeUnit_maskInput_hi[8367:8352]},
     {storeUnit_maskInput_hi[8351:8336]},
     {storeUnit_maskInput_hi[8335:8320]},
     {storeUnit_maskInput_hi[8319:8304]},
     {storeUnit_maskInput_hi[8303:8288]},
     {storeUnit_maskInput_hi[8287:8272]},
     {storeUnit_maskInput_hi[8271:8256]},
     {storeUnit_maskInput_hi[8255:8240]},
     {storeUnit_maskInput_hi[8239:8224]},
     {storeUnit_maskInput_hi[8223:8208]},
     {storeUnit_maskInput_hi[8207:8192]},
     {storeUnit_maskInput_hi[8191:8176]},
     {storeUnit_maskInput_hi[8175:8160]},
     {storeUnit_maskInput_hi[8159:8144]},
     {storeUnit_maskInput_hi[8143:8128]},
     {storeUnit_maskInput_hi[8127:8112]},
     {storeUnit_maskInput_hi[8111:8096]},
     {storeUnit_maskInput_hi[8095:8080]},
     {storeUnit_maskInput_hi[8079:8064]},
     {storeUnit_maskInput_hi[8063:8048]},
     {storeUnit_maskInput_hi[8047:8032]},
     {storeUnit_maskInput_hi[8031:8016]},
     {storeUnit_maskInput_hi[8015:8000]},
     {storeUnit_maskInput_hi[7999:7984]},
     {storeUnit_maskInput_hi[7983:7968]},
     {storeUnit_maskInput_hi[7967:7952]},
     {storeUnit_maskInput_hi[7951:7936]},
     {storeUnit_maskInput_hi[7935:7920]},
     {storeUnit_maskInput_hi[7919:7904]},
     {storeUnit_maskInput_hi[7903:7888]},
     {storeUnit_maskInput_hi[7887:7872]},
     {storeUnit_maskInput_hi[7871:7856]},
     {storeUnit_maskInput_hi[7855:7840]},
     {storeUnit_maskInput_hi[7839:7824]},
     {storeUnit_maskInput_hi[7823:7808]},
     {storeUnit_maskInput_hi[7807:7792]},
     {storeUnit_maskInput_hi[7791:7776]},
     {storeUnit_maskInput_hi[7775:7760]},
     {storeUnit_maskInput_hi[7759:7744]},
     {storeUnit_maskInput_hi[7743:7728]},
     {storeUnit_maskInput_hi[7727:7712]},
     {storeUnit_maskInput_hi[7711:7696]},
     {storeUnit_maskInput_hi[7695:7680]},
     {storeUnit_maskInput_hi[7679:7664]},
     {storeUnit_maskInput_hi[7663:7648]},
     {storeUnit_maskInput_hi[7647:7632]},
     {storeUnit_maskInput_hi[7631:7616]},
     {storeUnit_maskInput_hi[7615:7600]},
     {storeUnit_maskInput_hi[7599:7584]},
     {storeUnit_maskInput_hi[7583:7568]},
     {storeUnit_maskInput_hi[7567:7552]},
     {storeUnit_maskInput_hi[7551:7536]},
     {storeUnit_maskInput_hi[7535:7520]},
     {storeUnit_maskInput_hi[7519:7504]},
     {storeUnit_maskInput_hi[7503:7488]},
     {storeUnit_maskInput_hi[7487:7472]},
     {storeUnit_maskInput_hi[7471:7456]},
     {storeUnit_maskInput_hi[7455:7440]},
     {storeUnit_maskInput_hi[7439:7424]},
     {storeUnit_maskInput_hi[7423:7408]},
     {storeUnit_maskInput_hi[7407:7392]},
     {storeUnit_maskInput_hi[7391:7376]},
     {storeUnit_maskInput_hi[7375:7360]},
     {storeUnit_maskInput_hi[7359:7344]},
     {storeUnit_maskInput_hi[7343:7328]},
     {storeUnit_maskInput_hi[7327:7312]},
     {storeUnit_maskInput_hi[7311:7296]},
     {storeUnit_maskInput_hi[7295:7280]},
     {storeUnit_maskInput_hi[7279:7264]},
     {storeUnit_maskInput_hi[7263:7248]},
     {storeUnit_maskInput_hi[7247:7232]},
     {storeUnit_maskInput_hi[7231:7216]},
     {storeUnit_maskInput_hi[7215:7200]},
     {storeUnit_maskInput_hi[7199:7184]},
     {storeUnit_maskInput_hi[7183:7168]},
     {storeUnit_maskInput_hi[7167:7152]},
     {storeUnit_maskInput_hi[7151:7136]},
     {storeUnit_maskInput_hi[7135:7120]},
     {storeUnit_maskInput_hi[7119:7104]},
     {storeUnit_maskInput_hi[7103:7088]},
     {storeUnit_maskInput_hi[7087:7072]},
     {storeUnit_maskInput_hi[7071:7056]},
     {storeUnit_maskInput_hi[7055:7040]},
     {storeUnit_maskInput_hi[7039:7024]},
     {storeUnit_maskInput_hi[7023:7008]},
     {storeUnit_maskInput_hi[7007:6992]},
     {storeUnit_maskInput_hi[6991:6976]},
     {storeUnit_maskInput_hi[6975:6960]},
     {storeUnit_maskInput_hi[6959:6944]},
     {storeUnit_maskInput_hi[6943:6928]},
     {storeUnit_maskInput_hi[6927:6912]},
     {storeUnit_maskInput_hi[6911:6896]},
     {storeUnit_maskInput_hi[6895:6880]},
     {storeUnit_maskInput_hi[6879:6864]},
     {storeUnit_maskInput_hi[6863:6848]},
     {storeUnit_maskInput_hi[6847:6832]},
     {storeUnit_maskInput_hi[6831:6816]},
     {storeUnit_maskInput_hi[6815:6800]},
     {storeUnit_maskInput_hi[6799:6784]},
     {storeUnit_maskInput_hi[6783:6768]},
     {storeUnit_maskInput_hi[6767:6752]},
     {storeUnit_maskInput_hi[6751:6736]},
     {storeUnit_maskInput_hi[6735:6720]},
     {storeUnit_maskInput_hi[6719:6704]},
     {storeUnit_maskInput_hi[6703:6688]},
     {storeUnit_maskInput_hi[6687:6672]},
     {storeUnit_maskInput_hi[6671:6656]},
     {storeUnit_maskInput_hi[6655:6640]},
     {storeUnit_maskInput_hi[6639:6624]},
     {storeUnit_maskInput_hi[6623:6608]},
     {storeUnit_maskInput_hi[6607:6592]},
     {storeUnit_maskInput_hi[6591:6576]},
     {storeUnit_maskInput_hi[6575:6560]},
     {storeUnit_maskInput_hi[6559:6544]},
     {storeUnit_maskInput_hi[6543:6528]},
     {storeUnit_maskInput_hi[6527:6512]},
     {storeUnit_maskInput_hi[6511:6496]},
     {storeUnit_maskInput_hi[6495:6480]},
     {storeUnit_maskInput_hi[6479:6464]},
     {storeUnit_maskInput_hi[6463:6448]},
     {storeUnit_maskInput_hi[6447:6432]},
     {storeUnit_maskInput_hi[6431:6416]},
     {storeUnit_maskInput_hi[6415:6400]},
     {storeUnit_maskInput_hi[6399:6384]},
     {storeUnit_maskInput_hi[6383:6368]},
     {storeUnit_maskInput_hi[6367:6352]},
     {storeUnit_maskInput_hi[6351:6336]},
     {storeUnit_maskInput_hi[6335:6320]},
     {storeUnit_maskInput_hi[6319:6304]},
     {storeUnit_maskInput_hi[6303:6288]},
     {storeUnit_maskInput_hi[6287:6272]},
     {storeUnit_maskInput_hi[6271:6256]},
     {storeUnit_maskInput_hi[6255:6240]},
     {storeUnit_maskInput_hi[6239:6224]},
     {storeUnit_maskInput_hi[6223:6208]},
     {storeUnit_maskInput_hi[6207:6192]},
     {storeUnit_maskInput_hi[6191:6176]},
     {storeUnit_maskInput_hi[6175:6160]},
     {storeUnit_maskInput_hi[6159:6144]},
     {storeUnit_maskInput_hi[6143:6128]},
     {storeUnit_maskInput_hi[6127:6112]},
     {storeUnit_maskInput_hi[6111:6096]},
     {storeUnit_maskInput_hi[6095:6080]},
     {storeUnit_maskInput_hi[6079:6064]},
     {storeUnit_maskInput_hi[6063:6048]},
     {storeUnit_maskInput_hi[6047:6032]},
     {storeUnit_maskInput_hi[6031:6016]},
     {storeUnit_maskInput_hi[6015:6000]},
     {storeUnit_maskInput_hi[5999:5984]},
     {storeUnit_maskInput_hi[5983:5968]},
     {storeUnit_maskInput_hi[5967:5952]},
     {storeUnit_maskInput_hi[5951:5936]},
     {storeUnit_maskInput_hi[5935:5920]},
     {storeUnit_maskInput_hi[5919:5904]},
     {storeUnit_maskInput_hi[5903:5888]},
     {storeUnit_maskInput_hi[5887:5872]},
     {storeUnit_maskInput_hi[5871:5856]},
     {storeUnit_maskInput_hi[5855:5840]},
     {storeUnit_maskInput_hi[5839:5824]},
     {storeUnit_maskInput_hi[5823:5808]},
     {storeUnit_maskInput_hi[5807:5792]},
     {storeUnit_maskInput_hi[5791:5776]},
     {storeUnit_maskInput_hi[5775:5760]},
     {storeUnit_maskInput_hi[5759:5744]},
     {storeUnit_maskInput_hi[5743:5728]},
     {storeUnit_maskInput_hi[5727:5712]},
     {storeUnit_maskInput_hi[5711:5696]},
     {storeUnit_maskInput_hi[5695:5680]},
     {storeUnit_maskInput_hi[5679:5664]},
     {storeUnit_maskInput_hi[5663:5648]},
     {storeUnit_maskInput_hi[5647:5632]},
     {storeUnit_maskInput_hi[5631:5616]},
     {storeUnit_maskInput_hi[5615:5600]},
     {storeUnit_maskInput_hi[5599:5584]},
     {storeUnit_maskInput_hi[5583:5568]},
     {storeUnit_maskInput_hi[5567:5552]},
     {storeUnit_maskInput_hi[5551:5536]},
     {storeUnit_maskInput_hi[5535:5520]},
     {storeUnit_maskInput_hi[5519:5504]},
     {storeUnit_maskInput_hi[5503:5488]},
     {storeUnit_maskInput_hi[5487:5472]},
     {storeUnit_maskInput_hi[5471:5456]},
     {storeUnit_maskInput_hi[5455:5440]},
     {storeUnit_maskInput_hi[5439:5424]},
     {storeUnit_maskInput_hi[5423:5408]},
     {storeUnit_maskInput_hi[5407:5392]},
     {storeUnit_maskInput_hi[5391:5376]},
     {storeUnit_maskInput_hi[5375:5360]},
     {storeUnit_maskInput_hi[5359:5344]},
     {storeUnit_maskInput_hi[5343:5328]},
     {storeUnit_maskInput_hi[5327:5312]},
     {storeUnit_maskInput_hi[5311:5296]},
     {storeUnit_maskInput_hi[5295:5280]},
     {storeUnit_maskInput_hi[5279:5264]},
     {storeUnit_maskInput_hi[5263:5248]},
     {storeUnit_maskInput_hi[5247:5232]},
     {storeUnit_maskInput_hi[5231:5216]},
     {storeUnit_maskInput_hi[5215:5200]},
     {storeUnit_maskInput_hi[5199:5184]},
     {storeUnit_maskInput_hi[5183:5168]},
     {storeUnit_maskInput_hi[5167:5152]},
     {storeUnit_maskInput_hi[5151:5136]},
     {storeUnit_maskInput_hi[5135:5120]},
     {storeUnit_maskInput_hi[5119:5104]},
     {storeUnit_maskInput_hi[5103:5088]},
     {storeUnit_maskInput_hi[5087:5072]},
     {storeUnit_maskInput_hi[5071:5056]},
     {storeUnit_maskInput_hi[5055:5040]},
     {storeUnit_maskInput_hi[5039:5024]},
     {storeUnit_maskInput_hi[5023:5008]},
     {storeUnit_maskInput_hi[5007:4992]},
     {storeUnit_maskInput_hi[4991:4976]},
     {storeUnit_maskInput_hi[4975:4960]},
     {storeUnit_maskInput_hi[4959:4944]},
     {storeUnit_maskInput_hi[4943:4928]},
     {storeUnit_maskInput_hi[4927:4912]},
     {storeUnit_maskInput_hi[4911:4896]},
     {storeUnit_maskInput_hi[4895:4880]},
     {storeUnit_maskInput_hi[4879:4864]},
     {storeUnit_maskInput_hi[4863:4848]},
     {storeUnit_maskInput_hi[4847:4832]},
     {storeUnit_maskInput_hi[4831:4816]},
     {storeUnit_maskInput_hi[4815:4800]},
     {storeUnit_maskInput_hi[4799:4784]},
     {storeUnit_maskInput_hi[4783:4768]},
     {storeUnit_maskInput_hi[4767:4752]},
     {storeUnit_maskInput_hi[4751:4736]},
     {storeUnit_maskInput_hi[4735:4720]},
     {storeUnit_maskInput_hi[4719:4704]},
     {storeUnit_maskInput_hi[4703:4688]},
     {storeUnit_maskInput_hi[4687:4672]},
     {storeUnit_maskInput_hi[4671:4656]},
     {storeUnit_maskInput_hi[4655:4640]},
     {storeUnit_maskInput_hi[4639:4624]},
     {storeUnit_maskInput_hi[4623:4608]},
     {storeUnit_maskInput_hi[4607:4592]},
     {storeUnit_maskInput_hi[4591:4576]},
     {storeUnit_maskInput_hi[4575:4560]},
     {storeUnit_maskInput_hi[4559:4544]},
     {storeUnit_maskInput_hi[4543:4528]},
     {storeUnit_maskInput_hi[4527:4512]},
     {storeUnit_maskInput_hi[4511:4496]},
     {storeUnit_maskInput_hi[4495:4480]},
     {storeUnit_maskInput_hi[4479:4464]},
     {storeUnit_maskInput_hi[4463:4448]},
     {storeUnit_maskInput_hi[4447:4432]},
     {storeUnit_maskInput_hi[4431:4416]},
     {storeUnit_maskInput_hi[4415:4400]},
     {storeUnit_maskInput_hi[4399:4384]},
     {storeUnit_maskInput_hi[4383:4368]},
     {storeUnit_maskInput_hi[4367:4352]},
     {storeUnit_maskInput_hi[4351:4336]},
     {storeUnit_maskInput_hi[4335:4320]},
     {storeUnit_maskInput_hi[4319:4304]},
     {storeUnit_maskInput_hi[4303:4288]},
     {storeUnit_maskInput_hi[4287:4272]},
     {storeUnit_maskInput_hi[4271:4256]},
     {storeUnit_maskInput_hi[4255:4240]},
     {storeUnit_maskInput_hi[4239:4224]},
     {storeUnit_maskInput_hi[4223:4208]},
     {storeUnit_maskInput_hi[4207:4192]},
     {storeUnit_maskInput_hi[4191:4176]},
     {storeUnit_maskInput_hi[4175:4160]},
     {storeUnit_maskInput_hi[4159:4144]},
     {storeUnit_maskInput_hi[4143:4128]},
     {storeUnit_maskInput_hi[4127:4112]},
     {storeUnit_maskInput_hi[4111:4096]},
     {storeUnit_maskInput_hi[4095:4080]},
     {storeUnit_maskInput_hi[4079:4064]},
     {storeUnit_maskInput_hi[4063:4048]},
     {storeUnit_maskInput_hi[4047:4032]},
     {storeUnit_maskInput_hi[4031:4016]},
     {storeUnit_maskInput_hi[4015:4000]},
     {storeUnit_maskInput_hi[3999:3984]},
     {storeUnit_maskInput_hi[3983:3968]},
     {storeUnit_maskInput_hi[3967:3952]},
     {storeUnit_maskInput_hi[3951:3936]},
     {storeUnit_maskInput_hi[3935:3920]},
     {storeUnit_maskInput_hi[3919:3904]},
     {storeUnit_maskInput_hi[3903:3888]},
     {storeUnit_maskInput_hi[3887:3872]},
     {storeUnit_maskInput_hi[3871:3856]},
     {storeUnit_maskInput_hi[3855:3840]},
     {storeUnit_maskInput_hi[3839:3824]},
     {storeUnit_maskInput_hi[3823:3808]},
     {storeUnit_maskInput_hi[3807:3792]},
     {storeUnit_maskInput_hi[3791:3776]},
     {storeUnit_maskInput_hi[3775:3760]},
     {storeUnit_maskInput_hi[3759:3744]},
     {storeUnit_maskInput_hi[3743:3728]},
     {storeUnit_maskInput_hi[3727:3712]},
     {storeUnit_maskInput_hi[3711:3696]},
     {storeUnit_maskInput_hi[3695:3680]},
     {storeUnit_maskInput_hi[3679:3664]},
     {storeUnit_maskInput_hi[3663:3648]},
     {storeUnit_maskInput_hi[3647:3632]},
     {storeUnit_maskInput_hi[3631:3616]},
     {storeUnit_maskInput_hi[3615:3600]},
     {storeUnit_maskInput_hi[3599:3584]},
     {storeUnit_maskInput_hi[3583:3568]},
     {storeUnit_maskInput_hi[3567:3552]},
     {storeUnit_maskInput_hi[3551:3536]},
     {storeUnit_maskInput_hi[3535:3520]},
     {storeUnit_maskInput_hi[3519:3504]},
     {storeUnit_maskInput_hi[3503:3488]},
     {storeUnit_maskInput_hi[3487:3472]},
     {storeUnit_maskInput_hi[3471:3456]},
     {storeUnit_maskInput_hi[3455:3440]},
     {storeUnit_maskInput_hi[3439:3424]},
     {storeUnit_maskInput_hi[3423:3408]},
     {storeUnit_maskInput_hi[3407:3392]},
     {storeUnit_maskInput_hi[3391:3376]},
     {storeUnit_maskInput_hi[3375:3360]},
     {storeUnit_maskInput_hi[3359:3344]},
     {storeUnit_maskInput_hi[3343:3328]},
     {storeUnit_maskInput_hi[3327:3312]},
     {storeUnit_maskInput_hi[3311:3296]},
     {storeUnit_maskInput_hi[3295:3280]},
     {storeUnit_maskInput_hi[3279:3264]},
     {storeUnit_maskInput_hi[3263:3248]},
     {storeUnit_maskInput_hi[3247:3232]},
     {storeUnit_maskInput_hi[3231:3216]},
     {storeUnit_maskInput_hi[3215:3200]},
     {storeUnit_maskInput_hi[3199:3184]},
     {storeUnit_maskInput_hi[3183:3168]},
     {storeUnit_maskInput_hi[3167:3152]},
     {storeUnit_maskInput_hi[3151:3136]},
     {storeUnit_maskInput_hi[3135:3120]},
     {storeUnit_maskInput_hi[3119:3104]},
     {storeUnit_maskInput_hi[3103:3088]},
     {storeUnit_maskInput_hi[3087:3072]},
     {storeUnit_maskInput_hi[3071:3056]},
     {storeUnit_maskInput_hi[3055:3040]},
     {storeUnit_maskInput_hi[3039:3024]},
     {storeUnit_maskInput_hi[3023:3008]},
     {storeUnit_maskInput_hi[3007:2992]},
     {storeUnit_maskInput_hi[2991:2976]},
     {storeUnit_maskInput_hi[2975:2960]},
     {storeUnit_maskInput_hi[2959:2944]},
     {storeUnit_maskInput_hi[2943:2928]},
     {storeUnit_maskInput_hi[2927:2912]},
     {storeUnit_maskInput_hi[2911:2896]},
     {storeUnit_maskInput_hi[2895:2880]},
     {storeUnit_maskInput_hi[2879:2864]},
     {storeUnit_maskInput_hi[2863:2848]},
     {storeUnit_maskInput_hi[2847:2832]},
     {storeUnit_maskInput_hi[2831:2816]},
     {storeUnit_maskInput_hi[2815:2800]},
     {storeUnit_maskInput_hi[2799:2784]},
     {storeUnit_maskInput_hi[2783:2768]},
     {storeUnit_maskInput_hi[2767:2752]},
     {storeUnit_maskInput_hi[2751:2736]},
     {storeUnit_maskInput_hi[2735:2720]},
     {storeUnit_maskInput_hi[2719:2704]},
     {storeUnit_maskInput_hi[2703:2688]},
     {storeUnit_maskInput_hi[2687:2672]},
     {storeUnit_maskInput_hi[2671:2656]},
     {storeUnit_maskInput_hi[2655:2640]},
     {storeUnit_maskInput_hi[2639:2624]},
     {storeUnit_maskInput_hi[2623:2608]},
     {storeUnit_maskInput_hi[2607:2592]},
     {storeUnit_maskInput_hi[2591:2576]},
     {storeUnit_maskInput_hi[2575:2560]},
     {storeUnit_maskInput_hi[2559:2544]},
     {storeUnit_maskInput_hi[2543:2528]},
     {storeUnit_maskInput_hi[2527:2512]},
     {storeUnit_maskInput_hi[2511:2496]},
     {storeUnit_maskInput_hi[2495:2480]},
     {storeUnit_maskInput_hi[2479:2464]},
     {storeUnit_maskInput_hi[2463:2448]},
     {storeUnit_maskInput_hi[2447:2432]},
     {storeUnit_maskInput_hi[2431:2416]},
     {storeUnit_maskInput_hi[2415:2400]},
     {storeUnit_maskInput_hi[2399:2384]},
     {storeUnit_maskInput_hi[2383:2368]},
     {storeUnit_maskInput_hi[2367:2352]},
     {storeUnit_maskInput_hi[2351:2336]},
     {storeUnit_maskInput_hi[2335:2320]},
     {storeUnit_maskInput_hi[2319:2304]},
     {storeUnit_maskInput_hi[2303:2288]},
     {storeUnit_maskInput_hi[2287:2272]},
     {storeUnit_maskInput_hi[2271:2256]},
     {storeUnit_maskInput_hi[2255:2240]},
     {storeUnit_maskInput_hi[2239:2224]},
     {storeUnit_maskInput_hi[2223:2208]},
     {storeUnit_maskInput_hi[2207:2192]},
     {storeUnit_maskInput_hi[2191:2176]},
     {storeUnit_maskInput_hi[2175:2160]},
     {storeUnit_maskInput_hi[2159:2144]},
     {storeUnit_maskInput_hi[2143:2128]},
     {storeUnit_maskInput_hi[2127:2112]},
     {storeUnit_maskInput_hi[2111:2096]},
     {storeUnit_maskInput_hi[2095:2080]},
     {storeUnit_maskInput_hi[2079:2064]},
     {storeUnit_maskInput_hi[2063:2048]},
     {storeUnit_maskInput_hi[2047:2032]},
     {storeUnit_maskInput_hi[2031:2016]},
     {storeUnit_maskInput_hi[2015:2000]},
     {storeUnit_maskInput_hi[1999:1984]},
     {storeUnit_maskInput_hi[1983:1968]},
     {storeUnit_maskInput_hi[1967:1952]},
     {storeUnit_maskInput_hi[1951:1936]},
     {storeUnit_maskInput_hi[1935:1920]},
     {storeUnit_maskInput_hi[1919:1904]},
     {storeUnit_maskInput_hi[1903:1888]},
     {storeUnit_maskInput_hi[1887:1872]},
     {storeUnit_maskInput_hi[1871:1856]},
     {storeUnit_maskInput_hi[1855:1840]},
     {storeUnit_maskInput_hi[1839:1824]},
     {storeUnit_maskInput_hi[1823:1808]},
     {storeUnit_maskInput_hi[1807:1792]},
     {storeUnit_maskInput_hi[1791:1776]},
     {storeUnit_maskInput_hi[1775:1760]},
     {storeUnit_maskInput_hi[1759:1744]},
     {storeUnit_maskInput_hi[1743:1728]},
     {storeUnit_maskInput_hi[1727:1712]},
     {storeUnit_maskInput_hi[1711:1696]},
     {storeUnit_maskInput_hi[1695:1680]},
     {storeUnit_maskInput_hi[1679:1664]},
     {storeUnit_maskInput_hi[1663:1648]},
     {storeUnit_maskInput_hi[1647:1632]},
     {storeUnit_maskInput_hi[1631:1616]},
     {storeUnit_maskInput_hi[1615:1600]},
     {storeUnit_maskInput_hi[1599:1584]},
     {storeUnit_maskInput_hi[1583:1568]},
     {storeUnit_maskInput_hi[1567:1552]},
     {storeUnit_maskInput_hi[1551:1536]},
     {storeUnit_maskInput_hi[1535:1520]},
     {storeUnit_maskInput_hi[1519:1504]},
     {storeUnit_maskInput_hi[1503:1488]},
     {storeUnit_maskInput_hi[1487:1472]},
     {storeUnit_maskInput_hi[1471:1456]},
     {storeUnit_maskInput_hi[1455:1440]},
     {storeUnit_maskInput_hi[1439:1424]},
     {storeUnit_maskInput_hi[1423:1408]},
     {storeUnit_maskInput_hi[1407:1392]},
     {storeUnit_maskInput_hi[1391:1376]},
     {storeUnit_maskInput_hi[1375:1360]},
     {storeUnit_maskInput_hi[1359:1344]},
     {storeUnit_maskInput_hi[1343:1328]},
     {storeUnit_maskInput_hi[1327:1312]},
     {storeUnit_maskInput_hi[1311:1296]},
     {storeUnit_maskInput_hi[1295:1280]},
     {storeUnit_maskInput_hi[1279:1264]},
     {storeUnit_maskInput_hi[1263:1248]},
     {storeUnit_maskInput_hi[1247:1232]},
     {storeUnit_maskInput_hi[1231:1216]},
     {storeUnit_maskInput_hi[1215:1200]},
     {storeUnit_maskInput_hi[1199:1184]},
     {storeUnit_maskInput_hi[1183:1168]},
     {storeUnit_maskInput_hi[1167:1152]},
     {storeUnit_maskInput_hi[1151:1136]},
     {storeUnit_maskInput_hi[1135:1120]},
     {storeUnit_maskInput_hi[1119:1104]},
     {storeUnit_maskInput_hi[1103:1088]},
     {storeUnit_maskInput_hi[1087:1072]},
     {storeUnit_maskInput_hi[1071:1056]},
     {storeUnit_maskInput_hi[1055:1040]},
     {storeUnit_maskInput_hi[1039:1024]},
     {storeUnit_maskInput_hi[1023:1008]},
     {storeUnit_maskInput_hi[1007:992]},
     {storeUnit_maskInput_hi[991:976]},
     {storeUnit_maskInput_hi[975:960]},
     {storeUnit_maskInput_hi[959:944]},
     {storeUnit_maskInput_hi[943:928]},
     {storeUnit_maskInput_hi[927:912]},
     {storeUnit_maskInput_hi[911:896]},
     {storeUnit_maskInput_hi[895:880]},
     {storeUnit_maskInput_hi[879:864]},
     {storeUnit_maskInput_hi[863:848]},
     {storeUnit_maskInput_hi[847:832]},
     {storeUnit_maskInput_hi[831:816]},
     {storeUnit_maskInput_hi[815:800]},
     {storeUnit_maskInput_hi[799:784]},
     {storeUnit_maskInput_hi[783:768]},
     {storeUnit_maskInput_hi[767:752]},
     {storeUnit_maskInput_hi[751:736]},
     {storeUnit_maskInput_hi[735:720]},
     {storeUnit_maskInput_hi[719:704]},
     {storeUnit_maskInput_hi[703:688]},
     {storeUnit_maskInput_hi[687:672]},
     {storeUnit_maskInput_hi[671:656]},
     {storeUnit_maskInput_hi[655:640]},
     {storeUnit_maskInput_hi[639:624]},
     {storeUnit_maskInput_hi[623:608]},
     {storeUnit_maskInput_hi[607:592]},
     {storeUnit_maskInput_hi[591:576]},
     {storeUnit_maskInput_hi[575:560]},
     {storeUnit_maskInput_hi[559:544]},
     {storeUnit_maskInput_hi[543:528]},
     {storeUnit_maskInput_hi[527:512]},
     {storeUnit_maskInput_hi[511:496]},
     {storeUnit_maskInput_hi[495:480]},
     {storeUnit_maskInput_hi[479:464]},
     {storeUnit_maskInput_hi[463:448]},
     {storeUnit_maskInput_hi[447:432]},
     {storeUnit_maskInput_hi[431:416]},
     {storeUnit_maskInput_hi[415:400]},
     {storeUnit_maskInput_hi[399:384]},
     {storeUnit_maskInput_hi[383:368]},
     {storeUnit_maskInput_hi[367:352]},
     {storeUnit_maskInput_hi[351:336]},
     {storeUnit_maskInput_hi[335:320]},
     {storeUnit_maskInput_hi[319:304]},
     {storeUnit_maskInput_hi[303:288]},
     {storeUnit_maskInput_hi[287:272]},
     {storeUnit_maskInput_hi[271:256]},
     {storeUnit_maskInput_hi[255:240]},
     {storeUnit_maskInput_hi[239:224]},
     {storeUnit_maskInput_hi[223:208]},
     {storeUnit_maskInput_hi[207:192]},
     {storeUnit_maskInput_hi[191:176]},
     {storeUnit_maskInput_hi[175:160]},
     {storeUnit_maskInput_hi[159:144]},
     {storeUnit_maskInput_hi[143:128]},
     {storeUnit_maskInput_hi[127:112]},
     {storeUnit_maskInput_hi[111:96]},
     {storeUnit_maskInput_hi[95:80]},
     {storeUnit_maskInput_hi[79:64]},
     {storeUnit_maskInput_hi[63:48]},
     {storeUnit_maskInput_hi[47:32]},
     {storeUnit_maskInput_hi[31:16]},
     {storeUnit_maskInput_hi[15:0]},
     {storeUnit_maskInput_lo[32767:32752]},
     {storeUnit_maskInput_lo[32751:32736]},
     {storeUnit_maskInput_lo[32735:32720]},
     {storeUnit_maskInput_lo[32719:32704]},
     {storeUnit_maskInput_lo[32703:32688]},
     {storeUnit_maskInput_lo[32687:32672]},
     {storeUnit_maskInput_lo[32671:32656]},
     {storeUnit_maskInput_lo[32655:32640]},
     {storeUnit_maskInput_lo[32639:32624]},
     {storeUnit_maskInput_lo[32623:32608]},
     {storeUnit_maskInput_lo[32607:32592]},
     {storeUnit_maskInput_lo[32591:32576]},
     {storeUnit_maskInput_lo[32575:32560]},
     {storeUnit_maskInput_lo[32559:32544]},
     {storeUnit_maskInput_lo[32543:32528]},
     {storeUnit_maskInput_lo[32527:32512]},
     {storeUnit_maskInput_lo[32511:32496]},
     {storeUnit_maskInput_lo[32495:32480]},
     {storeUnit_maskInput_lo[32479:32464]},
     {storeUnit_maskInput_lo[32463:32448]},
     {storeUnit_maskInput_lo[32447:32432]},
     {storeUnit_maskInput_lo[32431:32416]},
     {storeUnit_maskInput_lo[32415:32400]},
     {storeUnit_maskInput_lo[32399:32384]},
     {storeUnit_maskInput_lo[32383:32368]},
     {storeUnit_maskInput_lo[32367:32352]},
     {storeUnit_maskInput_lo[32351:32336]},
     {storeUnit_maskInput_lo[32335:32320]},
     {storeUnit_maskInput_lo[32319:32304]},
     {storeUnit_maskInput_lo[32303:32288]},
     {storeUnit_maskInput_lo[32287:32272]},
     {storeUnit_maskInput_lo[32271:32256]},
     {storeUnit_maskInput_lo[32255:32240]},
     {storeUnit_maskInput_lo[32239:32224]},
     {storeUnit_maskInput_lo[32223:32208]},
     {storeUnit_maskInput_lo[32207:32192]},
     {storeUnit_maskInput_lo[32191:32176]},
     {storeUnit_maskInput_lo[32175:32160]},
     {storeUnit_maskInput_lo[32159:32144]},
     {storeUnit_maskInput_lo[32143:32128]},
     {storeUnit_maskInput_lo[32127:32112]},
     {storeUnit_maskInput_lo[32111:32096]},
     {storeUnit_maskInput_lo[32095:32080]},
     {storeUnit_maskInput_lo[32079:32064]},
     {storeUnit_maskInput_lo[32063:32048]},
     {storeUnit_maskInput_lo[32047:32032]},
     {storeUnit_maskInput_lo[32031:32016]},
     {storeUnit_maskInput_lo[32015:32000]},
     {storeUnit_maskInput_lo[31999:31984]},
     {storeUnit_maskInput_lo[31983:31968]},
     {storeUnit_maskInput_lo[31967:31952]},
     {storeUnit_maskInput_lo[31951:31936]},
     {storeUnit_maskInput_lo[31935:31920]},
     {storeUnit_maskInput_lo[31919:31904]},
     {storeUnit_maskInput_lo[31903:31888]},
     {storeUnit_maskInput_lo[31887:31872]},
     {storeUnit_maskInput_lo[31871:31856]},
     {storeUnit_maskInput_lo[31855:31840]},
     {storeUnit_maskInput_lo[31839:31824]},
     {storeUnit_maskInput_lo[31823:31808]},
     {storeUnit_maskInput_lo[31807:31792]},
     {storeUnit_maskInput_lo[31791:31776]},
     {storeUnit_maskInput_lo[31775:31760]},
     {storeUnit_maskInput_lo[31759:31744]},
     {storeUnit_maskInput_lo[31743:31728]},
     {storeUnit_maskInput_lo[31727:31712]},
     {storeUnit_maskInput_lo[31711:31696]},
     {storeUnit_maskInput_lo[31695:31680]},
     {storeUnit_maskInput_lo[31679:31664]},
     {storeUnit_maskInput_lo[31663:31648]},
     {storeUnit_maskInput_lo[31647:31632]},
     {storeUnit_maskInput_lo[31631:31616]},
     {storeUnit_maskInput_lo[31615:31600]},
     {storeUnit_maskInput_lo[31599:31584]},
     {storeUnit_maskInput_lo[31583:31568]},
     {storeUnit_maskInput_lo[31567:31552]},
     {storeUnit_maskInput_lo[31551:31536]},
     {storeUnit_maskInput_lo[31535:31520]},
     {storeUnit_maskInput_lo[31519:31504]},
     {storeUnit_maskInput_lo[31503:31488]},
     {storeUnit_maskInput_lo[31487:31472]},
     {storeUnit_maskInput_lo[31471:31456]},
     {storeUnit_maskInput_lo[31455:31440]},
     {storeUnit_maskInput_lo[31439:31424]},
     {storeUnit_maskInput_lo[31423:31408]},
     {storeUnit_maskInput_lo[31407:31392]},
     {storeUnit_maskInput_lo[31391:31376]},
     {storeUnit_maskInput_lo[31375:31360]},
     {storeUnit_maskInput_lo[31359:31344]},
     {storeUnit_maskInput_lo[31343:31328]},
     {storeUnit_maskInput_lo[31327:31312]},
     {storeUnit_maskInput_lo[31311:31296]},
     {storeUnit_maskInput_lo[31295:31280]},
     {storeUnit_maskInput_lo[31279:31264]},
     {storeUnit_maskInput_lo[31263:31248]},
     {storeUnit_maskInput_lo[31247:31232]},
     {storeUnit_maskInput_lo[31231:31216]},
     {storeUnit_maskInput_lo[31215:31200]},
     {storeUnit_maskInput_lo[31199:31184]},
     {storeUnit_maskInput_lo[31183:31168]},
     {storeUnit_maskInput_lo[31167:31152]},
     {storeUnit_maskInput_lo[31151:31136]},
     {storeUnit_maskInput_lo[31135:31120]},
     {storeUnit_maskInput_lo[31119:31104]},
     {storeUnit_maskInput_lo[31103:31088]},
     {storeUnit_maskInput_lo[31087:31072]},
     {storeUnit_maskInput_lo[31071:31056]},
     {storeUnit_maskInput_lo[31055:31040]},
     {storeUnit_maskInput_lo[31039:31024]},
     {storeUnit_maskInput_lo[31023:31008]},
     {storeUnit_maskInput_lo[31007:30992]},
     {storeUnit_maskInput_lo[30991:30976]},
     {storeUnit_maskInput_lo[30975:30960]},
     {storeUnit_maskInput_lo[30959:30944]},
     {storeUnit_maskInput_lo[30943:30928]},
     {storeUnit_maskInput_lo[30927:30912]},
     {storeUnit_maskInput_lo[30911:30896]},
     {storeUnit_maskInput_lo[30895:30880]},
     {storeUnit_maskInput_lo[30879:30864]},
     {storeUnit_maskInput_lo[30863:30848]},
     {storeUnit_maskInput_lo[30847:30832]},
     {storeUnit_maskInput_lo[30831:30816]},
     {storeUnit_maskInput_lo[30815:30800]},
     {storeUnit_maskInput_lo[30799:30784]},
     {storeUnit_maskInput_lo[30783:30768]},
     {storeUnit_maskInput_lo[30767:30752]},
     {storeUnit_maskInput_lo[30751:30736]},
     {storeUnit_maskInput_lo[30735:30720]},
     {storeUnit_maskInput_lo[30719:30704]},
     {storeUnit_maskInput_lo[30703:30688]},
     {storeUnit_maskInput_lo[30687:30672]},
     {storeUnit_maskInput_lo[30671:30656]},
     {storeUnit_maskInput_lo[30655:30640]},
     {storeUnit_maskInput_lo[30639:30624]},
     {storeUnit_maskInput_lo[30623:30608]},
     {storeUnit_maskInput_lo[30607:30592]},
     {storeUnit_maskInput_lo[30591:30576]},
     {storeUnit_maskInput_lo[30575:30560]},
     {storeUnit_maskInput_lo[30559:30544]},
     {storeUnit_maskInput_lo[30543:30528]},
     {storeUnit_maskInput_lo[30527:30512]},
     {storeUnit_maskInput_lo[30511:30496]},
     {storeUnit_maskInput_lo[30495:30480]},
     {storeUnit_maskInput_lo[30479:30464]},
     {storeUnit_maskInput_lo[30463:30448]},
     {storeUnit_maskInput_lo[30447:30432]},
     {storeUnit_maskInput_lo[30431:30416]},
     {storeUnit_maskInput_lo[30415:30400]},
     {storeUnit_maskInput_lo[30399:30384]},
     {storeUnit_maskInput_lo[30383:30368]},
     {storeUnit_maskInput_lo[30367:30352]},
     {storeUnit_maskInput_lo[30351:30336]},
     {storeUnit_maskInput_lo[30335:30320]},
     {storeUnit_maskInput_lo[30319:30304]},
     {storeUnit_maskInput_lo[30303:30288]},
     {storeUnit_maskInput_lo[30287:30272]},
     {storeUnit_maskInput_lo[30271:30256]},
     {storeUnit_maskInput_lo[30255:30240]},
     {storeUnit_maskInput_lo[30239:30224]},
     {storeUnit_maskInput_lo[30223:30208]},
     {storeUnit_maskInput_lo[30207:30192]},
     {storeUnit_maskInput_lo[30191:30176]},
     {storeUnit_maskInput_lo[30175:30160]},
     {storeUnit_maskInput_lo[30159:30144]},
     {storeUnit_maskInput_lo[30143:30128]},
     {storeUnit_maskInput_lo[30127:30112]},
     {storeUnit_maskInput_lo[30111:30096]},
     {storeUnit_maskInput_lo[30095:30080]},
     {storeUnit_maskInput_lo[30079:30064]},
     {storeUnit_maskInput_lo[30063:30048]},
     {storeUnit_maskInput_lo[30047:30032]},
     {storeUnit_maskInput_lo[30031:30016]},
     {storeUnit_maskInput_lo[30015:30000]},
     {storeUnit_maskInput_lo[29999:29984]},
     {storeUnit_maskInput_lo[29983:29968]},
     {storeUnit_maskInput_lo[29967:29952]},
     {storeUnit_maskInput_lo[29951:29936]},
     {storeUnit_maskInput_lo[29935:29920]},
     {storeUnit_maskInput_lo[29919:29904]},
     {storeUnit_maskInput_lo[29903:29888]},
     {storeUnit_maskInput_lo[29887:29872]},
     {storeUnit_maskInput_lo[29871:29856]},
     {storeUnit_maskInput_lo[29855:29840]},
     {storeUnit_maskInput_lo[29839:29824]},
     {storeUnit_maskInput_lo[29823:29808]},
     {storeUnit_maskInput_lo[29807:29792]},
     {storeUnit_maskInput_lo[29791:29776]},
     {storeUnit_maskInput_lo[29775:29760]},
     {storeUnit_maskInput_lo[29759:29744]},
     {storeUnit_maskInput_lo[29743:29728]},
     {storeUnit_maskInput_lo[29727:29712]},
     {storeUnit_maskInput_lo[29711:29696]},
     {storeUnit_maskInput_lo[29695:29680]},
     {storeUnit_maskInput_lo[29679:29664]},
     {storeUnit_maskInput_lo[29663:29648]},
     {storeUnit_maskInput_lo[29647:29632]},
     {storeUnit_maskInput_lo[29631:29616]},
     {storeUnit_maskInput_lo[29615:29600]},
     {storeUnit_maskInput_lo[29599:29584]},
     {storeUnit_maskInput_lo[29583:29568]},
     {storeUnit_maskInput_lo[29567:29552]},
     {storeUnit_maskInput_lo[29551:29536]},
     {storeUnit_maskInput_lo[29535:29520]},
     {storeUnit_maskInput_lo[29519:29504]},
     {storeUnit_maskInput_lo[29503:29488]},
     {storeUnit_maskInput_lo[29487:29472]},
     {storeUnit_maskInput_lo[29471:29456]},
     {storeUnit_maskInput_lo[29455:29440]},
     {storeUnit_maskInput_lo[29439:29424]},
     {storeUnit_maskInput_lo[29423:29408]},
     {storeUnit_maskInput_lo[29407:29392]},
     {storeUnit_maskInput_lo[29391:29376]},
     {storeUnit_maskInput_lo[29375:29360]},
     {storeUnit_maskInput_lo[29359:29344]},
     {storeUnit_maskInput_lo[29343:29328]},
     {storeUnit_maskInput_lo[29327:29312]},
     {storeUnit_maskInput_lo[29311:29296]},
     {storeUnit_maskInput_lo[29295:29280]},
     {storeUnit_maskInput_lo[29279:29264]},
     {storeUnit_maskInput_lo[29263:29248]},
     {storeUnit_maskInput_lo[29247:29232]},
     {storeUnit_maskInput_lo[29231:29216]},
     {storeUnit_maskInput_lo[29215:29200]},
     {storeUnit_maskInput_lo[29199:29184]},
     {storeUnit_maskInput_lo[29183:29168]},
     {storeUnit_maskInput_lo[29167:29152]},
     {storeUnit_maskInput_lo[29151:29136]},
     {storeUnit_maskInput_lo[29135:29120]},
     {storeUnit_maskInput_lo[29119:29104]},
     {storeUnit_maskInput_lo[29103:29088]},
     {storeUnit_maskInput_lo[29087:29072]},
     {storeUnit_maskInput_lo[29071:29056]},
     {storeUnit_maskInput_lo[29055:29040]},
     {storeUnit_maskInput_lo[29039:29024]},
     {storeUnit_maskInput_lo[29023:29008]},
     {storeUnit_maskInput_lo[29007:28992]},
     {storeUnit_maskInput_lo[28991:28976]},
     {storeUnit_maskInput_lo[28975:28960]},
     {storeUnit_maskInput_lo[28959:28944]},
     {storeUnit_maskInput_lo[28943:28928]},
     {storeUnit_maskInput_lo[28927:28912]},
     {storeUnit_maskInput_lo[28911:28896]},
     {storeUnit_maskInput_lo[28895:28880]},
     {storeUnit_maskInput_lo[28879:28864]},
     {storeUnit_maskInput_lo[28863:28848]},
     {storeUnit_maskInput_lo[28847:28832]},
     {storeUnit_maskInput_lo[28831:28816]},
     {storeUnit_maskInput_lo[28815:28800]},
     {storeUnit_maskInput_lo[28799:28784]},
     {storeUnit_maskInput_lo[28783:28768]},
     {storeUnit_maskInput_lo[28767:28752]},
     {storeUnit_maskInput_lo[28751:28736]},
     {storeUnit_maskInput_lo[28735:28720]},
     {storeUnit_maskInput_lo[28719:28704]},
     {storeUnit_maskInput_lo[28703:28688]},
     {storeUnit_maskInput_lo[28687:28672]},
     {storeUnit_maskInput_lo[28671:28656]},
     {storeUnit_maskInput_lo[28655:28640]},
     {storeUnit_maskInput_lo[28639:28624]},
     {storeUnit_maskInput_lo[28623:28608]},
     {storeUnit_maskInput_lo[28607:28592]},
     {storeUnit_maskInput_lo[28591:28576]},
     {storeUnit_maskInput_lo[28575:28560]},
     {storeUnit_maskInput_lo[28559:28544]},
     {storeUnit_maskInput_lo[28543:28528]},
     {storeUnit_maskInput_lo[28527:28512]},
     {storeUnit_maskInput_lo[28511:28496]},
     {storeUnit_maskInput_lo[28495:28480]},
     {storeUnit_maskInput_lo[28479:28464]},
     {storeUnit_maskInput_lo[28463:28448]},
     {storeUnit_maskInput_lo[28447:28432]},
     {storeUnit_maskInput_lo[28431:28416]},
     {storeUnit_maskInput_lo[28415:28400]},
     {storeUnit_maskInput_lo[28399:28384]},
     {storeUnit_maskInput_lo[28383:28368]},
     {storeUnit_maskInput_lo[28367:28352]},
     {storeUnit_maskInput_lo[28351:28336]},
     {storeUnit_maskInput_lo[28335:28320]},
     {storeUnit_maskInput_lo[28319:28304]},
     {storeUnit_maskInput_lo[28303:28288]},
     {storeUnit_maskInput_lo[28287:28272]},
     {storeUnit_maskInput_lo[28271:28256]},
     {storeUnit_maskInput_lo[28255:28240]},
     {storeUnit_maskInput_lo[28239:28224]},
     {storeUnit_maskInput_lo[28223:28208]},
     {storeUnit_maskInput_lo[28207:28192]},
     {storeUnit_maskInput_lo[28191:28176]},
     {storeUnit_maskInput_lo[28175:28160]},
     {storeUnit_maskInput_lo[28159:28144]},
     {storeUnit_maskInput_lo[28143:28128]},
     {storeUnit_maskInput_lo[28127:28112]},
     {storeUnit_maskInput_lo[28111:28096]},
     {storeUnit_maskInput_lo[28095:28080]},
     {storeUnit_maskInput_lo[28079:28064]},
     {storeUnit_maskInput_lo[28063:28048]},
     {storeUnit_maskInput_lo[28047:28032]},
     {storeUnit_maskInput_lo[28031:28016]},
     {storeUnit_maskInput_lo[28015:28000]},
     {storeUnit_maskInput_lo[27999:27984]},
     {storeUnit_maskInput_lo[27983:27968]},
     {storeUnit_maskInput_lo[27967:27952]},
     {storeUnit_maskInput_lo[27951:27936]},
     {storeUnit_maskInput_lo[27935:27920]},
     {storeUnit_maskInput_lo[27919:27904]},
     {storeUnit_maskInput_lo[27903:27888]},
     {storeUnit_maskInput_lo[27887:27872]},
     {storeUnit_maskInput_lo[27871:27856]},
     {storeUnit_maskInput_lo[27855:27840]},
     {storeUnit_maskInput_lo[27839:27824]},
     {storeUnit_maskInput_lo[27823:27808]},
     {storeUnit_maskInput_lo[27807:27792]},
     {storeUnit_maskInput_lo[27791:27776]},
     {storeUnit_maskInput_lo[27775:27760]},
     {storeUnit_maskInput_lo[27759:27744]},
     {storeUnit_maskInput_lo[27743:27728]},
     {storeUnit_maskInput_lo[27727:27712]},
     {storeUnit_maskInput_lo[27711:27696]},
     {storeUnit_maskInput_lo[27695:27680]},
     {storeUnit_maskInput_lo[27679:27664]},
     {storeUnit_maskInput_lo[27663:27648]},
     {storeUnit_maskInput_lo[27647:27632]},
     {storeUnit_maskInput_lo[27631:27616]},
     {storeUnit_maskInput_lo[27615:27600]},
     {storeUnit_maskInput_lo[27599:27584]},
     {storeUnit_maskInput_lo[27583:27568]},
     {storeUnit_maskInput_lo[27567:27552]},
     {storeUnit_maskInput_lo[27551:27536]},
     {storeUnit_maskInput_lo[27535:27520]},
     {storeUnit_maskInput_lo[27519:27504]},
     {storeUnit_maskInput_lo[27503:27488]},
     {storeUnit_maskInput_lo[27487:27472]},
     {storeUnit_maskInput_lo[27471:27456]},
     {storeUnit_maskInput_lo[27455:27440]},
     {storeUnit_maskInput_lo[27439:27424]},
     {storeUnit_maskInput_lo[27423:27408]},
     {storeUnit_maskInput_lo[27407:27392]},
     {storeUnit_maskInput_lo[27391:27376]},
     {storeUnit_maskInput_lo[27375:27360]},
     {storeUnit_maskInput_lo[27359:27344]},
     {storeUnit_maskInput_lo[27343:27328]},
     {storeUnit_maskInput_lo[27327:27312]},
     {storeUnit_maskInput_lo[27311:27296]},
     {storeUnit_maskInput_lo[27295:27280]},
     {storeUnit_maskInput_lo[27279:27264]},
     {storeUnit_maskInput_lo[27263:27248]},
     {storeUnit_maskInput_lo[27247:27232]},
     {storeUnit_maskInput_lo[27231:27216]},
     {storeUnit_maskInput_lo[27215:27200]},
     {storeUnit_maskInput_lo[27199:27184]},
     {storeUnit_maskInput_lo[27183:27168]},
     {storeUnit_maskInput_lo[27167:27152]},
     {storeUnit_maskInput_lo[27151:27136]},
     {storeUnit_maskInput_lo[27135:27120]},
     {storeUnit_maskInput_lo[27119:27104]},
     {storeUnit_maskInput_lo[27103:27088]},
     {storeUnit_maskInput_lo[27087:27072]},
     {storeUnit_maskInput_lo[27071:27056]},
     {storeUnit_maskInput_lo[27055:27040]},
     {storeUnit_maskInput_lo[27039:27024]},
     {storeUnit_maskInput_lo[27023:27008]},
     {storeUnit_maskInput_lo[27007:26992]},
     {storeUnit_maskInput_lo[26991:26976]},
     {storeUnit_maskInput_lo[26975:26960]},
     {storeUnit_maskInput_lo[26959:26944]},
     {storeUnit_maskInput_lo[26943:26928]},
     {storeUnit_maskInput_lo[26927:26912]},
     {storeUnit_maskInput_lo[26911:26896]},
     {storeUnit_maskInput_lo[26895:26880]},
     {storeUnit_maskInput_lo[26879:26864]},
     {storeUnit_maskInput_lo[26863:26848]},
     {storeUnit_maskInput_lo[26847:26832]},
     {storeUnit_maskInput_lo[26831:26816]},
     {storeUnit_maskInput_lo[26815:26800]},
     {storeUnit_maskInput_lo[26799:26784]},
     {storeUnit_maskInput_lo[26783:26768]},
     {storeUnit_maskInput_lo[26767:26752]},
     {storeUnit_maskInput_lo[26751:26736]},
     {storeUnit_maskInput_lo[26735:26720]},
     {storeUnit_maskInput_lo[26719:26704]},
     {storeUnit_maskInput_lo[26703:26688]},
     {storeUnit_maskInput_lo[26687:26672]},
     {storeUnit_maskInput_lo[26671:26656]},
     {storeUnit_maskInput_lo[26655:26640]},
     {storeUnit_maskInput_lo[26639:26624]},
     {storeUnit_maskInput_lo[26623:26608]},
     {storeUnit_maskInput_lo[26607:26592]},
     {storeUnit_maskInput_lo[26591:26576]},
     {storeUnit_maskInput_lo[26575:26560]},
     {storeUnit_maskInput_lo[26559:26544]},
     {storeUnit_maskInput_lo[26543:26528]},
     {storeUnit_maskInput_lo[26527:26512]},
     {storeUnit_maskInput_lo[26511:26496]},
     {storeUnit_maskInput_lo[26495:26480]},
     {storeUnit_maskInput_lo[26479:26464]},
     {storeUnit_maskInput_lo[26463:26448]},
     {storeUnit_maskInput_lo[26447:26432]},
     {storeUnit_maskInput_lo[26431:26416]},
     {storeUnit_maskInput_lo[26415:26400]},
     {storeUnit_maskInput_lo[26399:26384]},
     {storeUnit_maskInput_lo[26383:26368]},
     {storeUnit_maskInput_lo[26367:26352]},
     {storeUnit_maskInput_lo[26351:26336]},
     {storeUnit_maskInput_lo[26335:26320]},
     {storeUnit_maskInput_lo[26319:26304]},
     {storeUnit_maskInput_lo[26303:26288]},
     {storeUnit_maskInput_lo[26287:26272]},
     {storeUnit_maskInput_lo[26271:26256]},
     {storeUnit_maskInput_lo[26255:26240]},
     {storeUnit_maskInput_lo[26239:26224]},
     {storeUnit_maskInput_lo[26223:26208]},
     {storeUnit_maskInput_lo[26207:26192]},
     {storeUnit_maskInput_lo[26191:26176]},
     {storeUnit_maskInput_lo[26175:26160]},
     {storeUnit_maskInput_lo[26159:26144]},
     {storeUnit_maskInput_lo[26143:26128]},
     {storeUnit_maskInput_lo[26127:26112]},
     {storeUnit_maskInput_lo[26111:26096]},
     {storeUnit_maskInput_lo[26095:26080]},
     {storeUnit_maskInput_lo[26079:26064]},
     {storeUnit_maskInput_lo[26063:26048]},
     {storeUnit_maskInput_lo[26047:26032]},
     {storeUnit_maskInput_lo[26031:26016]},
     {storeUnit_maskInput_lo[26015:26000]},
     {storeUnit_maskInput_lo[25999:25984]},
     {storeUnit_maskInput_lo[25983:25968]},
     {storeUnit_maskInput_lo[25967:25952]},
     {storeUnit_maskInput_lo[25951:25936]},
     {storeUnit_maskInput_lo[25935:25920]},
     {storeUnit_maskInput_lo[25919:25904]},
     {storeUnit_maskInput_lo[25903:25888]},
     {storeUnit_maskInput_lo[25887:25872]},
     {storeUnit_maskInput_lo[25871:25856]},
     {storeUnit_maskInput_lo[25855:25840]},
     {storeUnit_maskInput_lo[25839:25824]},
     {storeUnit_maskInput_lo[25823:25808]},
     {storeUnit_maskInput_lo[25807:25792]},
     {storeUnit_maskInput_lo[25791:25776]},
     {storeUnit_maskInput_lo[25775:25760]},
     {storeUnit_maskInput_lo[25759:25744]},
     {storeUnit_maskInput_lo[25743:25728]},
     {storeUnit_maskInput_lo[25727:25712]},
     {storeUnit_maskInput_lo[25711:25696]},
     {storeUnit_maskInput_lo[25695:25680]},
     {storeUnit_maskInput_lo[25679:25664]},
     {storeUnit_maskInput_lo[25663:25648]},
     {storeUnit_maskInput_lo[25647:25632]},
     {storeUnit_maskInput_lo[25631:25616]},
     {storeUnit_maskInput_lo[25615:25600]},
     {storeUnit_maskInput_lo[25599:25584]},
     {storeUnit_maskInput_lo[25583:25568]},
     {storeUnit_maskInput_lo[25567:25552]},
     {storeUnit_maskInput_lo[25551:25536]},
     {storeUnit_maskInput_lo[25535:25520]},
     {storeUnit_maskInput_lo[25519:25504]},
     {storeUnit_maskInput_lo[25503:25488]},
     {storeUnit_maskInput_lo[25487:25472]},
     {storeUnit_maskInput_lo[25471:25456]},
     {storeUnit_maskInput_lo[25455:25440]},
     {storeUnit_maskInput_lo[25439:25424]},
     {storeUnit_maskInput_lo[25423:25408]},
     {storeUnit_maskInput_lo[25407:25392]},
     {storeUnit_maskInput_lo[25391:25376]},
     {storeUnit_maskInput_lo[25375:25360]},
     {storeUnit_maskInput_lo[25359:25344]},
     {storeUnit_maskInput_lo[25343:25328]},
     {storeUnit_maskInput_lo[25327:25312]},
     {storeUnit_maskInput_lo[25311:25296]},
     {storeUnit_maskInput_lo[25295:25280]},
     {storeUnit_maskInput_lo[25279:25264]},
     {storeUnit_maskInput_lo[25263:25248]},
     {storeUnit_maskInput_lo[25247:25232]},
     {storeUnit_maskInput_lo[25231:25216]},
     {storeUnit_maskInput_lo[25215:25200]},
     {storeUnit_maskInput_lo[25199:25184]},
     {storeUnit_maskInput_lo[25183:25168]},
     {storeUnit_maskInput_lo[25167:25152]},
     {storeUnit_maskInput_lo[25151:25136]},
     {storeUnit_maskInput_lo[25135:25120]},
     {storeUnit_maskInput_lo[25119:25104]},
     {storeUnit_maskInput_lo[25103:25088]},
     {storeUnit_maskInput_lo[25087:25072]},
     {storeUnit_maskInput_lo[25071:25056]},
     {storeUnit_maskInput_lo[25055:25040]},
     {storeUnit_maskInput_lo[25039:25024]},
     {storeUnit_maskInput_lo[25023:25008]},
     {storeUnit_maskInput_lo[25007:24992]},
     {storeUnit_maskInput_lo[24991:24976]},
     {storeUnit_maskInput_lo[24975:24960]},
     {storeUnit_maskInput_lo[24959:24944]},
     {storeUnit_maskInput_lo[24943:24928]},
     {storeUnit_maskInput_lo[24927:24912]},
     {storeUnit_maskInput_lo[24911:24896]},
     {storeUnit_maskInput_lo[24895:24880]},
     {storeUnit_maskInput_lo[24879:24864]},
     {storeUnit_maskInput_lo[24863:24848]},
     {storeUnit_maskInput_lo[24847:24832]},
     {storeUnit_maskInput_lo[24831:24816]},
     {storeUnit_maskInput_lo[24815:24800]},
     {storeUnit_maskInput_lo[24799:24784]},
     {storeUnit_maskInput_lo[24783:24768]},
     {storeUnit_maskInput_lo[24767:24752]},
     {storeUnit_maskInput_lo[24751:24736]},
     {storeUnit_maskInput_lo[24735:24720]},
     {storeUnit_maskInput_lo[24719:24704]},
     {storeUnit_maskInput_lo[24703:24688]},
     {storeUnit_maskInput_lo[24687:24672]},
     {storeUnit_maskInput_lo[24671:24656]},
     {storeUnit_maskInput_lo[24655:24640]},
     {storeUnit_maskInput_lo[24639:24624]},
     {storeUnit_maskInput_lo[24623:24608]},
     {storeUnit_maskInput_lo[24607:24592]},
     {storeUnit_maskInput_lo[24591:24576]},
     {storeUnit_maskInput_lo[24575:24560]},
     {storeUnit_maskInput_lo[24559:24544]},
     {storeUnit_maskInput_lo[24543:24528]},
     {storeUnit_maskInput_lo[24527:24512]},
     {storeUnit_maskInput_lo[24511:24496]},
     {storeUnit_maskInput_lo[24495:24480]},
     {storeUnit_maskInput_lo[24479:24464]},
     {storeUnit_maskInput_lo[24463:24448]},
     {storeUnit_maskInput_lo[24447:24432]},
     {storeUnit_maskInput_lo[24431:24416]},
     {storeUnit_maskInput_lo[24415:24400]},
     {storeUnit_maskInput_lo[24399:24384]},
     {storeUnit_maskInput_lo[24383:24368]},
     {storeUnit_maskInput_lo[24367:24352]},
     {storeUnit_maskInput_lo[24351:24336]},
     {storeUnit_maskInput_lo[24335:24320]},
     {storeUnit_maskInput_lo[24319:24304]},
     {storeUnit_maskInput_lo[24303:24288]},
     {storeUnit_maskInput_lo[24287:24272]},
     {storeUnit_maskInput_lo[24271:24256]},
     {storeUnit_maskInput_lo[24255:24240]},
     {storeUnit_maskInput_lo[24239:24224]},
     {storeUnit_maskInput_lo[24223:24208]},
     {storeUnit_maskInput_lo[24207:24192]},
     {storeUnit_maskInput_lo[24191:24176]},
     {storeUnit_maskInput_lo[24175:24160]},
     {storeUnit_maskInput_lo[24159:24144]},
     {storeUnit_maskInput_lo[24143:24128]},
     {storeUnit_maskInput_lo[24127:24112]},
     {storeUnit_maskInput_lo[24111:24096]},
     {storeUnit_maskInput_lo[24095:24080]},
     {storeUnit_maskInput_lo[24079:24064]},
     {storeUnit_maskInput_lo[24063:24048]},
     {storeUnit_maskInput_lo[24047:24032]},
     {storeUnit_maskInput_lo[24031:24016]},
     {storeUnit_maskInput_lo[24015:24000]},
     {storeUnit_maskInput_lo[23999:23984]},
     {storeUnit_maskInput_lo[23983:23968]},
     {storeUnit_maskInput_lo[23967:23952]},
     {storeUnit_maskInput_lo[23951:23936]},
     {storeUnit_maskInput_lo[23935:23920]},
     {storeUnit_maskInput_lo[23919:23904]},
     {storeUnit_maskInput_lo[23903:23888]},
     {storeUnit_maskInput_lo[23887:23872]},
     {storeUnit_maskInput_lo[23871:23856]},
     {storeUnit_maskInput_lo[23855:23840]},
     {storeUnit_maskInput_lo[23839:23824]},
     {storeUnit_maskInput_lo[23823:23808]},
     {storeUnit_maskInput_lo[23807:23792]},
     {storeUnit_maskInput_lo[23791:23776]},
     {storeUnit_maskInput_lo[23775:23760]},
     {storeUnit_maskInput_lo[23759:23744]},
     {storeUnit_maskInput_lo[23743:23728]},
     {storeUnit_maskInput_lo[23727:23712]},
     {storeUnit_maskInput_lo[23711:23696]},
     {storeUnit_maskInput_lo[23695:23680]},
     {storeUnit_maskInput_lo[23679:23664]},
     {storeUnit_maskInput_lo[23663:23648]},
     {storeUnit_maskInput_lo[23647:23632]},
     {storeUnit_maskInput_lo[23631:23616]},
     {storeUnit_maskInput_lo[23615:23600]},
     {storeUnit_maskInput_lo[23599:23584]},
     {storeUnit_maskInput_lo[23583:23568]},
     {storeUnit_maskInput_lo[23567:23552]},
     {storeUnit_maskInput_lo[23551:23536]},
     {storeUnit_maskInput_lo[23535:23520]},
     {storeUnit_maskInput_lo[23519:23504]},
     {storeUnit_maskInput_lo[23503:23488]},
     {storeUnit_maskInput_lo[23487:23472]},
     {storeUnit_maskInput_lo[23471:23456]},
     {storeUnit_maskInput_lo[23455:23440]},
     {storeUnit_maskInput_lo[23439:23424]},
     {storeUnit_maskInput_lo[23423:23408]},
     {storeUnit_maskInput_lo[23407:23392]},
     {storeUnit_maskInput_lo[23391:23376]},
     {storeUnit_maskInput_lo[23375:23360]},
     {storeUnit_maskInput_lo[23359:23344]},
     {storeUnit_maskInput_lo[23343:23328]},
     {storeUnit_maskInput_lo[23327:23312]},
     {storeUnit_maskInput_lo[23311:23296]},
     {storeUnit_maskInput_lo[23295:23280]},
     {storeUnit_maskInput_lo[23279:23264]},
     {storeUnit_maskInput_lo[23263:23248]},
     {storeUnit_maskInput_lo[23247:23232]},
     {storeUnit_maskInput_lo[23231:23216]},
     {storeUnit_maskInput_lo[23215:23200]},
     {storeUnit_maskInput_lo[23199:23184]},
     {storeUnit_maskInput_lo[23183:23168]},
     {storeUnit_maskInput_lo[23167:23152]},
     {storeUnit_maskInput_lo[23151:23136]},
     {storeUnit_maskInput_lo[23135:23120]},
     {storeUnit_maskInput_lo[23119:23104]},
     {storeUnit_maskInput_lo[23103:23088]},
     {storeUnit_maskInput_lo[23087:23072]},
     {storeUnit_maskInput_lo[23071:23056]},
     {storeUnit_maskInput_lo[23055:23040]},
     {storeUnit_maskInput_lo[23039:23024]},
     {storeUnit_maskInput_lo[23023:23008]},
     {storeUnit_maskInput_lo[23007:22992]},
     {storeUnit_maskInput_lo[22991:22976]},
     {storeUnit_maskInput_lo[22975:22960]},
     {storeUnit_maskInput_lo[22959:22944]},
     {storeUnit_maskInput_lo[22943:22928]},
     {storeUnit_maskInput_lo[22927:22912]},
     {storeUnit_maskInput_lo[22911:22896]},
     {storeUnit_maskInput_lo[22895:22880]},
     {storeUnit_maskInput_lo[22879:22864]},
     {storeUnit_maskInput_lo[22863:22848]},
     {storeUnit_maskInput_lo[22847:22832]},
     {storeUnit_maskInput_lo[22831:22816]},
     {storeUnit_maskInput_lo[22815:22800]},
     {storeUnit_maskInput_lo[22799:22784]},
     {storeUnit_maskInput_lo[22783:22768]},
     {storeUnit_maskInput_lo[22767:22752]},
     {storeUnit_maskInput_lo[22751:22736]},
     {storeUnit_maskInput_lo[22735:22720]},
     {storeUnit_maskInput_lo[22719:22704]},
     {storeUnit_maskInput_lo[22703:22688]},
     {storeUnit_maskInput_lo[22687:22672]},
     {storeUnit_maskInput_lo[22671:22656]},
     {storeUnit_maskInput_lo[22655:22640]},
     {storeUnit_maskInput_lo[22639:22624]},
     {storeUnit_maskInput_lo[22623:22608]},
     {storeUnit_maskInput_lo[22607:22592]},
     {storeUnit_maskInput_lo[22591:22576]},
     {storeUnit_maskInput_lo[22575:22560]},
     {storeUnit_maskInput_lo[22559:22544]},
     {storeUnit_maskInput_lo[22543:22528]},
     {storeUnit_maskInput_lo[22527:22512]},
     {storeUnit_maskInput_lo[22511:22496]},
     {storeUnit_maskInput_lo[22495:22480]},
     {storeUnit_maskInput_lo[22479:22464]},
     {storeUnit_maskInput_lo[22463:22448]},
     {storeUnit_maskInput_lo[22447:22432]},
     {storeUnit_maskInput_lo[22431:22416]},
     {storeUnit_maskInput_lo[22415:22400]},
     {storeUnit_maskInput_lo[22399:22384]},
     {storeUnit_maskInput_lo[22383:22368]},
     {storeUnit_maskInput_lo[22367:22352]},
     {storeUnit_maskInput_lo[22351:22336]},
     {storeUnit_maskInput_lo[22335:22320]},
     {storeUnit_maskInput_lo[22319:22304]},
     {storeUnit_maskInput_lo[22303:22288]},
     {storeUnit_maskInput_lo[22287:22272]},
     {storeUnit_maskInput_lo[22271:22256]},
     {storeUnit_maskInput_lo[22255:22240]},
     {storeUnit_maskInput_lo[22239:22224]},
     {storeUnit_maskInput_lo[22223:22208]},
     {storeUnit_maskInput_lo[22207:22192]},
     {storeUnit_maskInput_lo[22191:22176]},
     {storeUnit_maskInput_lo[22175:22160]},
     {storeUnit_maskInput_lo[22159:22144]},
     {storeUnit_maskInput_lo[22143:22128]},
     {storeUnit_maskInput_lo[22127:22112]},
     {storeUnit_maskInput_lo[22111:22096]},
     {storeUnit_maskInput_lo[22095:22080]},
     {storeUnit_maskInput_lo[22079:22064]},
     {storeUnit_maskInput_lo[22063:22048]},
     {storeUnit_maskInput_lo[22047:22032]},
     {storeUnit_maskInput_lo[22031:22016]},
     {storeUnit_maskInput_lo[22015:22000]},
     {storeUnit_maskInput_lo[21999:21984]},
     {storeUnit_maskInput_lo[21983:21968]},
     {storeUnit_maskInput_lo[21967:21952]},
     {storeUnit_maskInput_lo[21951:21936]},
     {storeUnit_maskInput_lo[21935:21920]},
     {storeUnit_maskInput_lo[21919:21904]},
     {storeUnit_maskInput_lo[21903:21888]},
     {storeUnit_maskInput_lo[21887:21872]},
     {storeUnit_maskInput_lo[21871:21856]},
     {storeUnit_maskInput_lo[21855:21840]},
     {storeUnit_maskInput_lo[21839:21824]},
     {storeUnit_maskInput_lo[21823:21808]},
     {storeUnit_maskInput_lo[21807:21792]},
     {storeUnit_maskInput_lo[21791:21776]},
     {storeUnit_maskInput_lo[21775:21760]},
     {storeUnit_maskInput_lo[21759:21744]},
     {storeUnit_maskInput_lo[21743:21728]},
     {storeUnit_maskInput_lo[21727:21712]},
     {storeUnit_maskInput_lo[21711:21696]},
     {storeUnit_maskInput_lo[21695:21680]},
     {storeUnit_maskInput_lo[21679:21664]},
     {storeUnit_maskInput_lo[21663:21648]},
     {storeUnit_maskInput_lo[21647:21632]},
     {storeUnit_maskInput_lo[21631:21616]},
     {storeUnit_maskInput_lo[21615:21600]},
     {storeUnit_maskInput_lo[21599:21584]},
     {storeUnit_maskInput_lo[21583:21568]},
     {storeUnit_maskInput_lo[21567:21552]},
     {storeUnit_maskInput_lo[21551:21536]},
     {storeUnit_maskInput_lo[21535:21520]},
     {storeUnit_maskInput_lo[21519:21504]},
     {storeUnit_maskInput_lo[21503:21488]},
     {storeUnit_maskInput_lo[21487:21472]},
     {storeUnit_maskInput_lo[21471:21456]},
     {storeUnit_maskInput_lo[21455:21440]},
     {storeUnit_maskInput_lo[21439:21424]},
     {storeUnit_maskInput_lo[21423:21408]},
     {storeUnit_maskInput_lo[21407:21392]},
     {storeUnit_maskInput_lo[21391:21376]},
     {storeUnit_maskInput_lo[21375:21360]},
     {storeUnit_maskInput_lo[21359:21344]},
     {storeUnit_maskInput_lo[21343:21328]},
     {storeUnit_maskInput_lo[21327:21312]},
     {storeUnit_maskInput_lo[21311:21296]},
     {storeUnit_maskInput_lo[21295:21280]},
     {storeUnit_maskInput_lo[21279:21264]},
     {storeUnit_maskInput_lo[21263:21248]},
     {storeUnit_maskInput_lo[21247:21232]},
     {storeUnit_maskInput_lo[21231:21216]},
     {storeUnit_maskInput_lo[21215:21200]},
     {storeUnit_maskInput_lo[21199:21184]},
     {storeUnit_maskInput_lo[21183:21168]},
     {storeUnit_maskInput_lo[21167:21152]},
     {storeUnit_maskInput_lo[21151:21136]},
     {storeUnit_maskInput_lo[21135:21120]},
     {storeUnit_maskInput_lo[21119:21104]},
     {storeUnit_maskInput_lo[21103:21088]},
     {storeUnit_maskInput_lo[21087:21072]},
     {storeUnit_maskInput_lo[21071:21056]},
     {storeUnit_maskInput_lo[21055:21040]},
     {storeUnit_maskInput_lo[21039:21024]},
     {storeUnit_maskInput_lo[21023:21008]},
     {storeUnit_maskInput_lo[21007:20992]},
     {storeUnit_maskInput_lo[20991:20976]},
     {storeUnit_maskInput_lo[20975:20960]},
     {storeUnit_maskInput_lo[20959:20944]},
     {storeUnit_maskInput_lo[20943:20928]},
     {storeUnit_maskInput_lo[20927:20912]},
     {storeUnit_maskInput_lo[20911:20896]},
     {storeUnit_maskInput_lo[20895:20880]},
     {storeUnit_maskInput_lo[20879:20864]},
     {storeUnit_maskInput_lo[20863:20848]},
     {storeUnit_maskInput_lo[20847:20832]},
     {storeUnit_maskInput_lo[20831:20816]},
     {storeUnit_maskInput_lo[20815:20800]},
     {storeUnit_maskInput_lo[20799:20784]},
     {storeUnit_maskInput_lo[20783:20768]},
     {storeUnit_maskInput_lo[20767:20752]},
     {storeUnit_maskInput_lo[20751:20736]},
     {storeUnit_maskInput_lo[20735:20720]},
     {storeUnit_maskInput_lo[20719:20704]},
     {storeUnit_maskInput_lo[20703:20688]},
     {storeUnit_maskInput_lo[20687:20672]},
     {storeUnit_maskInput_lo[20671:20656]},
     {storeUnit_maskInput_lo[20655:20640]},
     {storeUnit_maskInput_lo[20639:20624]},
     {storeUnit_maskInput_lo[20623:20608]},
     {storeUnit_maskInput_lo[20607:20592]},
     {storeUnit_maskInput_lo[20591:20576]},
     {storeUnit_maskInput_lo[20575:20560]},
     {storeUnit_maskInput_lo[20559:20544]},
     {storeUnit_maskInput_lo[20543:20528]},
     {storeUnit_maskInput_lo[20527:20512]},
     {storeUnit_maskInput_lo[20511:20496]},
     {storeUnit_maskInput_lo[20495:20480]},
     {storeUnit_maskInput_lo[20479:20464]},
     {storeUnit_maskInput_lo[20463:20448]},
     {storeUnit_maskInput_lo[20447:20432]},
     {storeUnit_maskInput_lo[20431:20416]},
     {storeUnit_maskInput_lo[20415:20400]},
     {storeUnit_maskInput_lo[20399:20384]},
     {storeUnit_maskInput_lo[20383:20368]},
     {storeUnit_maskInput_lo[20367:20352]},
     {storeUnit_maskInput_lo[20351:20336]},
     {storeUnit_maskInput_lo[20335:20320]},
     {storeUnit_maskInput_lo[20319:20304]},
     {storeUnit_maskInput_lo[20303:20288]},
     {storeUnit_maskInput_lo[20287:20272]},
     {storeUnit_maskInput_lo[20271:20256]},
     {storeUnit_maskInput_lo[20255:20240]},
     {storeUnit_maskInput_lo[20239:20224]},
     {storeUnit_maskInput_lo[20223:20208]},
     {storeUnit_maskInput_lo[20207:20192]},
     {storeUnit_maskInput_lo[20191:20176]},
     {storeUnit_maskInput_lo[20175:20160]},
     {storeUnit_maskInput_lo[20159:20144]},
     {storeUnit_maskInput_lo[20143:20128]},
     {storeUnit_maskInput_lo[20127:20112]},
     {storeUnit_maskInput_lo[20111:20096]},
     {storeUnit_maskInput_lo[20095:20080]},
     {storeUnit_maskInput_lo[20079:20064]},
     {storeUnit_maskInput_lo[20063:20048]},
     {storeUnit_maskInput_lo[20047:20032]},
     {storeUnit_maskInput_lo[20031:20016]},
     {storeUnit_maskInput_lo[20015:20000]},
     {storeUnit_maskInput_lo[19999:19984]},
     {storeUnit_maskInput_lo[19983:19968]},
     {storeUnit_maskInput_lo[19967:19952]},
     {storeUnit_maskInput_lo[19951:19936]},
     {storeUnit_maskInput_lo[19935:19920]},
     {storeUnit_maskInput_lo[19919:19904]},
     {storeUnit_maskInput_lo[19903:19888]},
     {storeUnit_maskInput_lo[19887:19872]},
     {storeUnit_maskInput_lo[19871:19856]},
     {storeUnit_maskInput_lo[19855:19840]},
     {storeUnit_maskInput_lo[19839:19824]},
     {storeUnit_maskInput_lo[19823:19808]},
     {storeUnit_maskInput_lo[19807:19792]},
     {storeUnit_maskInput_lo[19791:19776]},
     {storeUnit_maskInput_lo[19775:19760]},
     {storeUnit_maskInput_lo[19759:19744]},
     {storeUnit_maskInput_lo[19743:19728]},
     {storeUnit_maskInput_lo[19727:19712]},
     {storeUnit_maskInput_lo[19711:19696]},
     {storeUnit_maskInput_lo[19695:19680]},
     {storeUnit_maskInput_lo[19679:19664]},
     {storeUnit_maskInput_lo[19663:19648]},
     {storeUnit_maskInput_lo[19647:19632]},
     {storeUnit_maskInput_lo[19631:19616]},
     {storeUnit_maskInput_lo[19615:19600]},
     {storeUnit_maskInput_lo[19599:19584]},
     {storeUnit_maskInput_lo[19583:19568]},
     {storeUnit_maskInput_lo[19567:19552]},
     {storeUnit_maskInput_lo[19551:19536]},
     {storeUnit_maskInput_lo[19535:19520]},
     {storeUnit_maskInput_lo[19519:19504]},
     {storeUnit_maskInput_lo[19503:19488]},
     {storeUnit_maskInput_lo[19487:19472]},
     {storeUnit_maskInput_lo[19471:19456]},
     {storeUnit_maskInput_lo[19455:19440]},
     {storeUnit_maskInput_lo[19439:19424]},
     {storeUnit_maskInput_lo[19423:19408]},
     {storeUnit_maskInput_lo[19407:19392]},
     {storeUnit_maskInput_lo[19391:19376]},
     {storeUnit_maskInput_lo[19375:19360]},
     {storeUnit_maskInput_lo[19359:19344]},
     {storeUnit_maskInput_lo[19343:19328]},
     {storeUnit_maskInput_lo[19327:19312]},
     {storeUnit_maskInput_lo[19311:19296]},
     {storeUnit_maskInput_lo[19295:19280]},
     {storeUnit_maskInput_lo[19279:19264]},
     {storeUnit_maskInput_lo[19263:19248]},
     {storeUnit_maskInput_lo[19247:19232]},
     {storeUnit_maskInput_lo[19231:19216]},
     {storeUnit_maskInput_lo[19215:19200]},
     {storeUnit_maskInput_lo[19199:19184]},
     {storeUnit_maskInput_lo[19183:19168]},
     {storeUnit_maskInput_lo[19167:19152]},
     {storeUnit_maskInput_lo[19151:19136]},
     {storeUnit_maskInput_lo[19135:19120]},
     {storeUnit_maskInput_lo[19119:19104]},
     {storeUnit_maskInput_lo[19103:19088]},
     {storeUnit_maskInput_lo[19087:19072]},
     {storeUnit_maskInput_lo[19071:19056]},
     {storeUnit_maskInput_lo[19055:19040]},
     {storeUnit_maskInput_lo[19039:19024]},
     {storeUnit_maskInput_lo[19023:19008]},
     {storeUnit_maskInput_lo[19007:18992]},
     {storeUnit_maskInput_lo[18991:18976]},
     {storeUnit_maskInput_lo[18975:18960]},
     {storeUnit_maskInput_lo[18959:18944]},
     {storeUnit_maskInput_lo[18943:18928]},
     {storeUnit_maskInput_lo[18927:18912]},
     {storeUnit_maskInput_lo[18911:18896]},
     {storeUnit_maskInput_lo[18895:18880]},
     {storeUnit_maskInput_lo[18879:18864]},
     {storeUnit_maskInput_lo[18863:18848]},
     {storeUnit_maskInput_lo[18847:18832]},
     {storeUnit_maskInput_lo[18831:18816]},
     {storeUnit_maskInput_lo[18815:18800]},
     {storeUnit_maskInput_lo[18799:18784]},
     {storeUnit_maskInput_lo[18783:18768]},
     {storeUnit_maskInput_lo[18767:18752]},
     {storeUnit_maskInput_lo[18751:18736]},
     {storeUnit_maskInput_lo[18735:18720]},
     {storeUnit_maskInput_lo[18719:18704]},
     {storeUnit_maskInput_lo[18703:18688]},
     {storeUnit_maskInput_lo[18687:18672]},
     {storeUnit_maskInput_lo[18671:18656]},
     {storeUnit_maskInput_lo[18655:18640]},
     {storeUnit_maskInput_lo[18639:18624]},
     {storeUnit_maskInput_lo[18623:18608]},
     {storeUnit_maskInput_lo[18607:18592]},
     {storeUnit_maskInput_lo[18591:18576]},
     {storeUnit_maskInput_lo[18575:18560]},
     {storeUnit_maskInput_lo[18559:18544]},
     {storeUnit_maskInput_lo[18543:18528]},
     {storeUnit_maskInput_lo[18527:18512]},
     {storeUnit_maskInput_lo[18511:18496]},
     {storeUnit_maskInput_lo[18495:18480]},
     {storeUnit_maskInput_lo[18479:18464]},
     {storeUnit_maskInput_lo[18463:18448]},
     {storeUnit_maskInput_lo[18447:18432]},
     {storeUnit_maskInput_lo[18431:18416]},
     {storeUnit_maskInput_lo[18415:18400]},
     {storeUnit_maskInput_lo[18399:18384]},
     {storeUnit_maskInput_lo[18383:18368]},
     {storeUnit_maskInput_lo[18367:18352]},
     {storeUnit_maskInput_lo[18351:18336]},
     {storeUnit_maskInput_lo[18335:18320]},
     {storeUnit_maskInput_lo[18319:18304]},
     {storeUnit_maskInput_lo[18303:18288]},
     {storeUnit_maskInput_lo[18287:18272]},
     {storeUnit_maskInput_lo[18271:18256]},
     {storeUnit_maskInput_lo[18255:18240]},
     {storeUnit_maskInput_lo[18239:18224]},
     {storeUnit_maskInput_lo[18223:18208]},
     {storeUnit_maskInput_lo[18207:18192]},
     {storeUnit_maskInput_lo[18191:18176]},
     {storeUnit_maskInput_lo[18175:18160]},
     {storeUnit_maskInput_lo[18159:18144]},
     {storeUnit_maskInput_lo[18143:18128]},
     {storeUnit_maskInput_lo[18127:18112]},
     {storeUnit_maskInput_lo[18111:18096]},
     {storeUnit_maskInput_lo[18095:18080]},
     {storeUnit_maskInput_lo[18079:18064]},
     {storeUnit_maskInput_lo[18063:18048]},
     {storeUnit_maskInput_lo[18047:18032]},
     {storeUnit_maskInput_lo[18031:18016]},
     {storeUnit_maskInput_lo[18015:18000]},
     {storeUnit_maskInput_lo[17999:17984]},
     {storeUnit_maskInput_lo[17983:17968]},
     {storeUnit_maskInput_lo[17967:17952]},
     {storeUnit_maskInput_lo[17951:17936]},
     {storeUnit_maskInput_lo[17935:17920]},
     {storeUnit_maskInput_lo[17919:17904]},
     {storeUnit_maskInput_lo[17903:17888]},
     {storeUnit_maskInput_lo[17887:17872]},
     {storeUnit_maskInput_lo[17871:17856]},
     {storeUnit_maskInput_lo[17855:17840]},
     {storeUnit_maskInput_lo[17839:17824]},
     {storeUnit_maskInput_lo[17823:17808]},
     {storeUnit_maskInput_lo[17807:17792]},
     {storeUnit_maskInput_lo[17791:17776]},
     {storeUnit_maskInput_lo[17775:17760]},
     {storeUnit_maskInput_lo[17759:17744]},
     {storeUnit_maskInput_lo[17743:17728]},
     {storeUnit_maskInput_lo[17727:17712]},
     {storeUnit_maskInput_lo[17711:17696]},
     {storeUnit_maskInput_lo[17695:17680]},
     {storeUnit_maskInput_lo[17679:17664]},
     {storeUnit_maskInput_lo[17663:17648]},
     {storeUnit_maskInput_lo[17647:17632]},
     {storeUnit_maskInput_lo[17631:17616]},
     {storeUnit_maskInput_lo[17615:17600]},
     {storeUnit_maskInput_lo[17599:17584]},
     {storeUnit_maskInput_lo[17583:17568]},
     {storeUnit_maskInput_lo[17567:17552]},
     {storeUnit_maskInput_lo[17551:17536]},
     {storeUnit_maskInput_lo[17535:17520]},
     {storeUnit_maskInput_lo[17519:17504]},
     {storeUnit_maskInput_lo[17503:17488]},
     {storeUnit_maskInput_lo[17487:17472]},
     {storeUnit_maskInput_lo[17471:17456]},
     {storeUnit_maskInput_lo[17455:17440]},
     {storeUnit_maskInput_lo[17439:17424]},
     {storeUnit_maskInput_lo[17423:17408]},
     {storeUnit_maskInput_lo[17407:17392]},
     {storeUnit_maskInput_lo[17391:17376]},
     {storeUnit_maskInput_lo[17375:17360]},
     {storeUnit_maskInput_lo[17359:17344]},
     {storeUnit_maskInput_lo[17343:17328]},
     {storeUnit_maskInput_lo[17327:17312]},
     {storeUnit_maskInput_lo[17311:17296]},
     {storeUnit_maskInput_lo[17295:17280]},
     {storeUnit_maskInput_lo[17279:17264]},
     {storeUnit_maskInput_lo[17263:17248]},
     {storeUnit_maskInput_lo[17247:17232]},
     {storeUnit_maskInput_lo[17231:17216]},
     {storeUnit_maskInput_lo[17215:17200]},
     {storeUnit_maskInput_lo[17199:17184]},
     {storeUnit_maskInput_lo[17183:17168]},
     {storeUnit_maskInput_lo[17167:17152]},
     {storeUnit_maskInput_lo[17151:17136]},
     {storeUnit_maskInput_lo[17135:17120]},
     {storeUnit_maskInput_lo[17119:17104]},
     {storeUnit_maskInput_lo[17103:17088]},
     {storeUnit_maskInput_lo[17087:17072]},
     {storeUnit_maskInput_lo[17071:17056]},
     {storeUnit_maskInput_lo[17055:17040]},
     {storeUnit_maskInput_lo[17039:17024]},
     {storeUnit_maskInput_lo[17023:17008]},
     {storeUnit_maskInput_lo[17007:16992]},
     {storeUnit_maskInput_lo[16991:16976]},
     {storeUnit_maskInput_lo[16975:16960]},
     {storeUnit_maskInput_lo[16959:16944]},
     {storeUnit_maskInput_lo[16943:16928]},
     {storeUnit_maskInput_lo[16927:16912]},
     {storeUnit_maskInput_lo[16911:16896]},
     {storeUnit_maskInput_lo[16895:16880]},
     {storeUnit_maskInput_lo[16879:16864]},
     {storeUnit_maskInput_lo[16863:16848]},
     {storeUnit_maskInput_lo[16847:16832]},
     {storeUnit_maskInput_lo[16831:16816]},
     {storeUnit_maskInput_lo[16815:16800]},
     {storeUnit_maskInput_lo[16799:16784]},
     {storeUnit_maskInput_lo[16783:16768]},
     {storeUnit_maskInput_lo[16767:16752]},
     {storeUnit_maskInput_lo[16751:16736]},
     {storeUnit_maskInput_lo[16735:16720]},
     {storeUnit_maskInput_lo[16719:16704]},
     {storeUnit_maskInput_lo[16703:16688]},
     {storeUnit_maskInput_lo[16687:16672]},
     {storeUnit_maskInput_lo[16671:16656]},
     {storeUnit_maskInput_lo[16655:16640]},
     {storeUnit_maskInput_lo[16639:16624]},
     {storeUnit_maskInput_lo[16623:16608]},
     {storeUnit_maskInput_lo[16607:16592]},
     {storeUnit_maskInput_lo[16591:16576]},
     {storeUnit_maskInput_lo[16575:16560]},
     {storeUnit_maskInput_lo[16559:16544]},
     {storeUnit_maskInput_lo[16543:16528]},
     {storeUnit_maskInput_lo[16527:16512]},
     {storeUnit_maskInput_lo[16511:16496]},
     {storeUnit_maskInput_lo[16495:16480]},
     {storeUnit_maskInput_lo[16479:16464]},
     {storeUnit_maskInput_lo[16463:16448]},
     {storeUnit_maskInput_lo[16447:16432]},
     {storeUnit_maskInput_lo[16431:16416]},
     {storeUnit_maskInput_lo[16415:16400]},
     {storeUnit_maskInput_lo[16399:16384]},
     {storeUnit_maskInput_lo[16383:16368]},
     {storeUnit_maskInput_lo[16367:16352]},
     {storeUnit_maskInput_lo[16351:16336]},
     {storeUnit_maskInput_lo[16335:16320]},
     {storeUnit_maskInput_lo[16319:16304]},
     {storeUnit_maskInput_lo[16303:16288]},
     {storeUnit_maskInput_lo[16287:16272]},
     {storeUnit_maskInput_lo[16271:16256]},
     {storeUnit_maskInput_lo[16255:16240]},
     {storeUnit_maskInput_lo[16239:16224]},
     {storeUnit_maskInput_lo[16223:16208]},
     {storeUnit_maskInput_lo[16207:16192]},
     {storeUnit_maskInput_lo[16191:16176]},
     {storeUnit_maskInput_lo[16175:16160]},
     {storeUnit_maskInput_lo[16159:16144]},
     {storeUnit_maskInput_lo[16143:16128]},
     {storeUnit_maskInput_lo[16127:16112]},
     {storeUnit_maskInput_lo[16111:16096]},
     {storeUnit_maskInput_lo[16095:16080]},
     {storeUnit_maskInput_lo[16079:16064]},
     {storeUnit_maskInput_lo[16063:16048]},
     {storeUnit_maskInput_lo[16047:16032]},
     {storeUnit_maskInput_lo[16031:16016]},
     {storeUnit_maskInput_lo[16015:16000]},
     {storeUnit_maskInput_lo[15999:15984]},
     {storeUnit_maskInput_lo[15983:15968]},
     {storeUnit_maskInput_lo[15967:15952]},
     {storeUnit_maskInput_lo[15951:15936]},
     {storeUnit_maskInput_lo[15935:15920]},
     {storeUnit_maskInput_lo[15919:15904]},
     {storeUnit_maskInput_lo[15903:15888]},
     {storeUnit_maskInput_lo[15887:15872]},
     {storeUnit_maskInput_lo[15871:15856]},
     {storeUnit_maskInput_lo[15855:15840]},
     {storeUnit_maskInput_lo[15839:15824]},
     {storeUnit_maskInput_lo[15823:15808]},
     {storeUnit_maskInput_lo[15807:15792]},
     {storeUnit_maskInput_lo[15791:15776]},
     {storeUnit_maskInput_lo[15775:15760]},
     {storeUnit_maskInput_lo[15759:15744]},
     {storeUnit_maskInput_lo[15743:15728]},
     {storeUnit_maskInput_lo[15727:15712]},
     {storeUnit_maskInput_lo[15711:15696]},
     {storeUnit_maskInput_lo[15695:15680]},
     {storeUnit_maskInput_lo[15679:15664]},
     {storeUnit_maskInput_lo[15663:15648]},
     {storeUnit_maskInput_lo[15647:15632]},
     {storeUnit_maskInput_lo[15631:15616]},
     {storeUnit_maskInput_lo[15615:15600]},
     {storeUnit_maskInput_lo[15599:15584]},
     {storeUnit_maskInput_lo[15583:15568]},
     {storeUnit_maskInput_lo[15567:15552]},
     {storeUnit_maskInput_lo[15551:15536]},
     {storeUnit_maskInput_lo[15535:15520]},
     {storeUnit_maskInput_lo[15519:15504]},
     {storeUnit_maskInput_lo[15503:15488]},
     {storeUnit_maskInput_lo[15487:15472]},
     {storeUnit_maskInput_lo[15471:15456]},
     {storeUnit_maskInput_lo[15455:15440]},
     {storeUnit_maskInput_lo[15439:15424]},
     {storeUnit_maskInput_lo[15423:15408]},
     {storeUnit_maskInput_lo[15407:15392]},
     {storeUnit_maskInput_lo[15391:15376]},
     {storeUnit_maskInput_lo[15375:15360]},
     {storeUnit_maskInput_lo[15359:15344]},
     {storeUnit_maskInput_lo[15343:15328]},
     {storeUnit_maskInput_lo[15327:15312]},
     {storeUnit_maskInput_lo[15311:15296]},
     {storeUnit_maskInput_lo[15295:15280]},
     {storeUnit_maskInput_lo[15279:15264]},
     {storeUnit_maskInput_lo[15263:15248]},
     {storeUnit_maskInput_lo[15247:15232]},
     {storeUnit_maskInput_lo[15231:15216]},
     {storeUnit_maskInput_lo[15215:15200]},
     {storeUnit_maskInput_lo[15199:15184]},
     {storeUnit_maskInput_lo[15183:15168]},
     {storeUnit_maskInput_lo[15167:15152]},
     {storeUnit_maskInput_lo[15151:15136]},
     {storeUnit_maskInput_lo[15135:15120]},
     {storeUnit_maskInput_lo[15119:15104]},
     {storeUnit_maskInput_lo[15103:15088]},
     {storeUnit_maskInput_lo[15087:15072]},
     {storeUnit_maskInput_lo[15071:15056]},
     {storeUnit_maskInput_lo[15055:15040]},
     {storeUnit_maskInput_lo[15039:15024]},
     {storeUnit_maskInput_lo[15023:15008]},
     {storeUnit_maskInput_lo[15007:14992]},
     {storeUnit_maskInput_lo[14991:14976]},
     {storeUnit_maskInput_lo[14975:14960]},
     {storeUnit_maskInput_lo[14959:14944]},
     {storeUnit_maskInput_lo[14943:14928]},
     {storeUnit_maskInput_lo[14927:14912]},
     {storeUnit_maskInput_lo[14911:14896]},
     {storeUnit_maskInput_lo[14895:14880]},
     {storeUnit_maskInput_lo[14879:14864]},
     {storeUnit_maskInput_lo[14863:14848]},
     {storeUnit_maskInput_lo[14847:14832]},
     {storeUnit_maskInput_lo[14831:14816]},
     {storeUnit_maskInput_lo[14815:14800]},
     {storeUnit_maskInput_lo[14799:14784]},
     {storeUnit_maskInput_lo[14783:14768]},
     {storeUnit_maskInput_lo[14767:14752]},
     {storeUnit_maskInput_lo[14751:14736]},
     {storeUnit_maskInput_lo[14735:14720]},
     {storeUnit_maskInput_lo[14719:14704]},
     {storeUnit_maskInput_lo[14703:14688]},
     {storeUnit_maskInput_lo[14687:14672]},
     {storeUnit_maskInput_lo[14671:14656]},
     {storeUnit_maskInput_lo[14655:14640]},
     {storeUnit_maskInput_lo[14639:14624]},
     {storeUnit_maskInput_lo[14623:14608]},
     {storeUnit_maskInput_lo[14607:14592]},
     {storeUnit_maskInput_lo[14591:14576]},
     {storeUnit_maskInput_lo[14575:14560]},
     {storeUnit_maskInput_lo[14559:14544]},
     {storeUnit_maskInput_lo[14543:14528]},
     {storeUnit_maskInput_lo[14527:14512]},
     {storeUnit_maskInput_lo[14511:14496]},
     {storeUnit_maskInput_lo[14495:14480]},
     {storeUnit_maskInput_lo[14479:14464]},
     {storeUnit_maskInput_lo[14463:14448]},
     {storeUnit_maskInput_lo[14447:14432]},
     {storeUnit_maskInput_lo[14431:14416]},
     {storeUnit_maskInput_lo[14415:14400]},
     {storeUnit_maskInput_lo[14399:14384]},
     {storeUnit_maskInput_lo[14383:14368]},
     {storeUnit_maskInput_lo[14367:14352]},
     {storeUnit_maskInput_lo[14351:14336]},
     {storeUnit_maskInput_lo[14335:14320]},
     {storeUnit_maskInput_lo[14319:14304]},
     {storeUnit_maskInput_lo[14303:14288]},
     {storeUnit_maskInput_lo[14287:14272]},
     {storeUnit_maskInput_lo[14271:14256]},
     {storeUnit_maskInput_lo[14255:14240]},
     {storeUnit_maskInput_lo[14239:14224]},
     {storeUnit_maskInput_lo[14223:14208]},
     {storeUnit_maskInput_lo[14207:14192]},
     {storeUnit_maskInput_lo[14191:14176]},
     {storeUnit_maskInput_lo[14175:14160]},
     {storeUnit_maskInput_lo[14159:14144]},
     {storeUnit_maskInput_lo[14143:14128]},
     {storeUnit_maskInput_lo[14127:14112]},
     {storeUnit_maskInput_lo[14111:14096]},
     {storeUnit_maskInput_lo[14095:14080]},
     {storeUnit_maskInput_lo[14079:14064]},
     {storeUnit_maskInput_lo[14063:14048]},
     {storeUnit_maskInput_lo[14047:14032]},
     {storeUnit_maskInput_lo[14031:14016]},
     {storeUnit_maskInput_lo[14015:14000]},
     {storeUnit_maskInput_lo[13999:13984]},
     {storeUnit_maskInput_lo[13983:13968]},
     {storeUnit_maskInput_lo[13967:13952]},
     {storeUnit_maskInput_lo[13951:13936]},
     {storeUnit_maskInput_lo[13935:13920]},
     {storeUnit_maskInput_lo[13919:13904]},
     {storeUnit_maskInput_lo[13903:13888]},
     {storeUnit_maskInput_lo[13887:13872]},
     {storeUnit_maskInput_lo[13871:13856]},
     {storeUnit_maskInput_lo[13855:13840]},
     {storeUnit_maskInput_lo[13839:13824]},
     {storeUnit_maskInput_lo[13823:13808]},
     {storeUnit_maskInput_lo[13807:13792]},
     {storeUnit_maskInput_lo[13791:13776]},
     {storeUnit_maskInput_lo[13775:13760]},
     {storeUnit_maskInput_lo[13759:13744]},
     {storeUnit_maskInput_lo[13743:13728]},
     {storeUnit_maskInput_lo[13727:13712]},
     {storeUnit_maskInput_lo[13711:13696]},
     {storeUnit_maskInput_lo[13695:13680]},
     {storeUnit_maskInput_lo[13679:13664]},
     {storeUnit_maskInput_lo[13663:13648]},
     {storeUnit_maskInput_lo[13647:13632]},
     {storeUnit_maskInput_lo[13631:13616]},
     {storeUnit_maskInput_lo[13615:13600]},
     {storeUnit_maskInput_lo[13599:13584]},
     {storeUnit_maskInput_lo[13583:13568]},
     {storeUnit_maskInput_lo[13567:13552]},
     {storeUnit_maskInput_lo[13551:13536]},
     {storeUnit_maskInput_lo[13535:13520]},
     {storeUnit_maskInput_lo[13519:13504]},
     {storeUnit_maskInput_lo[13503:13488]},
     {storeUnit_maskInput_lo[13487:13472]},
     {storeUnit_maskInput_lo[13471:13456]},
     {storeUnit_maskInput_lo[13455:13440]},
     {storeUnit_maskInput_lo[13439:13424]},
     {storeUnit_maskInput_lo[13423:13408]},
     {storeUnit_maskInput_lo[13407:13392]},
     {storeUnit_maskInput_lo[13391:13376]},
     {storeUnit_maskInput_lo[13375:13360]},
     {storeUnit_maskInput_lo[13359:13344]},
     {storeUnit_maskInput_lo[13343:13328]},
     {storeUnit_maskInput_lo[13327:13312]},
     {storeUnit_maskInput_lo[13311:13296]},
     {storeUnit_maskInput_lo[13295:13280]},
     {storeUnit_maskInput_lo[13279:13264]},
     {storeUnit_maskInput_lo[13263:13248]},
     {storeUnit_maskInput_lo[13247:13232]},
     {storeUnit_maskInput_lo[13231:13216]},
     {storeUnit_maskInput_lo[13215:13200]},
     {storeUnit_maskInput_lo[13199:13184]},
     {storeUnit_maskInput_lo[13183:13168]},
     {storeUnit_maskInput_lo[13167:13152]},
     {storeUnit_maskInput_lo[13151:13136]},
     {storeUnit_maskInput_lo[13135:13120]},
     {storeUnit_maskInput_lo[13119:13104]},
     {storeUnit_maskInput_lo[13103:13088]},
     {storeUnit_maskInput_lo[13087:13072]},
     {storeUnit_maskInput_lo[13071:13056]},
     {storeUnit_maskInput_lo[13055:13040]},
     {storeUnit_maskInput_lo[13039:13024]},
     {storeUnit_maskInput_lo[13023:13008]},
     {storeUnit_maskInput_lo[13007:12992]},
     {storeUnit_maskInput_lo[12991:12976]},
     {storeUnit_maskInput_lo[12975:12960]},
     {storeUnit_maskInput_lo[12959:12944]},
     {storeUnit_maskInput_lo[12943:12928]},
     {storeUnit_maskInput_lo[12927:12912]},
     {storeUnit_maskInput_lo[12911:12896]},
     {storeUnit_maskInput_lo[12895:12880]},
     {storeUnit_maskInput_lo[12879:12864]},
     {storeUnit_maskInput_lo[12863:12848]},
     {storeUnit_maskInput_lo[12847:12832]},
     {storeUnit_maskInput_lo[12831:12816]},
     {storeUnit_maskInput_lo[12815:12800]},
     {storeUnit_maskInput_lo[12799:12784]},
     {storeUnit_maskInput_lo[12783:12768]},
     {storeUnit_maskInput_lo[12767:12752]},
     {storeUnit_maskInput_lo[12751:12736]},
     {storeUnit_maskInput_lo[12735:12720]},
     {storeUnit_maskInput_lo[12719:12704]},
     {storeUnit_maskInput_lo[12703:12688]},
     {storeUnit_maskInput_lo[12687:12672]},
     {storeUnit_maskInput_lo[12671:12656]},
     {storeUnit_maskInput_lo[12655:12640]},
     {storeUnit_maskInput_lo[12639:12624]},
     {storeUnit_maskInput_lo[12623:12608]},
     {storeUnit_maskInput_lo[12607:12592]},
     {storeUnit_maskInput_lo[12591:12576]},
     {storeUnit_maskInput_lo[12575:12560]},
     {storeUnit_maskInput_lo[12559:12544]},
     {storeUnit_maskInput_lo[12543:12528]},
     {storeUnit_maskInput_lo[12527:12512]},
     {storeUnit_maskInput_lo[12511:12496]},
     {storeUnit_maskInput_lo[12495:12480]},
     {storeUnit_maskInput_lo[12479:12464]},
     {storeUnit_maskInput_lo[12463:12448]},
     {storeUnit_maskInput_lo[12447:12432]},
     {storeUnit_maskInput_lo[12431:12416]},
     {storeUnit_maskInput_lo[12415:12400]},
     {storeUnit_maskInput_lo[12399:12384]},
     {storeUnit_maskInput_lo[12383:12368]},
     {storeUnit_maskInput_lo[12367:12352]},
     {storeUnit_maskInput_lo[12351:12336]},
     {storeUnit_maskInput_lo[12335:12320]},
     {storeUnit_maskInput_lo[12319:12304]},
     {storeUnit_maskInput_lo[12303:12288]},
     {storeUnit_maskInput_lo[12287:12272]},
     {storeUnit_maskInput_lo[12271:12256]},
     {storeUnit_maskInput_lo[12255:12240]},
     {storeUnit_maskInput_lo[12239:12224]},
     {storeUnit_maskInput_lo[12223:12208]},
     {storeUnit_maskInput_lo[12207:12192]},
     {storeUnit_maskInput_lo[12191:12176]},
     {storeUnit_maskInput_lo[12175:12160]},
     {storeUnit_maskInput_lo[12159:12144]},
     {storeUnit_maskInput_lo[12143:12128]},
     {storeUnit_maskInput_lo[12127:12112]},
     {storeUnit_maskInput_lo[12111:12096]},
     {storeUnit_maskInput_lo[12095:12080]},
     {storeUnit_maskInput_lo[12079:12064]},
     {storeUnit_maskInput_lo[12063:12048]},
     {storeUnit_maskInput_lo[12047:12032]},
     {storeUnit_maskInput_lo[12031:12016]},
     {storeUnit_maskInput_lo[12015:12000]},
     {storeUnit_maskInput_lo[11999:11984]},
     {storeUnit_maskInput_lo[11983:11968]},
     {storeUnit_maskInput_lo[11967:11952]},
     {storeUnit_maskInput_lo[11951:11936]},
     {storeUnit_maskInput_lo[11935:11920]},
     {storeUnit_maskInput_lo[11919:11904]},
     {storeUnit_maskInput_lo[11903:11888]},
     {storeUnit_maskInput_lo[11887:11872]},
     {storeUnit_maskInput_lo[11871:11856]},
     {storeUnit_maskInput_lo[11855:11840]},
     {storeUnit_maskInput_lo[11839:11824]},
     {storeUnit_maskInput_lo[11823:11808]},
     {storeUnit_maskInput_lo[11807:11792]},
     {storeUnit_maskInput_lo[11791:11776]},
     {storeUnit_maskInput_lo[11775:11760]},
     {storeUnit_maskInput_lo[11759:11744]},
     {storeUnit_maskInput_lo[11743:11728]},
     {storeUnit_maskInput_lo[11727:11712]},
     {storeUnit_maskInput_lo[11711:11696]},
     {storeUnit_maskInput_lo[11695:11680]},
     {storeUnit_maskInput_lo[11679:11664]},
     {storeUnit_maskInput_lo[11663:11648]},
     {storeUnit_maskInput_lo[11647:11632]},
     {storeUnit_maskInput_lo[11631:11616]},
     {storeUnit_maskInput_lo[11615:11600]},
     {storeUnit_maskInput_lo[11599:11584]},
     {storeUnit_maskInput_lo[11583:11568]},
     {storeUnit_maskInput_lo[11567:11552]},
     {storeUnit_maskInput_lo[11551:11536]},
     {storeUnit_maskInput_lo[11535:11520]},
     {storeUnit_maskInput_lo[11519:11504]},
     {storeUnit_maskInput_lo[11503:11488]},
     {storeUnit_maskInput_lo[11487:11472]},
     {storeUnit_maskInput_lo[11471:11456]},
     {storeUnit_maskInput_lo[11455:11440]},
     {storeUnit_maskInput_lo[11439:11424]},
     {storeUnit_maskInput_lo[11423:11408]},
     {storeUnit_maskInput_lo[11407:11392]},
     {storeUnit_maskInput_lo[11391:11376]},
     {storeUnit_maskInput_lo[11375:11360]},
     {storeUnit_maskInput_lo[11359:11344]},
     {storeUnit_maskInput_lo[11343:11328]},
     {storeUnit_maskInput_lo[11327:11312]},
     {storeUnit_maskInput_lo[11311:11296]},
     {storeUnit_maskInput_lo[11295:11280]},
     {storeUnit_maskInput_lo[11279:11264]},
     {storeUnit_maskInput_lo[11263:11248]},
     {storeUnit_maskInput_lo[11247:11232]},
     {storeUnit_maskInput_lo[11231:11216]},
     {storeUnit_maskInput_lo[11215:11200]},
     {storeUnit_maskInput_lo[11199:11184]},
     {storeUnit_maskInput_lo[11183:11168]},
     {storeUnit_maskInput_lo[11167:11152]},
     {storeUnit_maskInput_lo[11151:11136]},
     {storeUnit_maskInput_lo[11135:11120]},
     {storeUnit_maskInput_lo[11119:11104]},
     {storeUnit_maskInput_lo[11103:11088]},
     {storeUnit_maskInput_lo[11087:11072]},
     {storeUnit_maskInput_lo[11071:11056]},
     {storeUnit_maskInput_lo[11055:11040]},
     {storeUnit_maskInput_lo[11039:11024]},
     {storeUnit_maskInput_lo[11023:11008]},
     {storeUnit_maskInput_lo[11007:10992]},
     {storeUnit_maskInput_lo[10991:10976]},
     {storeUnit_maskInput_lo[10975:10960]},
     {storeUnit_maskInput_lo[10959:10944]},
     {storeUnit_maskInput_lo[10943:10928]},
     {storeUnit_maskInput_lo[10927:10912]},
     {storeUnit_maskInput_lo[10911:10896]},
     {storeUnit_maskInput_lo[10895:10880]},
     {storeUnit_maskInput_lo[10879:10864]},
     {storeUnit_maskInput_lo[10863:10848]},
     {storeUnit_maskInput_lo[10847:10832]},
     {storeUnit_maskInput_lo[10831:10816]},
     {storeUnit_maskInput_lo[10815:10800]},
     {storeUnit_maskInput_lo[10799:10784]},
     {storeUnit_maskInput_lo[10783:10768]},
     {storeUnit_maskInput_lo[10767:10752]},
     {storeUnit_maskInput_lo[10751:10736]},
     {storeUnit_maskInput_lo[10735:10720]},
     {storeUnit_maskInput_lo[10719:10704]},
     {storeUnit_maskInput_lo[10703:10688]},
     {storeUnit_maskInput_lo[10687:10672]},
     {storeUnit_maskInput_lo[10671:10656]},
     {storeUnit_maskInput_lo[10655:10640]},
     {storeUnit_maskInput_lo[10639:10624]},
     {storeUnit_maskInput_lo[10623:10608]},
     {storeUnit_maskInput_lo[10607:10592]},
     {storeUnit_maskInput_lo[10591:10576]},
     {storeUnit_maskInput_lo[10575:10560]},
     {storeUnit_maskInput_lo[10559:10544]},
     {storeUnit_maskInput_lo[10543:10528]},
     {storeUnit_maskInput_lo[10527:10512]},
     {storeUnit_maskInput_lo[10511:10496]},
     {storeUnit_maskInput_lo[10495:10480]},
     {storeUnit_maskInput_lo[10479:10464]},
     {storeUnit_maskInput_lo[10463:10448]},
     {storeUnit_maskInput_lo[10447:10432]},
     {storeUnit_maskInput_lo[10431:10416]},
     {storeUnit_maskInput_lo[10415:10400]},
     {storeUnit_maskInput_lo[10399:10384]},
     {storeUnit_maskInput_lo[10383:10368]},
     {storeUnit_maskInput_lo[10367:10352]},
     {storeUnit_maskInput_lo[10351:10336]},
     {storeUnit_maskInput_lo[10335:10320]},
     {storeUnit_maskInput_lo[10319:10304]},
     {storeUnit_maskInput_lo[10303:10288]},
     {storeUnit_maskInput_lo[10287:10272]},
     {storeUnit_maskInput_lo[10271:10256]},
     {storeUnit_maskInput_lo[10255:10240]},
     {storeUnit_maskInput_lo[10239:10224]},
     {storeUnit_maskInput_lo[10223:10208]},
     {storeUnit_maskInput_lo[10207:10192]},
     {storeUnit_maskInput_lo[10191:10176]},
     {storeUnit_maskInput_lo[10175:10160]},
     {storeUnit_maskInput_lo[10159:10144]},
     {storeUnit_maskInput_lo[10143:10128]},
     {storeUnit_maskInput_lo[10127:10112]},
     {storeUnit_maskInput_lo[10111:10096]},
     {storeUnit_maskInput_lo[10095:10080]},
     {storeUnit_maskInput_lo[10079:10064]},
     {storeUnit_maskInput_lo[10063:10048]},
     {storeUnit_maskInput_lo[10047:10032]},
     {storeUnit_maskInput_lo[10031:10016]},
     {storeUnit_maskInput_lo[10015:10000]},
     {storeUnit_maskInput_lo[9999:9984]},
     {storeUnit_maskInput_lo[9983:9968]},
     {storeUnit_maskInput_lo[9967:9952]},
     {storeUnit_maskInput_lo[9951:9936]},
     {storeUnit_maskInput_lo[9935:9920]},
     {storeUnit_maskInput_lo[9919:9904]},
     {storeUnit_maskInput_lo[9903:9888]},
     {storeUnit_maskInput_lo[9887:9872]},
     {storeUnit_maskInput_lo[9871:9856]},
     {storeUnit_maskInput_lo[9855:9840]},
     {storeUnit_maskInput_lo[9839:9824]},
     {storeUnit_maskInput_lo[9823:9808]},
     {storeUnit_maskInput_lo[9807:9792]},
     {storeUnit_maskInput_lo[9791:9776]},
     {storeUnit_maskInput_lo[9775:9760]},
     {storeUnit_maskInput_lo[9759:9744]},
     {storeUnit_maskInput_lo[9743:9728]},
     {storeUnit_maskInput_lo[9727:9712]},
     {storeUnit_maskInput_lo[9711:9696]},
     {storeUnit_maskInput_lo[9695:9680]},
     {storeUnit_maskInput_lo[9679:9664]},
     {storeUnit_maskInput_lo[9663:9648]},
     {storeUnit_maskInput_lo[9647:9632]},
     {storeUnit_maskInput_lo[9631:9616]},
     {storeUnit_maskInput_lo[9615:9600]},
     {storeUnit_maskInput_lo[9599:9584]},
     {storeUnit_maskInput_lo[9583:9568]},
     {storeUnit_maskInput_lo[9567:9552]},
     {storeUnit_maskInput_lo[9551:9536]},
     {storeUnit_maskInput_lo[9535:9520]},
     {storeUnit_maskInput_lo[9519:9504]},
     {storeUnit_maskInput_lo[9503:9488]},
     {storeUnit_maskInput_lo[9487:9472]},
     {storeUnit_maskInput_lo[9471:9456]},
     {storeUnit_maskInput_lo[9455:9440]},
     {storeUnit_maskInput_lo[9439:9424]},
     {storeUnit_maskInput_lo[9423:9408]},
     {storeUnit_maskInput_lo[9407:9392]},
     {storeUnit_maskInput_lo[9391:9376]},
     {storeUnit_maskInput_lo[9375:9360]},
     {storeUnit_maskInput_lo[9359:9344]},
     {storeUnit_maskInput_lo[9343:9328]},
     {storeUnit_maskInput_lo[9327:9312]},
     {storeUnit_maskInput_lo[9311:9296]},
     {storeUnit_maskInput_lo[9295:9280]},
     {storeUnit_maskInput_lo[9279:9264]},
     {storeUnit_maskInput_lo[9263:9248]},
     {storeUnit_maskInput_lo[9247:9232]},
     {storeUnit_maskInput_lo[9231:9216]},
     {storeUnit_maskInput_lo[9215:9200]},
     {storeUnit_maskInput_lo[9199:9184]},
     {storeUnit_maskInput_lo[9183:9168]},
     {storeUnit_maskInput_lo[9167:9152]},
     {storeUnit_maskInput_lo[9151:9136]},
     {storeUnit_maskInput_lo[9135:9120]},
     {storeUnit_maskInput_lo[9119:9104]},
     {storeUnit_maskInput_lo[9103:9088]},
     {storeUnit_maskInput_lo[9087:9072]},
     {storeUnit_maskInput_lo[9071:9056]},
     {storeUnit_maskInput_lo[9055:9040]},
     {storeUnit_maskInput_lo[9039:9024]},
     {storeUnit_maskInput_lo[9023:9008]},
     {storeUnit_maskInput_lo[9007:8992]},
     {storeUnit_maskInput_lo[8991:8976]},
     {storeUnit_maskInput_lo[8975:8960]},
     {storeUnit_maskInput_lo[8959:8944]},
     {storeUnit_maskInput_lo[8943:8928]},
     {storeUnit_maskInput_lo[8927:8912]},
     {storeUnit_maskInput_lo[8911:8896]},
     {storeUnit_maskInput_lo[8895:8880]},
     {storeUnit_maskInput_lo[8879:8864]},
     {storeUnit_maskInput_lo[8863:8848]},
     {storeUnit_maskInput_lo[8847:8832]},
     {storeUnit_maskInput_lo[8831:8816]},
     {storeUnit_maskInput_lo[8815:8800]},
     {storeUnit_maskInput_lo[8799:8784]},
     {storeUnit_maskInput_lo[8783:8768]},
     {storeUnit_maskInput_lo[8767:8752]},
     {storeUnit_maskInput_lo[8751:8736]},
     {storeUnit_maskInput_lo[8735:8720]},
     {storeUnit_maskInput_lo[8719:8704]},
     {storeUnit_maskInput_lo[8703:8688]},
     {storeUnit_maskInput_lo[8687:8672]},
     {storeUnit_maskInput_lo[8671:8656]},
     {storeUnit_maskInput_lo[8655:8640]},
     {storeUnit_maskInput_lo[8639:8624]},
     {storeUnit_maskInput_lo[8623:8608]},
     {storeUnit_maskInput_lo[8607:8592]},
     {storeUnit_maskInput_lo[8591:8576]},
     {storeUnit_maskInput_lo[8575:8560]},
     {storeUnit_maskInput_lo[8559:8544]},
     {storeUnit_maskInput_lo[8543:8528]},
     {storeUnit_maskInput_lo[8527:8512]},
     {storeUnit_maskInput_lo[8511:8496]},
     {storeUnit_maskInput_lo[8495:8480]},
     {storeUnit_maskInput_lo[8479:8464]},
     {storeUnit_maskInput_lo[8463:8448]},
     {storeUnit_maskInput_lo[8447:8432]},
     {storeUnit_maskInput_lo[8431:8416]},
     {storeUnit_maskInput_lo[8415:8400]},
     {storeUnit_maskInput_lo[8399:8384]},
     {storeUnit_maskInput_lo[8383:8368]},
     {storeUnit_maskInput_lo[8367:8352]},
     {storeUnit_maskInput_lo[8351:8336]},
     {storeUnit_maskInput_lo[8335:8320]},
     {storeUnit_maskInput_lo[8319:8304]},
     {storeUnit_maskInput_lo[8303:8288]},
     {storeUnit_maskInput_lo[8287:8272]},
     {storeUnit_maskInput_lo[8271:8256]},
     {storeUnit_maskInput_lo[8255:8240]},
     {storeUnit_maskInput_lo[8239:8224]},
     {storeUnit_maskInput_lo[8223:8208]},
     {storeUnit_maskInput_lo[8207:8192]},
     {storeUnit_maskInput_lo[8191:8176]},
     {storeUnit_maskInput_lo[8175:8160]},
     {storeUnit_maskInput_lo[8159:8144]},
     {storeUnit_maskInput_lo[8143:8128]},
     {storeUnit_maskInput_lo[8127:8112]},
     {storeUnit_maskInput_lo[8111:8096]},
     {storeUnit_maskInput_lo[8095:8080]},
     {storeUnit_maskInput_lo[8079:8064]},
     {storeUnit_maskInput_lo[8063:8048]},
     {storeUnit_maskInput_lo[8047:8032]},
     {storeUnit_maskInput_lo[8031:8016]},
     {storeUnit_maskInput_lo[8015:8000]},
     {storeUnit_maskInput_lo[7999:7984]},
     {storeUnit_maskInput_lo[7983:7968]},
     {storeUnit_maskInput_lo[7967:7952]},
     {storeUnit_maskInput_lo[7951:7936]},
     {storeUnit_maskInput_lo[7935:7920]},
     {storeUnit_maskInput_lo[7919:7904]},
     {storeUnit_maskInput_lo[7903:7888]},
     {storeUnit_maskInput_lo[7887:7872]},
     {storeUnit_maskInput_lo[7871:7856]},
     {storeUnit_maskInput_lo[7855:7840]},
     {storeUnit_maskInput_lo[7839:7824]},
     {storeUnit_maskInput_lo[7823:7808]},
     {storeUnit_maskInput_lo[7807:7792]},
     {storeUnit_maskInput_lo[7791:7776]},
     {storeUnit_maskInput_lo[7775:7760]},
     {storeUnit_maskInput_lo[7759:7744]},
     {storeUnit_maskInput_lo[7743:7728]},
     {storeUnit_maskInput_lo[7727:7712]},
     {storeUnit_maskInput_lo[7711:7696]},
     {storeUnit_maskInput_lo[7695:7680]},
     {storeUnit_maskInput_lo[7679:7664]},
     {storeUnit_maskInput_lo[7663:7648]},
     {storeUnit_maskInput_lo[7647:7632]},
     {storeUnit_maskInput_lo[7631:7616]},
     {storeUnit_maskInput_lo[7615:7600]},
     {storeUnit_maskInput_lo[7599:7584]},
     {storeUnit_maskInput_lo[7583:7568]},
     {storeUnit_maskInput_lo[7567:7552]},
     {storeUnit_maskInput_lo[7551:7536]},
     {storeUnit_maskInput_lo[7535:7520]},
     {storeUnit_maskInput_lo[7519:7504]},
     {storeUnit_maskInput_lo[7503:7488]},
     {storeUnit_maskInput_lo[7487:7472]},
     {storeUnit_maskInput_lo[7471:7456]},
     {storeUnit_maskInput_lo[7455:7440]},
     {storeUnit_maskInput_lo[7439:7424]},
     {storeUnit_maskInput_lo[7423:7408]},
     {storeUnit_maskInput_lo[7407:7392]},
     {storeUnit_maskInput_lo[7391:7376]},
     {storeUnit_maskInput_lo[7375:7360]},
     {storeUnit_maskInput_lo[7359:7344]},
     {storeUnit_maskInput_lo[7343:7328]},
     {storeUnit_maskInput_lo[7327:7312]},
     {storeUnit_maskInput_lo[7311:7296]},
     {storeUnit_maskInput_lo[7295:7280]},
     {storeUnit_maskInput_lo[7279:7264]},
     {storeUnit_maskInput_lo[7263:7248]},
     {storeUnit_maskInput_lo[7247:7232]},
     {storeUnit_maskInput_lo[7231:7216]},
     {storeUnit_maskInput_lo[7215:7200]},
     {storeUnit_maskInput_lo[7199:7184]},
     {storeUnit_maskInput_lo[7183:7168]},
     {storeUnit_maskInput_lo[7167:7152]},
     {storeUnit_maskInput_lo[7151:7136]},
     {storeUnit_maskInput_lo[7135:7120]},
     {storeUnit_maskInput_lo[7119:7104]},
     {storeUnit_maskInput_lo[7103:7088]},
     {storeUnit_maskInput_lo[7087:7072]},
     {storeUnit_maskInput_lo[7071:7056]},
     {storeUnit_maskInput_lo[7055:7040]},
     {storeUnit_maskInput_lo[7039:7024]},
     {storeUnit_maskInput_lo[7023:7008]},
     {storeUnit_maskInput_lo[7007:6992]},
     {storeUnit_maskInput_lo[6991:6976]},
     {storeUnit_maskInput_lo[6975:6960]},
     {storeUnit_maskInput_lo[6959:6944]},
     {storeUnit_maskInput_lo[6943:6928]},
     {storeUnit_maskInput_lo[6927:6912]},
     {storeUnit_maskInput_lo[6911:6896]},
     {storeUnit_maskInput_lo[6895:6880]},
     {storeUnit_maskInput_lo[6879:6864]},
     {storeUnit_maskInput_lo[6863:6848]},
     {storeUnit_maskInput_lo[6847:6832]},
     {storeUnit_maskInput_lo[6831:6816]},
     {storeUnit_maskInput_lo[6815:6800]},
     {storeUnit_maskInput_lo[6799:6784]},
     {storeUnit_maskInput_lo[6783:6768]},
     {storeUnit_maskInput_lo[6767:6752]},
     {storeUnit_maskInput_lo[6751:6736]},
     {storeUnit_maskInput_lo[6735:6720]},
     {storeUnit_maskInput_lo[6719:6704]},
     {storeUnit_maskInput_lo[6703:6688]},
     {storeUnit_maskInput_lo[6687:6672]},
     {storeUnit_maskInput_lo[6671:6656]},
     {storeUnit_maskInput_lo[6655:6640]},
     {storeUnit_maskInput_lo[6639:6624]},
     {storeUnit_maskInput_lo[6623:6608]},
     {storeUnit_maskInput_lo[6607:6592]},
     {storeUnit_maskInput_lo[6591:6576]},
     {storeUnit_maskInput_lo[6575:6560]},
     {storeUnit_maskInput_lo[6559:6544]},
     {storeUnit_maskInput_lo[6543:6528]},
     {storeUnit_maskInput_lo[6527:6512]},
     {storeUnit_maskInput_lo[6511:6496]},
     {storeUnit_maskInput_lo[6495:6480]},
     {storeUnit_maskInput_lo[6479:6464]},
     {storeUnit_maskInput_lo[6463:6448]},
     {storeUnit_maskInput_lo[6447:6432]},
     {storeUnit_maskInput_lo[6431:6416]},
     {storeUnit_maskInput_lo[6415:6400]},
     {storeUnit_maskInput_lo[6399:6384]},
     {storeUnit_maskInput_lo[6383:6368]},
     {storeUnit_maskInput_lo[6367:6352]},
     {storeUnit_maskInput_lo[6351:6336]},
     {storeUnit_maskInput_lo[6335:6320]},
     {storeUnit_maskInput_lo[6319:6304]},
     {storeUnit_maskInput_lo[6303:6288]},
     {storeUnit_maskInput_lo[6287:6272]},
     {storeUnit_maskInput_lo[6271:6256]},
     {storeUnit_maskInput_lo[6255:6240]},
     {storeUnit_maskInput_lo[6239:6224]},
     {storeUnit_maskInput_lo[6223:6208]},
     {storeUnit_maskInput_lo[6207:6192]},
     {storeUnit_maskInput_lo[6191:6176]},
     {storeUnit_maskInput_lo[6175:6160]},
     {storeUnit_maskInput_lo[6159:6144]},
     {storeUnit_maskInput_lo[6143:6128]},
     {storeUnit_maskInput_lo[6127:6112]},
     {storeUnit_maskInput_lo[6111:6096]},
     {storeUnit_maskInput_lo[6095:6080]},
     {storeUnit_maskInput_lo[6079:6064]},
     {storeUnit_maskInput_lo[6063:6048]},
     {storeUnit_maskInput_lo[6047:6032]},
     {storeUnit_maskInput_lo[6031:6016]},
     {storeUnit_maskInput_lo[6015:6000]},
     {storeUnit_maskInput_lo[5999:5984]},
     {storeUnit_maskInput_lo[5983:5968]},
     {storeUnit_maskInput_lo[5967:5952]},
     {storeUnit_maskInput_lo[5951:5936]},
     {storeUnit_maskInput_lo[5935:5920]},
     {storeUnit_maskInput_lo[5919:5904]},
     {storeUnit_maskInput_lo[5903:5888]},
     {storeUnit_maskInput_lo[5887:5872]},
     {storeUnit_maskInput_lo[5871:5856]},
     {storeUnit_maskInput_lo[5855:5840]},
     {storeUnit_maskInput_lo[5839:5824]},
     {storeUnit_maskInput_lo[5823:5808]},
     {storeUnit_maskInput_lo[5807:5792]},
     {storeUnit_maskInput_lo[5791:5776]},
     {storeUnit_maskInput_lo[5775:5760]},
     {storeUnit_maskInput_lo[5759:5744]},
     {storeUnit_maskInput_lo[5743:5728]},
     {storeUnit_maskInput_lo[5727:5712]},
     {storeUnit_maskInput_lo[5711:5696]},
     {storeUnit_maskInput_lo[5695:5680]},
     {storeUnit_maskInput_lo[5679:5664]},
     {storeUnit_maskInput_lo[5663:5648]},
     {storeUnit_maskInput_lo[5647:5632]},
     {storeUnit_maskInput_lo[5631:5616]},
     {storeUnit_maskInput_lo[5615:5600]},
     {storeUnit_maskInput_lo[5599:5584]},
     {storeUnit_maskInput_lo[5583:5568]},
     {storeUnit_maskInput_lo[5567:5552]},
     {storeUnit_maskInput_lo[5551:5536]},
     {storeUnit_maskInput_lo[5535:5520]},
     {storeUnit_maskInput_lo[5519:5504]},
     {storeUnit_maskInput_lo[5503:5488]},
     {storeUnit_maskInput_lo[5487:5472]},
     {storeUnit_maskInput_lo[5471:5456]},
     {storeUnit_maskInput_lo[5455:5440]},
     {storeUnit_maskInput_lo[5439:5424]},
     {storeUnit_maskInput_lo[5423:5408]},
     {storeUnit_maskInput_lo[5407:5392]},
     {storeUnit_maskInput_lo[5391:5376]},
     {storeUnit_maskInput_lo[5375:5360]},
     {storeUnit_maskInput_lo[5359:5344]},
     {storeUnit_maskInput_lo[5343:5328]},
     {storeUnit_maskInput_lo[5327:5312]},
     {storeUnit_maskInput_lo[5311:5296]},
     {storeUnit_maskInput_lo[5295:5280]},
     {storeUnit_maskInput_lo[5279:5264]},
     {storeUnit_maskInput_lo[5263:5248]},
     {storeUnit_maskInput_lo[5247:5232]},
     {storeUnit_maskInput_lo[5231:5216]},
     {storeUnit_maskInput_lo[5215:5200]},
     {storeUnit_maskInput_lo[5199:5184]},
     {storeUnit_maskInput_lo[5183:5168]},
     {storeUnit_maskInput_lo[5167:5152]},
     {storeUnit_maskInput_lo[5151:5136]},
     {storeUnit_maskInput_lo[5135:5120]},
     {storeUnit_maskInput_lo[5119:5104]},
     {storeUnit_maskInput_lo[5103:5088]},
     {storeUnit_maskInput_lo[5087:5072]},
     {storeUnit_maskInput_lo[5071:5056]},
     {storeUnit_maskInput_lo[5055:5040]},
     {storeUnit_maskInput_lo[5039:5024]},
     {storeUnit_maskInput_lo[5023:5008]},
     {storeUnit_maskInput_lo[5007:4992]},
     {storeUnit_maskInput_lo[4991:4976]},
     {storeUnit_maskInput_lo[4975:4960]},
     {storeUnit_maskInput_lo[4959:4944]},
     {storeUnit_maskInput_lo[4943:4928]},
     {storeUnit_maskInput_lo[4927:4912]},
     {storeUnit_maskInput_lo[4911:4896]},
     {storeUnit_maskInput_lo[4895:4880]},
     {storeUnit_maskInput_lo[4879:4864]},
     {storeUnit_maskInput_lo[4863:4848]},
     {storeUnit_maskInput_lo[4847:4832]},
     {storeUnit_maskInput_lo[4831:4816]},
     {storeUnit_maskInput_lo[4815:4800]},
     {storeUnit_maskInput_lo[4799:4784]},
     {storeUnit_maskInput_lo[4783:4768]},
     {storeUnit_maskInput_lo[4767:4752]},
     {storeUnit_maskInput_lo[4751:4736]},
     {storeUnit_maskInput_lo[4735:4720]},
     {storeUnit_maskInput_lo[4719:4704]},
     {storeUnit_maskInput_lo[4703:4688]},
     {storeUnit_maskInput_lo[4687:4672]},
     {storeUnit_maskInput_lo[4671:4656]},
     {storeUnit_maskInput_lo[4655:4640]},
     {storeUnit_maskInput_lo[4639:4624]},
     {storeUnit_maskInput_lo[4623:4608]},
     {storeUnit_maskInput_lo[4607:4592]},
     {storeUnit_maskInput_lo[4591:4576]},
     {storeUnit_maskInput_lo[4575:4560]},
     {storeUnit_maskInput_lo[4559:4544]},
     {storeUnit_maskInput_lo[4543:4528]},
     {storeUnit_maskInput_lo[4527:4512]},
     {storeUnit_maskInput_lo[4511:4496]},
     {storeUnit_maskInput_lo[4495:4480]},
     {storeUnit_maskInput_lo[4479:4464]},
     {storeUnit_maskInput_lo[4463:4448]},
     {storeUnit_maskInput_lo[4447:4432]},
     {storeUnit_maskInput_lo[4431:4416]},
     {storeUnit_maskInput_lo[4415:4400]},
     {storeUnit_maskInput_lo[4399:4384]},
     {storeUnit_maskInput_lo[4383:4368]},
     {storeUnit_maskInput_lo[4367:4352]},
     {storeUnit_maskInput_lo[4351:4336]},
     {storeUnit_maskInput_lo[4335:4320]},
     {storeUnit_maskInput_lo[4319:4304]},
     {storeUnit_maskInput_lo[4303:4288]},
     {storeUnit_maskInput_lo[4287:4272]},
     {storeUnit_maskInput_lo[4271:4256]},
     {storeUnit_maskInput_lo[4255:4240]},
     {storeUnit_maskInput_lo[4239:4224]},
     {storeUnit_maskInput_lo[4223:4208]},
     {storeUnit_maskInput_lo[4207:4192]},
     {storeUnit_maskInput_lo[4191:4176]},
     {storeUnit_maskInput_lo[4175:4160]},
     {storeUnit_maskInput_lo[4159:4144]},
     {storeUnit_maskInput_lo[4143:4128]},
     {storeUnit_maskInput_lo[4127:4112]},
     {storeUnit_maskInput_lo[4111:4096]},
     {storeUnit_maskInput_lo[4095:4080]},
     {storeUnit_maskInput_lo[4079:4064]},
     {storeUnit_maskInput_lo[4063:4048]},
     {storeUnit_maskInput_lo[4047:4032]},
     {storeUnit_maskInput_lo[4031:4016]},
     {storeUnit_maskInput_lo[4015:4000]},
     {storeUnit_maskInput_lo[3999:3984]},
     {storeUnit_maskInput_lo[3983:3968]},
     {storeUnit_maskInput_lo[3967:3952]},
     {storeUnit_maskInput_lo[3951:3936]},
     {storeUnit_maskInput_lo[3935:3920]},
     {storeUnit_maskInput_lo[3919:3904]},
     {storeUnit_maskInput_lo[3903:3888]},
     {storeUnit_maskInput_lo[3887:3872]},
     {storeUnit_maskInput_lo[3871:3856]},
     {storeUnit_maskInput_lo[3855:3840]},
     {storeUnit_maskInput_lo[3839:3824]},
     {storeUnit_maskInput_lo[3823:3808]},
     {storeUnit_maskInput_lo[3807:3792]},
     {storeUnit_maskInput_lo[3791:3776]},
     {storeUnit_maskInput_lo[3775:3760]},
     {storeUnit_maskInput_lo[3759:3744]},
     {storeUnit_maskInput_lo[3743:3728]},
     {storeUnit_maskInput_lo[3727:3712]},
     {storeUnit_maskInput_lo[3711:3696]},
     {storeUnit_maskInput_lo[3695:3680]},
     {storeUnit_maskInput_lo[3679:3664]},
     {storeUnit_maskInput_lo[3663:3648]},
     {storeUnit_maskInput_lo[3647:3632]},
     {storeUnit_maskInput_lo[3631:3616]},
     {storeUnit_maskInput_lo[3615:3600]},
     {storeUnit_maskInput_lo[3599:3584]},
     {storeUnit_maskInput_lo[3583:3568]},
     {storeUnit_maskInput_lo[3567:3552]},
     {storeUnit_maskInput_lo[3551:3536]},
     {storeUnit_maskInput_lo[3535:3520]},
     {storeUnit_maskInput_lo[3519:3504]},
     {storeUnit_maskInput_lo[3503:3488]},
     {storeUnit_maskInput_lo[3487:3472]},
     {storeUnit_maskInput_lo[3471:3456]},
     {storeUnit_maskInput_lo[3455:3440]},
     {storeUnit_maskInput_lo[3439:3424]},
     {storeUnit_maskInput_lo[3423:3408]},
     {storeUnit_maskInput_lo[3407:3392]},
     {storeUnit_maskInput_lo[3391:3376]},
     {storeUnit_maskInput_lo[3375:3360]},
     {storeUnit_maskInput_lo[3359:3344]},
     {storeUnit_maskInput_lo[3343:3328]},
     {storeUnit_maskInput_lo[3327:3312]},
     {storeUnit_maskInput_lo[3311:3296]},
     {storeUnit_maskInput_lo[3295:3280]},
     {storeUnit_maskInput_lo[3279:3264]},
     {storeUnit_maskInput_lo[3263:3248]},
     {storeUnit_maskInput_lo[3247:3232]},
     {storeUnit_maskInput_lo[3231:3216]},
     {storeUnit_maskInput_lo[3215:3200]},
     {storeUnit_maskInput_lo[3199:3184]},
     {storeUnit_maskInput_lo[3183:3168]},
     {storeUnit_maskInput_lo[3167:3152]},
     {storeUnit_maskInput_lo[3151:3136]},
     {storeUnit_maskInput_lo[3135:3120]},
     {storeUnit_maskInput_lo[3119:3104]},
     {storeUnit_maskInput_lo[3103:3088]},
     {storeUnit_maskInput_lo[3087:3072]},
     {storeUnit_maskInput_lo[3071:3056]},
     {storeUnit_maskInput_lo[3055:3040]},
     {storeUnit_maskInput_lo[3039:3024]},
     {storeUnit_maskInput_lo[3023:3008]},
     {storeUnit_maskInput_lo[3007:2992]},
     {storeUnit_maskInput_lo[2991:2976]},
     {storeUnit_maskInput_lo[2975:2960]},
     {storeUnit_maskInput_lo[2959:2944]},
     {storeUnit_maskInput_lo[2943:2928]},
     {storeUnit_maskInput_lo[2927:2912]},
     {storeUnit_maskInput_lo[2911:2896]},
     {storeUnit_maskInput_lo[2895:2880]},
     {storeUnit_maskInput_lo[2879:2864]},
     {storeUnit_maskInput_lo[2863:2848]},
     {storeUnit_maskInput_lo[2847:2832]},
     {storeUnit_maskInput_lo[2831:2816]},
     {storeUnit_maskInput_lo[2815:2800]},
     {storeUnit_maskInput_lo[2799:2784]},
     {storeUnit_maskInput_lo[2783:2768]},
     {storeUnit_maskInput_lo[2767:2752]},
     {storeUnit_maskInput_lo[2751:2736]},
     {storeUnit_maskInput_lo[2735:2720]},
     {storeUnit_maskInput_lo[2719:2704]},
     {storeUnit_maskInput_lo[2703:2688]},
     {storeUnit_maskInput_lo[2687:2672]},
     {storeUnit_maskInput_lo[2671:2656]},
     {storeUnit_maskInput_lo[2655:2640]},
     {storeUnit_maskInput_lo[2639:2624]},
     {storeUnit_maskInput_lo[2623:2608]},
     {storeUnit_maskInput_lo[2607:2592]},
     {storeUnit_maskInput_lo[2591:2576]},
     {storeUnit_maskInput_lo[2575:2560]},
     {storeUnit_maskInput_lo[2559:2544]},
     {storeUnit_maskInput_lo[2543:2528]},
     {storeUnit_maskInput_lo[2527:2512]},
     {storeUnit_maskInput_lo[2511:2496]},
     {storeUnit_maskInput_lo[2495:2480]},
     {storeUnit_maskInput_lo[2479:2464]},
     {storeUnit_maskInput_lo[2463:2448]},
     {storeUnit_maskInput_lo[2447:2432]},
     {storeUnit_maskInput_lo[2431:2416]},
     {storeUnit_maskInput_lo[2415:2400]},
     {storeUnit_maskInput_lo[2399:2384]},
     {storeUnit_maskInput_lo[2383:2368]},
     {storeUnit_maskInput_lo[2367:2352]},
     {storeUnit_maskInput_lo[2351:2336]},
     {storeUnit_maskInput_lo[2335:2320]},
     {storeUnit_maskInput_lo[2319:2304]},
     {storeUnit_maskInput_lo[2303:2288]},
     {storeUnit_maskInput_lo[2287:2272]},
     {storeUnit_maskInput_lo[2271:2256]},
     {storeUnit_maskInput_lo[2255:2240]},
     {storeUnit_maskInput_lo[2239:2224]},
     {storeUnit_maskInput_lo[2223:2208]},
     {storeUnit_maskInput_lo[2207:2192]},
     {storeUnit_maskInput_lo[2191:2176]},
     {storeUnit_maskInput_lo[2175:2160]},
     {storeUnit_maskInput_lo[2159:2144]},
     {storeUnit_maskInput_lo[2143:2128]},
     {storeUnit_maskInput_lo[2127:2112]},
     {storeUnit_maskInput_lo[2111:2096]},
     {storeUnit_maskInput_lo[2095:2080]},
     {storeUnit_maskInput_lo[2079:2064]},
     {storeUnit_maskInput_lo[2063:2048]},
     {storeUnit_maskInput_lo[2047:2032]},
     {storeUnit_maskInput_lo[2031:2016]},
     {storeUnit_maskInput_lo[2015:2000]},
     {storeUnit_maskInput_lo[1999:1984]},
     {storeUnit_maskInput_lo[1983:1968]},
     {storeUnit_maskInput_lo[1967:1952]},
     {storeUnit_maskInput_lo[1951:1936]},
     {storeUnit_maskInput_lo[1935:1920]},
     {storeUnit_maskInput_lo[1919:1904]},
     {storeUnit_maskInput_lo[1903:1888]},
     {storeUnit_maskInput_lo[1887:1872]},
     {storeUnit_maskInput_lo[1871:1856]},
     {storeUnit_maskInput_lo[1855:1840]},
     {storeUnit_maskInput_lo[1839:1824]},
     {storeUnit_maskInput_lo[1823:1808]},
     {storeUnit_maskInput_lo[1807:1792]},
     {storeUnit_maskInput_lo[1791:1776]},
     {storeUnit_maskInput_lo[1775:1760]},
     {storeUnit_maskInput_lo[1759:1744]},
     {storeUnit_maskInput_lo[1743:1728]},
     {storeUnit_maskInput_lo[1727:1712]},
     {storeUnit_maskInput_lo[1711:1696]},
     {storeUnit_maskInput_lo[1695:1680]},
     {storeUnit_maskInput_lo[1679:1664]},
     {storeUnit_maskInput_lo[1663:1648]},
     {storeUnit_maskInput_lo[1647:1632]},
     {storeUnit_maskInput_lo[1631:1616]},
     {storeUnit_maskInput_lo[1615:1600]},
     {storeUnit_maskInput_lo[1599:1584]},
     {storeUnit_maskInput_lo[1583:1568]},
     {storeUnit_maskInput_lo[1567:1552]},
     {storeUnit_maskInput_lo[1551:1536]},
     {storeUnit_maskInput_lo[1535:1520]},
     {storeUnit_maskInput_lo[1519:1504]},
     {storeUnit_maskInput_lo[1503:1488]},
     {storeUnit_maskInput_lo[1487:1472]},
     {storeUnit_maskInput_lo[1471:1456]},
     {storeUnit_maskInput_lo[1455:1440]},
     {storeUnit_maskInput_lo[1439:1424]},
     {storeUnit_maskInput_lo[1423:1408]},
     {storeUnit_maskInput_lo[1407:1392]},
     {storeUnit_maskInput_lo[1391:1376]},
     {storeUnit_maskInput_lo[1375:1360]},
     {storeUnit_maskInput_lo[1359:1344]},
     {storeUnit_maskInput_lo[1343:1328]},
     {storeUnit_maskInput_lo[1327:1312]},
     {storeUnit_maskInput_lo[1311:1296]},
     {storeUnit_maskInput_lo[1295:1280]},
     {storeUnit_maskInput_lo[1279:1264]},
     {storeUnit_maskInput_lo[1263:1248]},
     {storeUnit_maskInput_lo[1247:1232]},
     {storeUnit_maskInput_lo[1231:1216]},
     {storeUnit_maskInput_lo[1215:1200]},
     {storeUnit_maskInput_lo[1199:1184]},
     {storeUnit_maskInput_lo[1183:1168]},
     {storeUnit_maskInput_lo[1167:1152]},
     {storeUnit_maskInput_lo[1151:1136]},
     {storeUnit_maskInput_lo[1135:1120]},
     {storeUnit_maskInput_lo[1119:1104]},
     {storeUnit_maskInput_lo[1103:1088]},
     {storeUnit_maskInput_lo[1087:1072]},
     {storeUnit_maskInput_lo[1071:1056]},
     {storeUnit_maskInput_lo[1055:1040]},
     {storeUnit_maskInput_lo[1039:1024]},
     {storeUnit_maskInput_lo[1023:1008]},
     {storeUnit_maskInput_lo[1007:992]},
     {storeUnit_maskInput_lo[991:976]},
     {storeUnit_maskInput_lo[975:960]},
     {storeUnit_maskInput_lo[959:944]},
     {storeUnit_maskInput_lo[943:928]},
     {storeUnit_maskInput_lo[927:912]},
     {storeUnit_maskInput_lo[911:896]},
     {storeUnit_maskInput_lo[895:880]},
     {storeUnit_maskInput_lo[879:864]},
     {storeUnit_maskInput_lo[863:848]},
     {storeUnit_maskInput_lo[847:832]},
     {storeUnit_maskInput_lo[831:816]},
     {storeUnit_maskInput_lo[815:800]},
     {storeUnit_maskInput_lo[799:784]},
     {storeUnit_maskInput_lo[783:768]},
     {storeUnit_maskInput_lo[767:752]},
     {storeUnit_maskInput_lo[751:736]},
     {storeUnit_maskInput_lo[735:720]},
     {storeUnit_maskInput_lo[719:704]},
     {storeUnit_maskInput_lo[703:688]},
     {storeUnit_maskInput_lo[687:672]},
     {storeUnit_maskInput_lo[671:656]},
     {storeUnit_maskInput_lo[655:640]},
     {storeUnit_maskInput_lo[639:624]},
     {storeUnit_maskInput_lo[623:608]},
     {storeUnit_maskInput_lo[607:592]},
     {storeUnit_maskInput_lo[591:576]},
     {storeUnit_maskInput_lo[575:560]},
     {storeUnit_maskInput_lo[559:544]},
     {storeUnit_maskInput_lo[543:528]},
     {storeUnit_maskInput_lo[527:512]},
     {storeUnit_maskInput_lo[511:496]},
     {storeUnit_maskInput_lo[495:480]},
     {storeUnit_maskInput_lo[479:464]},
     {storeUnit_maskInput_lo[463:448]},
     {storeUnit_maskInput_lo[447:432]},
     {storeUnit_maskInput_lo[431:416]},
     {storeUnit_maskInput_lo[415:400]},
     {storeUnit_maskInput_lo[399:384]},
     {storeUnit_maskInput_lo[383:368]},
     {storeUnit_maskInput_lo[367:352]},
     {storeUnit_maskInput_lo[351:336]},
     {storeUnit_maskInput_lo[335:320]},
     {storeUnit_maskInput_lo[319:304]},
     {storeUnit_maskInput_lo[303:288]},
     {storeUnit_maskInput_lo[287:272]},
     {storeUnit_maskInput_lo[271:256]},
     {storeUnit_maskInput_lo[255:240]},
     {storeUnit_maskInput_lo[239:224]},
     {storeUnit_maskInput_lo[223:208]},
     {storeUnit_maskInput_lo[207:192]},
     {storeUnit_maskInput_lo[191:176]},
     {storeUnit_maskInput_lo[175:160]},
     {storeUnit_maskInput_lo[159:144]},
     {storeUnit_maskInput_lo[143:128]},
     {storeUnit_maskInput_lo[127:112]},
     {storeUnit_maskInput_lo[111:96]},
     {storeUnit_maskInput_lo[95:80]},
     {storeUnit_maskInput_lo[79:64]},
     {storeUnit_maskInput_lo[63:48]},
     {storeUnit_maskInput_lo[47:32]},
     {storeUnit_maskInput_lo[31:16]},
     {storeUnit_maskInput_lo[15:0]}};
  wire [11:0]         maskSelect_2 = _otherUnit_maskSelect_valid ? _otherUnit_maskSelect_bits : 12'h0;
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi = {otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo = {otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi = {otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi = {otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo = {otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi = {otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo = {otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo = {otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi = {otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi = {otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi = {otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_lo_lo_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi = {otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo = {otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo = {otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi = {otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi = {otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo = {otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo = {otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi = {otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo = {otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo = {otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi = {otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi = {otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi = {otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_lo_lo_lo_lo_hi = {otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo};
  wire [2047:0]       otherUnit_maskInput_lo_lo_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi = {otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo = {otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi = {otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi = {otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo = {otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo = {otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi = {otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo = {otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo = {otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi = {otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi = {otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi = {otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_lo_lo_lo_hi_lo = {otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi = {otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo = {otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo = {otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi = {otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi = {otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo = {otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo = {otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi = {otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo = {otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo = {otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi = {otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi = {otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi = {otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_lo_lo_lo_hi_hi = {otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo};
  wire [2047:0]       otherUnit_maskInput_lo_lo_lo_lo_hi = {otherUnit_maskInput_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_lo};
  wire [4095:0]       otherUnit_maskInput_lo_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi = {otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo = {otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi = {otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi = {otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo = {otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi = {otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo = {otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo = {otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi = {otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi = {otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi = {otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_lo_lo_hi_lo_lo = {otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi = {otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo = {otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo = {otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi = {otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi = {otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo = {otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo = {otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi = {otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo = {otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo = {otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi = {otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi = {otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi = {otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_lo_lo_hi_lo_hi = {otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo};
  wire [2047:0]       otherUnit_maskInput_lo_lo_lo_hi_lo = {otherUnit_maskInput_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi = {otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo = {otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi = {otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi = {otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo = {otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo = {otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi = {otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo = {otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo = {otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi = {otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi = {otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi = {otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_lo_lo_hi_hi_lo = {otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi = {otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo = {otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo = {otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi = {otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi = {otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo = {otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo = {otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi = {otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo = {otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo = {otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi = {otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi = {otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi = {otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_lo_lo_hi_hi_hi = {otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo};
  wire [2047:0]       otherUnit_maskInput_lo_lo_lo_hi_hi = {otherUnit_maskInput_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_lo};
  wire [4095:0]       otherUnit_maskInput_lo_lo_lo_hi = {otherUnit_maskInput_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_lo};
  wire [8191:0]       otherUnit_maskInput_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo = {otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi = {otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo = {otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo = {otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi = {otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi = {otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo = {otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo = {otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi = {otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo = {otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo = {otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi = {otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi = {otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi = {otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_lo_hi_lo_lo_lo = {otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo = {otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi = {otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo = {otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo = {otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi = {otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi = {otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo = {otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo = {otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi = {otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo = {otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo = {otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi = {otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi = {otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi = {otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_lo_hi_lo_lo_hi = {otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo};
  wire [2047:0]       otherUnit_maskInput_lo_lo_hi_lo_lo = {otherUnit_maskInput_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo = {otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi = {otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo = {otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo = {otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi = {otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi = {otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo = {otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo = {otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi = {otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo = {otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo = {otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi = {otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi = {otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi = {otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_lo_hi_lo_hi_lo = {otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo = {otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi = {otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo = {otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo = {otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi = {otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi = {otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo = {otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo = {otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi = {otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo = {otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo = {otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi = {otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi = {otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi = {otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_lo_hi_lo_hi_hi = {otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo};
  wire [2047:0]       otherUnit_maskInput_lo_lo_hi_lo_hi = {otherUnit_maskInput_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_lo};
  wire [4095:0]       otherUnit_maskInput_lo_lo_hi_lo = {otherUnit_maskInput_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo = {otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi = {otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo = {otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo = {otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi = {otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi = {otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo = {otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo = {otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi = {otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo = {otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo = {otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi = {otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi = {otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi = {otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_lo_hi_hi_lo_lo = {otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo = {otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi = {otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo = {otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo = {otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi = {otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi = {otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo = {otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo = {otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi = {otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo = {otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo = {otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi = {otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi = {otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi = {otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_lo_hi_hi_lo_hi = {otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo};
  wire [2047:0]       otherUnit_maskInput_lo_lo_hi_hi_lo = {otherUnit_maskInput_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo = {otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi = {otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo = {otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo = {otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi = {otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi = {otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo = {otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo = {otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi = {otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo = {otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo = {otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi = {otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi = {otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi = {otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_lo_hi_hi_hi_lo = {otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo = {otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi = {otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo = {otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo = {otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi = {otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi = {otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo = {otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo = {otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi = {otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo = {otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo = {otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi = {otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi = {otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi = {otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_lo_hi_hi_hi_hi = {otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo};
  wire [2047:0]       otherUnit_maskInput_lo_lo_hi_hi_hi = {otherUnit_maskInput_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_lo};
  wire [4095:0]       otherUnit_maskInput_lo_lo_hi_hi = {otherUnit_maskInput_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_lo};
  wire [8191:0]       otherUnit_maskInput_lo_lo_hi = {otherUnit_maskInput_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo};
  wire [16383:0]      otherUnit_maskInput_lo_lo = {otherUnit_maskInput_lo_lo_hi, otherUnit_maskInput_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo = {otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi = {otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo = {otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi = {otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi = {otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo = {otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo = {otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi = {otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo = {otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi = {otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi = {otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi = {otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_hi_lo_lo_lo_lo = {otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo = {otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi = {otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo = {otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi = {otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi = {otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo = {otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi = {otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo = {otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo = {otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi = {otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi = {otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi = {otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_hi_lo_lo_lo_hi = {otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo};
  wire [2047:0]       otherUnit_maskInput_lo_hi_lo_lo_lo = {otherUnit_maskInput_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo = {otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi = {otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo = {otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi = {otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi = {otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo = {otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo = {otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi = {otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo = {otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi = {otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi = {otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi = {otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_hi_lo_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo = {otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi = {otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo = {otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi = {otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi = {otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo = {otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo = {otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi = {otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo = {otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo = {otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi = {otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi = {otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi = {otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_hi_lo_lo_hi_hi = {otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo};
  wire [2047:0]       otherUnit_maskInput_lo_hi_lo_lo_hi = {otherUnit_maskInput_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_lo};
  wire [4095:0]       otherUnit_maskInput_lo_hi_lo_lo = {otherUnit_maskInput_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo = {otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi = {otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo = {otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi = {otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi = {otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo = {otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo = {otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi = {otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi = {otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi = {otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi = {otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_hi_lo_hi_lo_lo = {otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo = {otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi = {otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo = {otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi = {otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi = {otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo = {otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi = {otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi = {otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi = {otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi = {otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_hi_lo_hi_lo_hi = {otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo};
  wire [2047:0]       otherUnit_maskInput_lo_hi_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo = {otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi = {otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo = {otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi = {otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi = {otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo = {otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo = {otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi = {otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi = {otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi = {otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi = {otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_hi_lo_hi_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo = {otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi = {otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo = {otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi = {otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi = {otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo = {otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi = {otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi = {otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi = {otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi = {otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_hi_lo_hi_hi_hi = {otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo};
  wire [2047:0]       otherUnit_maskInput_lo_hi_lo_hi_hi = {otherUnit_maskInput_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_lo};
  wire [4095:0]       otherUnit_maskInput_lo_hi_lo_hi = {otherUnit_maskInput_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_lo};
  wire [8191:0]       otherUnit_maskInput_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo = {otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi = {otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo = {otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo = {otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi = {otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi = {otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo = {otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo = {otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi = {otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo = {otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo = {otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi = {otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi = {otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi = {otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_hi_hi_lo_lo_lo = {otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo = {otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi = {otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo = {otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo = {otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi = {otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi = {otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo = {otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo = {otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi = {otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo = {otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo = {otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi = {otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi = {otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi = {otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_hi_hi_lo_lo_hi = {otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo};
  wire [2047:0]       otherUnit_maskInput_lo_hi_hi_lo_lo = {otherUnit_maskInput_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo = {otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi = {otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo = {otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo = {otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi = {otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi = {otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo = {otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo = {otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi = {otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo = {otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo = {otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi = {otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi = {otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi = {otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_hi_hi_lo_hi_lo = {otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo = {otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi = {otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo = {otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo = {otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi = {otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi = {otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo = {otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo = {otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi = {otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo = {otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo = {otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi = {otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi = {otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi = {otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_hi_hi_lo_hi_hi = {otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo};
  wire [2047:0]       otherUnit_maskInput_lo_hi_hi_lo_hi = {otherUnit_maskInput_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_lo};
  wire [4095:0]       otherUnit_maskInput_lo_hi_hi_lo = {otherUnit_maskInput_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo = {otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi = {otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo = {otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo = {otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi = {otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo = {otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo = {otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi = {otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo = {otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo = {otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi = {otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_hi_hi_hi_lo_lo = {otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo = {otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi = {otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo = {otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo = {otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi = {otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo = {otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo = {otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi = {otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo = {otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo = {otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_hi_hi_hi_lo_hi = {otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo};
  wire [2047:0]       otherUnit_maskInput_lo_hi_hi_hi_lo = {otherUnit_maskInput_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo = {otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi = {otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo = {otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo = {otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi = {otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo = {otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo = {otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi = {otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo = {otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo = {otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi = {otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_hi_hi_hi_hi_lo = {otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo = {otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi = {otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo = {otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo = {otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi = {otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo = {otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo = {otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi = {otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo = {otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo = {otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_hi_hi_hi_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo};
  wire [2047:0]       otherUnit_maskInput_lo_hi_hi_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_lo};
  wire [4095:0]       otherUnit_maskInput_lo_hi_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_lo};
  wire [8191:0]       otherUnit_maskInput_lo_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_lo};
  wire [16383:0]      otherUnit_maskInput_lo_hi = {otherUnit_maskInput_lo_hi_hi, otherUnit_maskInput_lo_hi_lo};
  wire [32767:0]      otherUnit_maskInput_lo = {otherUnit_maskInput_lo_hi, otherUnit_maskInput_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo = {otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi = {otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo = {otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo = {otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi = {otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi = {otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo = {otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo = {otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi = {otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo = {otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo = {otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi = {otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi = {otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi = {otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_lo_lo_lo_lo_lo = {otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo = {otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi = {otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo = {otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo = {otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi = {otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi = {otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo = {otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo = {otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi = {otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo = {otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo = {otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi = {otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi = {otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi = {otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_lo_lo_lo_lo_hi = {otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo};
  wire [2047:0]       otherUnit_maskInput_hi_lo_lo_lo_lo = {otherUnit_maskInput_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo = {otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi = {otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo = {otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo = {otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi = {otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi = {otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo = {otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo = {otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi = {otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo = {otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo = {otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi = {otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi = {otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi = {otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_lo_lo_lo_hi_lo = {otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo = {otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi = {otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo = {otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo = {otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi = {otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi = {otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo = {otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo = {otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi = {otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo = {otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo = {otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi = {otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi = {otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi = {otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_lo_lo_lo_hi_hi = {otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo};
  wire [2047:0]       otherUnit_maskInput_hi_lo_lo_lo_hi = {otherUnit_maskInput_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_lo};
  wire [4095:0]       otherUnit_maskInput_hi_lo_lo_lo = {otherUnit_maskInput_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo = {otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi = {otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo = {otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo = {otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi = {otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi = {otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo = {otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo = {otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi = {otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo = {otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo = {otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi = {otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi = {otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi = {otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_lo_lo_hi_lo_lo = {otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo = {otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi = {otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo = {otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo = {otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi = {otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi = {otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo = {otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo = {otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi = {otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo = {otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo = {otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi = {otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi = {otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi = {otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_lo_lo_hi_lo_hi = {otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo};
  wire [2047:0]       otherUnit_maskInput_hi_lo_lo_hi_lo = {otherUnit_maskInput_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo = {otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi = {otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo = {otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo = {otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi = {otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi = {otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo = {otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo = {otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi = {otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo = {otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo = {otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi = {otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi = {otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi = {otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_lo_lo_hi_hi_lo = {otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo = {otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi = {otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo = {otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo = {otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi = {otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi = {otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo = {otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo = {otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi = {otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo = {otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo = {otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi = {otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi = {otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi = {otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_lo_lo_hi_hi_hi = {otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo};
  wire [2047:0]       otherUnit_maskInput_hi_lo_lo_hi_hi = {otherUnit_maskInput_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_lo};
  wire [4095:0]       otherUnit_maskInput_hi_lo_lo_hi = {otherUnit_maskInput_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_lo};
  wire [8191:0]       otherUnit_maskInput_hi_lo_lo = {otherUnit_maskInput_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo = {otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi = {otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo = {otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo = {otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi = {otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi = {otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo = {otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo = {otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo = {otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo = {otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi = {otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi = {otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi = {otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_lo_hi_lo_lo_lo = {otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo = {otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi = {otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo = {otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo = {otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi = {otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo = {otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo = {otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo = {otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo = {otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi = {otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi = {otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi = {otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_lo_hi_lo_lo_hi = {otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo};
  wire [2047:0]       otherUnit_maskInput_hi_lo_hi_lo_lo = {otherUnit_maskInput_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo = {otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi = {otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo = {otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo = {otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi = {otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi = {otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo = {otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo = {otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo = {otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo = {otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi = {otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi = {otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_lo_hi_lo_hi_lo = {otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo = {otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi = {otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo = {otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo = {otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi = {otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo = {otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo = {otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo = {otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo = {otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi = {otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi = {otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi = {otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_lo_hi_lo_hi_hi = {otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo};
  wire [2047:0]       otherUnit_maskInput_hi_lo_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_lo};
  wire [4095:0]       otherUnit_maskInput_hi_lo_hi_lo = {otherUnit_maskInput_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo = {otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi = {otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo = {otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo = {otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi = {otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi = {otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo = {otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo = {otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo = {otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo = {otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi = {otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi = {otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi = {otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_lo_hi_hi_lo_lo = {otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo = {otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi = {otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo = {otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo = {otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi = {otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo = {otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo = {otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo = {otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo = {otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi = {otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi = {otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi = {otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_lo_hi_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo};
  wire [2047:0]       otherUnit_maskInput_hi_lo_hi_hi_lo = {otherUnit_maskInput_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo = {otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi = {otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo = {otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo = {otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi = {otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi = {otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo = {otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo = {otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo = {otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo = {otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi = {otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi = {otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_lo_hi_hi_hi_lo = {otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo = {otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi = {otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo = {otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo = {otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi = {otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo = {otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo = {otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo = {otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo = {otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi = {otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi = {otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi = {otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_lo_hi_hi_hi_hi = {otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo};
  wire [2047:0]       otherUnit_maskInput_hi_lo_hi_hi_hi = {otherUnit_maskInput_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_lo};
  wire [4095:0]       otherUnit_maskInput_hi_lo_hi_hi = {otherUnit_maskInput_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_lo};
  wire [8191:0]       otherUnit_maskInput_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo};
  wire [16383:0]      otherUnit_maskInput_hi_lo = {otherUnit_maskInput_hi_lo_hi, otherUnit_maskInput_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo = {otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi = {otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo = {otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo = {otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi = {otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi = {otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo = {otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo = {otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi = {otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo = {otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo = {otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi = {otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi = {otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi = {otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_hi_lo_lo_lo_lo = {otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo = {otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi = {otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo = {otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo = {otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi = {otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi = {otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo = {otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo = {otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi = {otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo = {otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo = {otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi = {otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi = {otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi = {otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_hi_lo_lo_lo_hi = {otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo};
  wire [2047:0]       otherUnit_maskInput_hi_hi_lo_lo_lo = {otherUnit_maskInput_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo = {otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi = {otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo = {otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo = {otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi = {otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi = {otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo = {otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo = {otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi = {otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo = {otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo = {otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi = {otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi = {otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi = {otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_hi_lo_lo_hi_lo = {otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo = {otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi = {otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo = {otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo = {otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi = {otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi = {otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo = {otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo = {otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi = {otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo = {otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo = {otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi = {otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi = {otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi = {otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_hi_lo_lo_hi_hi = {otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo};
  wire [2047:0]       otherUnit_maskInput_hi_hi_lo_lo_hi = {otherUnit_maskInput_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_lo};
  wire [4095:0]       otherUnit_maskInput_hi_hi_lo_lo = {otherUnit_maskInput_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo = {otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi = {otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo = {otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi = {otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi = {otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo = {otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo = {otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi = {otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi = {otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi = {otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi = {otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_hi_lo_hi_lo_lo = {otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo = {otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi = {otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo = {otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi = {otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi = {otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo = {otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi = {otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi = {otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi = {otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi = {otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_hi_lo_hi_lo_hi = {otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo};
  wire [2047:0]       otherUnit_maskInput_hi_hi_lo_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo = {otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi = {otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo = {otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi = {otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi = {otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo = {otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo = {otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi = {otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi = {otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi = {otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi = {otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_hi_lo_hi_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo = {otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi = {otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo = {otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi = {otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi = {otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo = {otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi = {otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi = {otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi = {otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi = {otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_hi_lo_hi_hi_hi = {otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo};
  wire [2047:0]       otherUnit_maskInput_hi_hi_lo_hi_hi = {otherUnit_maskInput_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_lo};
  wire [4095:0]       otherUnit_maskInput_hi_hi_lo_hi = {otherUnit_maskInput_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_lo};
  wire [8191:0]       otherUnit_maskInput_hi_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo = {otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi = {otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo = {otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo = {otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi = {otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi = {otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo = {otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo = {otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi = {otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo = {otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo = {otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi = {otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi = {otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_hi_hi_lo_lo_lo = {otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo = {otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi = {otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo = {otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo = {otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi = {otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi = {otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo = {otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo = {otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi = {otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo = {otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo = {otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi = {otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_hi_hi_lo_lo_hi = {otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo};
  wire [2047:0]       otherUnit_maskInput_hi_hi_hi_lo_lo = {otherUnit_maskInput_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo = {otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi = {otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo = {otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo = {otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi = {otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi = {otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo = {otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo = {otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi = {otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo = {otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo = {otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi = {otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi = {otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_hi_hi_lo_hi_lo = {otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo = {otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi = {otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo = {otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo = {otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi = {otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi = {otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo = {otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo = {otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi = {otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo = {otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo = {otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_hi_hi_lo_hi_hi = {otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo};
  wire [2047:0]       otherUnit_maskInput_hi_hi_hi_lo_hi = {otherUnit_maskInput_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_lo};
  wire [4095:0]       otherUnit_maskInput_hi_hi_hi_lo = {otherUnit_maskInput_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo = {otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi = {otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo = {otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo = {otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi = {otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo = {otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo = {otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi = {otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo = {otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo = {otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi = {otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_hi_hi_hi_lo_lo = {otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo = {otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi = {otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo = {otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo = {otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi = {otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo = {otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo = {otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi = {otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo = {otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo = {otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_hi_hi_hi_lo_hi = {otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo};
  wire [2047:0]       otherUnit_maskInput_hi_hi_hi_hi_lo = {otherUnit_maskInput_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo = {otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi = {otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo = {otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo = {otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi = {otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo = {otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo = {otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi = {otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo = {otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo = {otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi = {otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_hi_hi_hi_hi_lo = {otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo = {otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi = {otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo = {otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo = {otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi = {otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo = {otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo = {otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi = {otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo = {otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo = {otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_hi_hi_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo};
  wire [2047:0]       otherUnit_maskInput_hi_hi_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_lo};
  wire [4095:0]       otherUnit_maskInput_hi_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_lo};
  wire [8191:0]       otherUnit_maskInput_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_lo};
  wire [16383:0]      otherUnit_maskInput_hi_hi = {otherUnit_maskInput_hi_hi_hi, otherUnit_maskInput_hi_hi_lo};
  wire [32767:0]      otherUnit_maskInput_hi = {otherUnit_maskInput_hi_hi, otherUnit_maskInput_hi_lo};
  wire [4095:0][15:0] _GEN_1025 =
    {{otherUnit_maskInput_hi[32767:32752]},
     {otherUnit_maskInput_hi[32751:32736]},
     {otherUnit_maskInput_hi[32735:32720]},
     {otherUnit_maskInput_hi[32719:32704]},
     {otherUnit_maskInput_hi[32703:32688]},
     {otherUnit_maskInput_hi[32687:32672]},
     {otherUnit_maskInput_hi[32671:32656]},
     {otherUnit_maskInput_hi[32655:32640]},
     {otherUnit_maskInput_hi[32639:32624]},
     {otherUnit_maskInput_hi[32623:32608]},
     {otherUnit_maskInput_hi[32607:32592]},
     {otherUnit_maskInput_hi[32591:32576]},
     {otherUnit_maskInput_hi[32575:32560]},
     {otherUnit_maskInput_hi[32559:32544]},
     {otherUnit_maskInput_hi[32543:32528]},
     {otherUnit_maskInput_hi[32527:32512]},
     {otherUnit_maskInput_hi[32511:32496]},
     {otherUnit_maskInput_hi[32495:32480]},
     {otherUnit_maskInput_hi[32479:32464]},
     {otherUnit_maskInput_hi[32463:32448]},
     {otherUnit_maskInput_hi[32447:32432]},
     {otherUnit_maskInput_hi[32431:32416]},
     {otherUnit_maskInput_hi[32415:32400]},
     {otherUnit_maskInput_hi[32399:32384]},
     {otherUnit_maskInput_hi[32383:32368]},
     {otherUnit_maskInput_hi[32367:32352]},
     {otherUnit_maskInput_hi[32351:32336]},
     {otherUnit_maskInput_hi[32335:32320]},
     {otherUnit_maskInput_hi[32319:32304]},
     {otherUnit_maskInput_hi[32303:32288]},
     {otherUnit_maskInput_hi[32287:32272]},
     {otherUnit_maskInput_hi[32271:32256]},
     {otherUnit_maskInput_hi[32255:32240]},
     {otherUnit_maskInput_hi[32239:32224]},
     {otherUnit_maskInput_hi[32223:32208]},
     {otherUnit_maskInput_hi[32207:32192]},
     {otherUnit_maskInput_hi[32191:32176]},
     {otherUnit_maskInput_hi[32175:32160]},
     {otherUnit_maskInput_hi[32159:32144]},
     {otherUnit_maskInput_hi[32143:32128]},
     {otherUnit_maskInput_hi[32127:32112]},
     {otherUnit_maskInput_hi[32111:32096]},
     {otherUnit_maskInput_hi[32095:32080]},
     {otherUnit_maskInput_hi[32079:32064]},
     {otherUnit_maskInput_hi[32063:32048]},
     {otherUnit_maskInput_hi[32047:32032]},
     {otherUnit_maskInput_hi[32031:32016]},
     {otherUnit_maskInput_hi[32015:32000]},
     {otherUnit_maskInput_hi[31999:31984]},
     {otherUnit_maskInput_hi[31983:31968]},
     {otherUnit_maskInput_hi[31967:31952]},
     {otherUnit_maskInput_hi[31951:31936]},
     {otherUnit_maskInput_hi[31935:31920]},
     {otherUnit_maskInput_hi[31919:31904]},
     {otherUnit_maskInput_hi[31903:31888]},
     {otherUnit_maskInput_hi[31887:31872]},
     {otherUnit_maskInput_hi[31871:31856]},
     {otherUnit_maskInput_hi[31855:31840]},
     {otherUnit_maskInput_hi[31839:31824]},
     {otherUnit_maskInput_hi[31823:31808]},
     {otherUnit_maskInput_hi[31807:31792]},
     {otherUnit_maskInput_hi[31791:31776]},
     {otherUnit_maskInput_hi[31775:31760]},
     {otherUnit_maskInput_hi[31759:31744]},
     {otherUnit_maskInput_hi[31743:31728]},
     {otherUnit_maskInput_hi[31727:31712]},
     {otherUnit_maskInput_hi[31711:31696]},
     {otherUnit_maskInput_hi[31695:31680]},
     {otherUnit_maskInput_hi[31679:31664]},
     {otherUnit_maskInput_hi[31663:31648]},
     {otherUnit_maskInput_hi[31647:31632]},
     {otherUnit_maskInput_hi[31631:31616]},
     {otherUnit_maskInput_hi[31615:31600]},
     {otherUnit_maskInput_hi[31599:31584]},
     {otherUnit_maskInput_hi[31583:31568]},
     {otherUnit_maskInput_hi[31567:31552]},
     {otherUnit_maskInput_hi[31551:31536]},
     {otherUnit_maskInput_hi[31535:31520]},
     {otherUnit_maskInput_hi[31519:31504]},
     {otherUnit_maskInput_hi[31503:31488]},
     {otherUnit_maskInput_hi[31487:31472]},
     {otherUnit_maskInput_hi[31471:31456]},
     {otherUnit_maskInput_hi[31455:31440]},
     {otherUnit_maskInput_hi[31439:31424]},
     {otherUnit_maskInput_hi[31423:31408]},
     {otherUnit_maskInput_hi[31407:31392]},
     {otherUnit_maskInput_hi[31391:31376]},
     {otherUnit_maskInput_hi[31375:31360]},
     {otherUnit_maskInput_hi[31359:31344]},
     {otherUnit_maskInput_hi[31343:31328]},
     {otherUnit_maskInput_hi[31327:31312]},
     {otherUnit_maskInput_hi[31311:31296]},
     {otherUnit_maskInput_hi[31295:31280]},
     {otherUnit_maskInput_hi[31279:31264]},
     {otherUnit_maskInput_hi[31263:31248]},
     {otherUnit_maskInput_hi[31247:31232]},
     {otherUnit_maskInput_hi[31231:31216]},
     {otherUnit_maskInput_hi[31215:31200]},
     {otherUnit_maskInput_hi[31199:31184]},
     {otherUnit_maskInput_hi[31183:31168]},
     {otherUnit_maskInput_hi[31167:31152]},
     {otherUnit_maskInput_hi[31151:31136]},
     {otherUnit_maskInput_hi[31135:31120]},
     {otherUnit_maskInput_hi[31119:31104]},
     {otherUnit_maskInput_hi[31103:31088]},
     {otherUnit_maskInput_hi[31087:31072]},
     {otherUnit_maskInput_hi[31071:31056]},
     {otherUnit_maskInput_hi[31055:31040]},
     {otherUnit_maskInput_hi[31039:31024]},
     {otherUnit_maskInput_hi[31023:31008]},
     {otherUnit_maskInput_hi[31007:30992]},
     {otherUnit_maskInput_hi[30991:30976]},
     {otherUnit_maskInput_hi[30975:30960]},
     {otherUnit_maskInput_hi[30959:30944]},
     {otherUnit_maskInput_hi[30943:30928]},
     {otherUnit_maskInput_hi[30927:30912]},
     {otherUnit_maskInput_hi[30911:30896]},
     {otherUnit_maskInput_hi[30895:30880]},
     {otherUnit_maskInput_hi[30879:30864]},
     {otherUnit_maskInput_hi[30863:30848]},
     {otherUnit_maskInput_hi[30847:30832]},
     {otherUnit_maskInput_hi[30831:30816]},
     {otherUnit_maskInput_hi[30815:30800]},
     {otherUnit_maskInput_hi[30799:30784]},
     {otherUnit_maskInput_hi[30783:30768]},
     {otherUnit_maskInput_hi[30767:30752]},
     {otherUnit_maskInput_hi[30751:30736]},
     {otherUnit_maskInput_hi[30735:30720]},
     {otherUnit_maskInput_hi[30719:30704]},
     {otherUnit_maskInput_hi[30703:30688]},
     {otherUnit_maskInput_hi[30687:30672]},
     {otherUnit_maskInput_hi[30671:30656]},
     {otherUnit_maskInput_hi[30655:30640]},
     {otherUnit_maskInput_hi[30639:30624]},
     {otherUnit_maskInput_hi[30623:30608]},
     {otherUnit_maskInput_hi[30607:30592]},
     {otherUnit_maskInput_hi[30591:30576]},
     {otherUnit_maskInput_hi[30575:30560]},
     {otherUnit_maskInput_hi[30559:30544]},
     {otherUnit_maskInput_hi[30543:30528]},
     {otherUnit_maskInput_hi[30527:30512]},
     {otherUnit_maskInput_hi[30511:30496]},
     {otherUnit_maskInput_hi[30495:30480]},
     {otherUnit_maskInput_hi[30479:30464]},
     {otherUnit_maskInput_hi[30463:30448]},
     {otherUnit_maskInput_hi[30447:30432]},
     {otherUnit_maskInput_hi[30431:30416]},
     {otherUnit_maskInput_hi[30415:30400]},
     {otherUnit_maskInput_hi[30399:30384]},
     {otherUnit_maskInput_hi[30383:30368]},
     {otherUnit_maskInput_hi[30367:30352]},
     {otherUnit_maskInput_hi[30351:30336]},
     {otherUnit_maskInput_hi[30335:30320]},
     {otherUnit_maskInput_hi[30319:30304]},
     {otherUnit_maskInput_hi[30303:30288]},
     {otherUnit_maskInput_hi[30287:30272]},
     {otherUnit_maskInput_hi[30271:30256]},
     {otherUnit_maskInput_hi[30255:30240]},
     {otherUnit_maskInput_hi[30239:30224]},
     {otherUnit_maskInput_hi[30223:30208]},
     {otherUnit_maskInput_hi[30207:30192]},
     {otherUnit_maskInput_hi[30191:30176]},
     {otherUnit_maskInput_hi[30175:30160]},
     {otherUnit_maskInput_hi[30159:30144]},
     {otherUnit_maskInput_hi[30143:30128]},
     {otherUnit_maskInput_hi[30127:30112]},
     {otherUnit_maskInput_hi[30111:30096]},
     {otherUnit_maskInput_hi[30095:30080]},
     {otherUnit_maskInput_hi[30079:30064]},
     {otherUnit_maskInput_hi[30063:30048]},
     {otherUnit_maskInput_hi[30047:30032]},
     {otherUnit_maskInput_hi[30031:30016]},
     {otherUnit_maskInput_hi[30015:30000]},
     {otherUnit_maskInput_hi[29999:29984]},
     {otherUnit_maskInput_hi[29983:29968]},
     {otherUnit_maskInput_hi[29967:29952]},
     {otherUnit_maskInput_hi[29951:29936]},
     {otherUnit_maskInput_hi[29935:29920]},
     {otherUnit_maskInput_hi[29919:29904]},
     {otherUnit_maskInput_hi[29903:29888]},
     {otherUnit_maskInput_hi[29887:29872]},
     {otherUnit_maskInput_hi[29871:29856]},
     {otherUnit_maskInput_hi[29855:29840]},
     {otherUnit_maskInput_hi[29839:29824]},
     {otherUnit_maskInput_hi[29823:29808]},
     {otherUnit_maskInput_hi[29807:29792]},
     {otherUnit_maskInput_hi[29791:29776]},
     {otherUnit_maskInput_hi[29775:29760]},
     {otherUnit_maskInput_hi[29759:29744]},
     {otherUnit_maskInput_hi[29743:29728]},
     {otherUnit_maskInput_hi[29727:29712]},
     {otherUnit_maskInput_hi[29711:29696]},
     {otherUnit_maskInput_hi[29695:29680]},
     {otherUnit_maskInput_hi[29679:29664]},
     {otherUnit_maskInput_hi[29663:29648]},
     {otherUnit_maskInput_hi[29647:29632]},
     {otherUnit_maskInput_hi[29631:29616]},
     {otherUnit_maskInput_hi[29615:29600]},
     {otherUnit_maskInput_hi[29599:29584]},
     {otherUnit_maskInput_hi[29583:29568]},
     {otherUnit_maskInput_hi[29567:29552]},
     {otherUnit_maskInput_hi[29551:29536]},
     {otherUnit_maskInput_hi[29535:29520]},
     {otherUnit_maskInput_hi[29519:29504]},
     {otherUnit_maskInput_hi[29503:29488]},
     {otherUnit_maskInput_hi[29487:29472]},
     {otherUnit_maskInput_hi[29471:29456]},
     {otherUnit_maskInput_hi[29455:29440]},
     {otherUnit_maskInput_hi[29439:29424]},
     {otherUnit_maskInput_hi[29423:29408]},
     {otherUnit_maskInput_hi[29407:29392]},
     {otherUnit_maskInput_hi[29391:29376]},
     {otherUnit_maskInput_hi[29375:29360]},
     {otherUnit_maskInput_hi[29359:29344]},
     {otherUnit_maskInput_hi[29343:29328]},
     {otherUnit_maskInput_hi[29327:29312]},
     {otherUnit_maskInput_hi[29311:29296]},
     {otherUnit_maskInput_hi[29295:29280]},
     {otherUnit_maskInput_hi[29279:29264]},
     {otherUnit_maskInput_hi[29263:29248]},
     {otherUnit_maskInput_hi[29247:29232]},
     {otherUnit_maskInput_hi[29231:29216]},
     {otherUnit_maskInput_hi[29215:29200]},
     {otherUnit_maskInput_hi[29199:29184]},
     {otherUnit_maskInput_hi[29183:29168]},
     {otherUnit_maskInput_hi[29167:29152]},
     {otherUnit_maskInput_hi[29151:29136]},
     {otherUnit_maskInput_hi[29135:29120]},
     {otherUnit_maskInput_hi[29119:29104]},
     {otherUnit_maskInput_hi[29103:29088]},
     {otherUnit_maskInput_hi[29087:29072]},
     {otherUnit_maskInput_hi[29071:29056]},
     {otherUnit_maskInput_hi[29055:29040]},
     {otherUnit_maskInput_hi[29039:29024]},
     {otherUnit_maskInput_hi[29023:29008]},
     {otherUnit_maskInput_hi[29007:28992]},
     {otherUnit_maskInput_hi[28991:28976]},
     {otherUnit_maskInput_hi[28975:28960]},
     {otherUnit_maskInput_hi[28959:28944]},
     {otherUnit_maskInput_hi[28943:28928]},
     {otherUnit_maskInput_hi[28927:28912]},
     {otherUnit_maskInput_hi[28911:28896]},
     {otherUnit_maskInput_hi[28895:28880]},
     {otherUnit_maskInput_hi[28879:28864]},
     {otherUnit_maskInput_hi[28863:28848]},
     {otherUnit_maskInput_hi[28847:28832]},
     {otherUnit_maskInput_hi[28831:28816]},
     {otherUnit_maskInput_hi[28815:28800]},
     {otherUnit_maskInput_hi[28799:28784]},
     {otherUnit_maskInput_hi[28783:28768]},
     {otherUnit_maskInput_hi[28767:28752]},
     {otherUnit_maskInput_hi[28751:28736]},
     {otherUnit_maskInput_hi[28735:28720]},
     {otherUnit_maskInput_hi[28719:28704]},
     {otherUnit_maskInput_hi[28703:28688]},
     {otherUnit_maskInput_hi[28687:28672]},
     {otherUnit_maskInput_hi[28671:28656]},
     {otherUnit_maskInput_hi[28655:28640]},
     {otherUnit_maskInput_hi[28639:28624]},
     {otherUnit_maskInput_hi[28623:28608]},
     {otherUnit_maskInput_hi[28607:28592]},
     {otherUnit_maskInput_hi[28591:28576]},
     {otherUnit_maskInput_hi[28575:28560]},
     {otherUnit_maskInput_hi[28559:28544]},
     {otherUnit_maskInput_hi[28543:28528]},
     {otherUnit_maskInput_hi[28527:28512]},
     {otherUnit_maskInput_hi[28511:28496]},
     {otherUnit_maskInput_hi[28495:28480]},
     {otherUnit_maskInput_hi[28479:28464]},
     {otherUnit_maskInput_hi[28463:28448]},
     {otherUnit_maskInput_hi[28447:28432]},
     {otherUnit_maskInput_hi[28431:28416]},
     {otherUnit_maskInput_hi[28415:28400]},
     {otherUnit_maskInput_hi[28399:28384]},
     {otherUnit_maskInput_hi[28383:28368]},
     {otherUnit_maskInput_hi[28367:28352]},
     {otherUnit_maskInput_hi[28351:28336]},
     {otherUnit_maskInput_hi[28335:28320]},
     {otherUnit_maskInput_hi[28319:28304]},
     {otherUnit_maskInput_hi[28303:28288]},
     {otherUnit_maskInput_hi[28287:28272]},
     {otherUnit_maskInput_hi[28271:28256]},
     {otherUnit_maskInput_hi[28255:28240]},
     {otherUnit_maskInput_hi[28239:28224]},
     {otherUnit_maskInput_hi[28223:28208]},
     {otherUnit_maskInput_hi[28207:28192]},
     {otherUnit_maskInput_hi[28191:28176]},
     {otherUnit_maskInput_hi[28175:28160]},
     {otherUnit_maskInput_hi[28159:28144]},
     {otherUnit_maskInput_hi[28143:28128]},
     {otherUnit_maskInput_hi[28127:28112]},
     {otherUnit_maskInput_hi[28111:28096]},
     {otherUnit_maskInput_hi[28095:28080]},
     {otherUnit_maskInput_hi[28079:28064]},
     {otherUnit_maskInput_hi[28063:28048]},
     {otherUnit_maskInput_hi[28047:28032]},
     {otherUnit_maskInput_hi[28031:28016]},
     {otherUnit_maskInput_hi[28015:28000]},
     {otherUnit_maskInput_hi[27999:27984]},
     {otherUnit_maskInput_hi[27983:27968]},
     {otherUnit_maskInput_hi[27967:27952]},
     {otherUnit_maskInput_hi[27951:27936]},
     {otherUnit_maskInput_hi[27935:27920]},
     {otherUnit_maskInput_hi[27919:27904]},
     {otherUnit_maskInput_hi[27903:27888]},
     {otherUnit_maskInput_hi[27887:27872]},
     {otherUnit_maskInput_hi[27871:27856]},
     {otherUnit_maskInput_hi[27855:27840]},
     {otherUnit_maskInput_hi[27839:27824]},
     {otherUnit_maskInput_hi[27823:27808]},
     {otherUnit_maskInput_hi[27807:27792]},
     {otherUnit_maskInput_hi[27791:27776]},
     {otherUnit_maskInput_hi[27775:27760]},
     {otherUnit_maskInput_hi[27759:27744]},
     {otherUnit_maskInput_hi[27743:27728]},
     {otherUnit_maskInput_hi[27727:27712]},
     {otherUnit_maskInput_hi[27711:27696]},
     {otherUnit_maskInput_hi[27695:27680]},
     {otherUnit_maskInput_hi[27679:27664]},
     {otherUnit_maskInput_hi[27663:27648]},
     {otherUnit_maskInput_hi[27647:27632]},
     {otherUnit_maskInput_hi[27631:27616]},
     {otherUnit_maskInput_hi[27615:27600]},
     {otherUnit_maskInput_hi[27599:27584]},
     {otherUnit_maskInput_hi[27583:27568]},
     {otherUnit_maskInput_hi[27567:27552]},
     {otherUnit_maskInput_hi[27551:27536]},
     {otherUnit_maskInput_hi[27535:27520]},
     {otherUnit_maskInput_hi[27519:27504]},
     {otherUnit_maskInput_hi[27503:27488]},
     {otherUnit_maskInput_hi[27487:27472]},
     {otherUnit_maskInput_hi[27471:27456]},
     {otherUnit_maskInput_hi[27455:27440]},
     {otherUnit_maskInput_hi[27439:27424]},
     {otherUnit_maskInput_hi[27423:27408]},
     {otherUnit_maskInput_hi[27407:27392]},
     {otherUnit_maskInput_hi[27391:27376]},
     {otherUnit_maskInput_hi[27375:27360]},
     {otherUnit_maskInput_hi[27359:27344]},
     {otherUnit_maskInput_hi[27343:27328]},
     {otherUnit_maskInput_hi[27327:27312]},
     {otherUnit_maskInput_hi[27311:27296]},
     {otherUnit_maskInput_hi[27295:27280]},
     {otherUnit_maskInput_hi[27279:27264]},
     {otherUnit_maskInput_hi[27263:27248]},
     {otherUnit_maskInput_hi[27247:27232]},
     {otherUnit_maskInput_hi[27231:27216]},
     {otherUnit_maskInput_hi[27215:27200]},
     {otherUnit_maskInput_hi[27199:27184]},
     {otherUnit_maskInput_hi[27183:27168]},
     {otherUnit_maskInput_hi[27167:27152]},
     {otherUnit_maskInput_hi[27151:27136]},
     {otherUnit_maskInput_hi[27135:27120]},
     {otherUnit_maskInput_hi[27119:27104]},
     {otherUnit_maskInput_hi[27103:27088]},
     {otherUnit_maskInput_hi[27087:27072]},
     {otherUnit_maskInput_hi[27071:27056]},
     {otherUnit_maskInput_hi[27055:27040]},
     {otherUnit_maskInput_hi[27039:27024]},
     {otherUnit_maskInput_hi[27023:27008]},
     {otherUnit_maskInput_hi[27007:26992]},
     {otherUnit_maskInput_hi[26991:26976]},
     {otherUnit_maskInput_hi[26975:26960]},
     {otherUnit_maskInput_hi[26959:26944]},
     {otherUnit_maskInput_hi[26943:26928]},
     {otherUnit_maskInput_hi[26927:26912]},
     {otherUnit_maskInput_hi[26911:26896]},
     {otherUnit_maskInput_hi[26895:26880]},
     {otherUnit_maskInput_hi[26879:26864]},
     {otherUnit_maskInput_hi[26863:26848]},
     {otherUnit_maskInput_hi[26847:26832]},
     {otherUnit_maskInput_hi[26831:26816]},
     {otherUnit_maskInput_hi[26815:26800]},
     {otherUnit_maskInput_hi[26799:26784]},
     {otherUnit_maskInput_hi[26783:26768]},
     {otherUnit_maskInput_hi[26767:26752]},
     {otherUnit_maskInput_hi[26751:26736]},
     {otherUnit_maskInput_hi[26735:26720]},
     {otherUnit_maskInput_hi[26719:26704]},
     {otherUnit_maskInput_hi[26703:26688]},
     {otherUnit_maskInput_hi[26687:26672]},
     {otherUnit_maskInput_hi[26671:26656]},
     {otherUnit_maskInput_hi[26655:26640]},
     {otherUnit_maskInput_hi[26639:26624]},
     {otherUnit_maskInput_hi[26623:26608]},
     {otherUnit_maskInput_hi[26607:26592]},
     {otherUnit_maskInput_hi[26591:26576]},
     {otherUnit_maskInput_hi[26575:26560]},
     {otherUnit_maskInput_hi[26559:26544]},
     {otherUnit_maskInput_hi[26543:26528]},
     {otherUnit_maskInput_hi[26527:26512]},
     {otherUnit_maskInput_hi[26511:26496]},
     {otherUnit_maskInput_hi[26495:26480]},
     {otherUnit_maskInput_hi[26479:26464]},
     {otherUnit_maskInput_hi[26463:26448]},
     {otherUnit_maskInput_hi[26447:26432]},
     {otherUnit_maskInput_hi[26431:26416]},
     {otherUnit_maskInput_hi[26415:26400]},
     {otherUnit_maskInput_hi[26399:26384]},
     {otherUnit_maskInput_hi[26383:26368]},
     {otherUnit_maskInput_hi[26367:26352]},
     {otherUnit_maskInput_hi[26351:26336]},
     {otherUnit_maskInput_hi[26335:26320]},
     {otherUnit_maskInput_hi[26319:26304]},
     {otherUnit_maskInput_hi[26303:26288]},
     {otherUnit_maskInput_hi[26287:26272]},
     {otherUnit_maskInput_hi[26271:26256]},
     {otherUnit_maskInput_hi[26255:26240]},
     {otherUnit_maskInput_hi[26239:26224]},
     {otherUnit_maskInput_hi[26223:26208]},
     {otherUnit_maskInput_hi[26207:26192]},
     {otherUnit_maskInput_hi[26191:26176]},
     {otherUnit_maskInput_hi[26175:26160]},
     {otherUnit_maskInput_hi[26159:26144]},
     {otherUnit_maskInput_hi[26143:26128]},
     {otherUnit_maskInput_hi[26127:26112]},
     {otherUnit_maskInput_hi[26111:26096]},
     {otherUnit_maskInput_hi[26095:26080]},
     {otherUnit_maskInput_hi[26079:26064]},
     {otherUnit_maskInput_hi[26063:26048]},
     {otherUnit_maskInput_hi[26047:26032]},
     {otherUnit_maskInput_hi[26031:26016]},
     {otherUnit_maskInput_hi[26015:26000]},
     {otherUnit_maskInput_hi[25999:25984]},
     {otherUnit_maskInput_hi[25983:25968]},
     {otherUnit_maskInput_hi[25967:25952]},
     {otherUnit_maskInput_hi[25951:25936]},
     {otherUnit_maskInput_hi[25935:25920]},
     {otherUnit_maskInput_hi[25919:25904]},
     {otherUnit_maskInput_hi[25903:25888]},
     {otherUnit_maskInput_hi[25887:25872]},
     {otherUnit_maskInput_hi[25871:25856]},
     {otherUnit_maskInput_hi[25855:25840]},
     {otherUnit_maskInput_hi[25839:25824]},
     {otherUnit_maskInput_hi[25823:25808]},
     {otherUnit_maskInput_hi[25807:25792]},
     {otherUnit_maskInput_hi[25791:25776]},
     {otherUnit_maskInput_hi[25775:25760]},
     {otherUnit_maskInput_hi[25759:25744]},
     {otherUnit_maskInput_hi[25743:25728]},
     {otherUnit_maskInput_hi[25727:25712]},
     {otherUnit_maskInput_hi[25711:25696]},
     {otherUnit_maskInput_hi[25695:25680]},
     {otherUnit_maskInput_hi[25679:25664]},
     {otherUnit_maskInput_hi[25663:25648]},
     {otherUnit_maskInput_hi[25647:25632]},
     {otherUnit_maskInput_hi[25631:25616]},
     {otherUnit_maskInput_hi[25615:25600]},
     {otherUnit_maskInput_hi[25599:25584]},
     {otherUnit_maskInput_hi[25583:25568]},
     {otherUnit_maskInput_hi[25567:25552]},
     {otherUnit_maskInput_hi[25551:25536]},
     {otherUnit_maskInput_hi[25535:25520]},
     {otherUnit_maskInput_hi[25519:25504]},
     {otherUnit_maskInput_hi[25503:25488]},
     {otherUnit_maskInput_hi[25487:25472]},
     {otherUnit_maskInput_hi[25471:25456]},
     {otherUnit_maskInput_hi[25455:25440]},
     {otherUnit_maskInput_hi[25439:25424]},
     {otherUnit_maskInput_hi[25423:25408]},
     {otherUnit_maskInput_hi[25407:25392]},
     {otherUnit_maskInput_hi[25391:25376]},
     {otherUnit_maskInput_hi[25375:25360]},
     {otherUnit_maskInput_hi[25359:25344]},
     {otherUnit_maskInput_hi[25343:25328]},
     {otherUnit_maskInput_hi[25327:25312]},
     {otherUnit_maskInput_hi[25311:25296]},
     {otherUnit_maskInput_hi[25295:25280]},
     {otherUnit_maskInput_hi[25279:25264]},
     {otherUnit_maskInput_hi[25263:25248]},
     {otherUnit_maskInput_hi[25247:25232]},
     {otherUnit_maskInput_hi[25231:25216]},
     {otherUnit_maskInput_hi[25215:25200]},
     {otherUnit_maskInput_hi[25199:25184]},
     {otherUnit_maskInput_hi[25183:25168]},
     {otherUnit_maskInput_hi[25167:25152]},
     {otherUnit_maskInput_hi[25151:25136]},
     {otherUnit_maskInput_hi[25135:25120]},
     {otherUnit_maskInput_hi[25119:25104]},
     {otherUnit_maskInput_hi[25103:25088]},
     {otherUnit_maskInput_hi[25087:25072]},
     {otherUnit_maskInput_hi[25071:25056]},
     {otherUnit_maskInput_hi[25055:25040]},
     {otherUnit_maskInput_hi[25039:25024]},
     {otherUnit_maskInput_hi[25023:25008]},
     {otherUnit_maskInput_hi[25007:24992]},
     {otherUnit_maskInput_hi[24991:24976]},
     {otherUnit_maskInput_hi[24975:24960]},
     {otherUnit_maskInput_hi[24959:24944]},
     {otherUnit_maskInput_hi[24943:24928]},
     {otherUnit_maskInput_hi[24927:24912]},
     {otherUnit_maskInput_hi[24911:24896]},
     {otherUnit_maskInput_hi[24895:24880]},
     {otherUnit_maskInput_hi[24879:24864]},
     {otherUnit_maskInput_hi[24863:24848]},
     {otherUnit_maskInput_hi[24847:24832]},
     {otherUnit_maskInput_hi[24831:24816]},
     {otherUnit_maskInput_hi[24815:24800]},
     {otherUnit_maskInput_hi[24799:24784]},
     {otherUnit_maskInput_hi[24783:24768]},
     {otherUnit_maskInput_hi[24767:24752]},
     {otherUnit_maskInput_hi[24751:24736]},
     {otherUnit_maskInput_hi[24735:24720]},
     {otherUnit_maskInput_hi[24719:24704]},
     {otherUnit_maskInput_hi[24703:24688]},
     {otherUnit_maskInput_hi[24687:24672]},
     {otherUnit_maskInput_hi[24671:24656]},
     {otherUnit_maskInput_hi[24655:24640]},
     {otherUnit_maskInput_hi[24639:24624]},
     {otherUnit_maskInput_hi[24623:24608]},
     {otherUnit_maskInput_hi[24607:24592]},
     {otherUnit_maskInput_hi[24591:24576]},
     {otherUnit_maskInput_hi[24575:24560]},
     {otherUnit_maskInput_hi[24559:24544]},
     {otherUnit_maskInput_hi[24543:24528]},
     {otherUnit_maskInput_hi[24527:24512]},
     {otherUnit_maskInput_hi[24511:24496]},
     {otherUnit_maskInput_hi[24495:24480]},
     {otherUnit_maskInput_hi[24479:24464]},
     {otherUnit_maskInput_hi[24463:24448]},
     {otherUnit_maskInput_hi[24447:24432]},
     {otherUnit_maskInput_hi[24431:24416]},
     {otherUnit_maskInput_hi[24415:24400]},
     {otherUnit_maskInput_hi[24399:24384]},
     {otherUnit_maskInput_hi[24383:24368]},
     {otherUnit_maskInput_hi[24367:24352]},
     {otherUnit_maskInput_hi[24351:24336]},
     {otherUnit_maskInput_hi[24335:24320]},
     {otherUnit_maskInput_hi[24319:24304]},
     {otherUnit_maskInput_hi[24303:24288]},
     {otherUnit_maskInput_hi[24287:24272]},
     {otherUnit_maskInput_hi[24271:24256]},
     {otherUnit_maskInput_hi[24255:24240]},
     {otherUnit_maskInput_hi[24239:24224]},
     {otherUnit_maskInput_hi[24223:24208]},
     {otherUnit_maskInput_hi[24207:24192]},
     {otherUnit_maskInput_hi[24191:24176]},
     {otherUnit_maskInput_hi[24175:24160]},
     {otherUnit_maskInput_hi[24159:24144]},
     {otherUnit_maskInput_hi[24143:24128]},
     {otherUnit_maskInput_hi[24127:24112]},
     {otherUnit_maskInput_hi[24111:24096]},
     {otherUnit_maskInput_hi[24095:24080]},
     {otherUnit_maskInput_hi[24079:24064]},
     {otherUnit_maskInput_hi[24063:24048]},
     {otherUnit_maskInput_hi[24047:24032]},
     {otherUnit_maskInput_hi[24031:24016]},
     {otherUnit_maskInput_hi[24015:24000]},
     {otherUnit_maskInput_hi[23999:23984]},
     {otherUnit_maskInput_hi[23983:23968]},
     {otherUnit_maskInput_hi[23967:23952]},
     {otherUnit_maskInput_hi[23951:23936]},
     {otherUnit_maskInput_hi[23935:23920]},
     {otherUnit_maskInput_hi[23919:23904]},
     {otherUnit_maskInput_hi[23903:23888]},
     {otherUnit_maskInput_hi[23887:23872]},
     {otherUnit_maskInput_hi[23871:23856]},
     {otherUnit_maskInput_hi[23855:23840]},
     {otherUnit_maskInput_hi[23839:23824]},
     {otherUnit_maskInput_hi[23823:23808]},
     {otherUnit_maskInput_hi[23807:23792]},
     {otherUnit_maskInput_hi[23791:23776]},
     {otherUnit_maskInput_hi[23775:23760]},
     {otherUnit_maskInput_hi[23759:23744]},
     {otherUnit_maskInput_hi[23743:23728]},
     {otherUnit_maskInput_hi[23727:23712]},
     {otherUnit_maskInput_hi[23711:23696]},
     {otherUnit_maskInput_hi[23695:23680]},
     {otherUnit_maskInput_hi[23679:23664]},
     {otherUnit_maskInput_hi[23663:23648]},
     {otherUnit_maskInput_hi[23647:23632]},
     {otherUnit_maskInput_hi[23631:23616]},
     {otherUnit_maskInput_hi[23615:23600]},
     {otherUnit_maskInput_hi[23599:23584]},
     {otherUnit_maskInput_hi[23583:23568]},
     {otherUnit_maskInput_hi[23567:23552]},
     {otherUnit_maskInput_hi[23551:23536]},
     {otherUnit_maskInput_hi[23535:23520]},
     {otherUnit_maskInput_hi[23519:23504]},
     {otherUnit_maskInput_hi[23503:23488]},
     {otherUnit_maskInput_hi[23487:23472]},
     {otherUnit_maskInput_hi[23471:23456]},
     {otherUnit_maskInput_hi[23455:23440]},
     {otherUnit_maskInput_hi[23439:23424]},
     {otherUnit_maskInput_hi[23423:23408]},
     {otherUnit_maskInput_hi[23407:23392]},
     {otherUnit_maskInput_hi[23391:23376]},
     {otherUnit_maskInput_hi[23375:23360]},
     {otherUnit_maskInput_hi[23359:23344]},
     {otherUnit_maskInput_hi[23343:23328]},
     {otherUnit_maskInput_hi[23327:23312]},
     {otherUnit_maskInput_hi[23311:23296]},
     {otherUnit_maskInput_hi[23295:23280]},
     {otherUnit_maskInput_hi[23279:23264]},
     {otherUnit_maskInput_hi[23263:23248]},
     {otherUnit_maskInput_hi[23247:23232]},
     {otherUnit_maskInput_hi[23231:23216]},
     {otherUnit_maskInput_hi[23215:23200]},
     {otherUnit_maskInput_hi[23199:23184]},
     {otherUnit_maskInput_hi[23183:23168]},
     {otherUnit_maskInput_hi[23167:23152]},
     {otherUnit_maskInput_hi[23151:23136]},
     {otherUnit_maskInput_hi[23135:23120]},
     {otherUnit_maskInput_hi[23119:23104]},
     {otherUnit_maskInput_hi[23103:23088]},
     {otherUnit_maskInput_hi[23087:23072]},
     {otherUnit_maskInput_hi[23071:23056]},
     {otherUnit_maskInput_hi[23055:23040]},
     {otherUnit_maskInput_hi[23039:23024]},
     {otherUnit_maskInput_hi[23023:23008]},
     {otherUnit_maskInput_hi[23007:22992]},
     {otherUnit_maskInput_hi[22991:22976]},
     {otherUnit_maskInput_hi[22975:22960]},
     {otherUnit_maskInput_hi[22959:22944]},
     {otherUnit_maskInput_hi[22943:22928]},
     {otherUnit_maskInput_hi[22927:22912]},
     {otherUnit_maskInput_hi[22911:22896]},
     {otherUnit_maskInput_hi[22895:22880]},
     {otherUnit_maskInput_hi[22879:22864]},
     {otherUnit_maskInput_hi[22863:22848]},
     {otherUnit_maskInput_hi[22847:22832]},
     {otherUnit_maskInput_hi[22831:22816]},
     {otherUnit_maskInput_hi[22815:22800]},
     {otherUnit_maskInput_hi[22799:22784]},
     {otherUnit_maskInput_hi[22783:22768]},
     {otherUnit_maskInput_hi[22767:22752]},
     {otherUnit_maskInput_hi[22751:22736]},
     {otherUnit_maskInput_hi[22735:22720]},
     {otherUnit_maskInput_hi[22719:22704]},
     {otherUnit_maskInput_hi[22703:22688]},
     {otherUnit_maskInput_hi[22687:22672]},
     {otherUnit_maskInput_hi[22671:22656]},
     {otherUnit_maskInput_hi[22655:22640]},
     {otherUnit_maskInput_hi[22639:22624]},
     {otherUnit_maskInput_hi[22623:22608]},
     {otherUnit_maskInput_hi[22607:22592]},
     {otherUnit_maskInput_hi[22591:22576]},
     {otherUnit_maskInput_hi[22575:22560]},
     {otherUnit_maskInput_hi[22559:22544]},
     {otherUnit_maskInput_hi[22543:22528]},
     {otherUnit_maskInput_hi[22527:22512]},
     {otherUnit_maskInput_hi[22511:22496]},
     {otherUnit_maskInput_hi[22495:22480]},
     {otherUnit_maskInput_hi[22479:22464]},
     {otherUnit_maskInput_hi[22463:22448]},
     {otherUnit_maskInput_hi[22447:22432]},
     {otherUnit_maskInput_hi[22431:22416]},
     {otherUnit_maskInput_hi[22415:22400]},
     {otherUnit_maskInput_hi[22399:22384]},
     {otherUnit_maskInput_hi[22383:22368]},
     {otherUnit_maskInput_hi[22367:22352]},
     {otherUnit_maskInput_hi[22351:22336]},
     {otherUnit_maskInput_hi[22335:22320]},
     {otherUnit_maskInput_hi[22319:22304]},
     {otherUnit_maskInput_hi[22303:22288]},
     {otherUnit_maskInput_hi[22287:22272]},
     {otherUnit_maskInput_hi[22271:22256]},
     {otherUnit_maskInput_hi[22255:22240]},
     {otherUnit_maskInput_hi[22239:22224]},
     {otherUnit_maskInput_hi[22223:22208]},
     {otherUnit_maskInput_hi[22207:22192]},
     {otherUnit_maskInput_hi[22191:22176]},
     {otherUnit_maskInput_hi[22175:22160]},
     {otherUnit_maskInput_hi[22159:22144]},
     {otherUnit_maskInput_hi[22143:22128]},
     {otherUnit_maskInput_hi[22127:22112]},
     {otherUnit_maskInput_hi[22111:22096]},
     {otherUnit_maskInput_hi[22095:22080]},
     {otherUnit_maskInput_hi[22079:22064]},
     {otherUnit_maskInput_hi[22063:22048]},
     {otherUnit_maskInput_hi[22047:22032]},
     {otherUnit_maskInput_hi[22031:22016]},
     {otherUnit_maskInput_hi[22015:22000]},
     {otherUnit_maskInput_hi[21999:21984]},
     {otherUnit_maskInput_hi[21983:21968]},
     {otherUnit_maskInput_hi[21967:21952]},
     {otherUnit_maskInput_hi[21951:21936]},
     {otherUnit_maskInput_hi[21935:21920]},
     {otherUnit_maskInput_hi[21919:21904]},
     {otherUnit_maskInput_hi[21903:21888]},
     {otherUnit_maskInput_hi[21887:21872]},
     {otherUnit_maskInput_hi[21871:21856]},
     {otherUnit_maskInput_hi[21855:21840]},
     {otherUnit_maskInput_hi[21839:21824]},
     {otherUnit_maskInput_hi[21823:21808]},
     {otherUnit_maskInput_hi[21807:21792]},
     {otherUnit_maskInput_hi[21791:21776]},
     {otherUnit_maskInput_hi[21775:21760]},
     {otherUnit_maskInput_hi[21759:21744]},
     {otherUnit_maskInput_hi[21743:21728]},
     {otherUnit_maskInput_hi[21727:21712]},
     {otherUnit_maskInput_hi[21711:21696]},
     {otherUnit_maskInput_hi[21695:21680]},
     {otherUnit_maskInput_hi[21679:21664]},
     {otherUnit_maskInput_hi[21663:21648]},
     {otherUnit_maskInput_hi[21647:21632]},
     {otherUnit_maskInput_hi[21631:21616]},
     {otherUnit_maskInput_hi[21615:21600]},
     {otherUnit_maskInput_hi[21599:21584]},
     {otherUnit_maskInput_hi[21583:21568]},
     {otherUnit_maskInput_hi[21567:21552]},
     {otherUnit_maskInput_hi[21551:21536]},
     {otherUnit_maskInput_hi[21535:21520]},
     {otherUnit_maskInput_hi[21519:21504]},
     {otherUnit_maskInput_hi[21503:21488]},
     {otherUnit_maskInput_hi[21487:21472]},
     {otherUnit_maskInput_hi[21471:21456]},
     {otherUnit_maskInput_hi[21455:21440]},
     {otherUnit_maskInput_hi[21439:21424]},
     {otherUnit_maskInput_hi[21423:21408]},
     {otherUnit_maskInput_hi[21407:21392]},
     {otherUnit_maskInput_hi[21391:21376]},
     {otherUnit_maskInput_hi[21375:21360]},
     {otherUnit_maskInput_hi[21359:21344]},
     {otherUnit_maskInput_hi[21343:21328]},
     {otherUnit_maskInput_hi[21327:21312]},
     {otherUnit_maskInput_hi[21311:21296]},
     {otherUnit_maskInput_hi[21295:21280]},
     {otherUnit_maskInput_hi[21279:21264]},
     {otherUnit_maskInput_hi[21263:21248]},
     {otherUnit_maskInput_hi[21247:21232]},
     {otherUnit_maskInput_hi[21231:21216]},
     {otherUnit_maskInput_hi[21215:21200]},
     {otherUnit_maskInput_hi[21199:21184]},
     {otherUnit_maskInput_hi[21183:21168]},
     {otherUnit_maskInput_hi[21167:21152]},
     {otherUnit_maskInput_hi[21151:21136]},
     {otherUnit_maskInput_hi[21135:21120]},
     {otherUnit_maskInput_hi[21119:21104]},
     {otherUnit_maskInput_hi[21103:21088]},
     {otherUnit_maskInput_hi[21087:21072]},
     {otherUnit_maskInput_hi[21071:21056]},
     {otherUnit_maskInput_hi[21055:21040]},
     {otherUnit_maskInput_hi[21039:21024]},
     {otherUnit_maskInput_hi[21023:21008]},
     {otherUnit_maskInput_hi[21007:20992]},
     {otherUnit_maskInput_hi[20991:20976]},
     {otherUnit_maskInput_hi[20975:20960]},
     {otherUnit_maskInput_hi[20959:20944]},
     {otherUnit_maskInput_hi[20943:20928]},
     {otherUnit_maskInput_hi[20927:20912]},
     {otherUnit_maskInput_hi[20911:20896]},
     {otherUnit_maskInput_hi[20895:20880]},
     {otherUnit_maskInput_hi[20879:20864]},
     {otherUnit_maskInput_hi[20863:20848]},
     {otherUnit_maskInput_hi[20847:20832]},
     {otherUnit_maskInput_hi[20831:20816]},
     {otherUnit_maskInput_hi[20815:20800]},
     {otherUnit_maskInput_hi[20799:20784]},
     {otherUnit_maskInput_hi[20783:20768]},
     {otherUnit_maskInput_hi[20767:20752]},
     {otherUnit_maskInput_hi[20751:20736]},
     {otherUnit_maskInput_hi[20735:20720]},
     {otherUnit_maskInput_hi[20719:20704]},
     {otherUnit_maskInput_hi[20703:20688]},
     {otherUnit_maskInput_hi[20687:20672]},
     {otherUnit_maskInput_hi[20671:20656]},
     {otherUnit_maskInput_hi[20655:20640]},
     {otherUnit_maskInput_hi[20639:20624]},
     {otherUnit_maskInput_hi[20623:20608]},
     {otherUnit_maskInput_hi[20607:20592]},
     {otherUnit_maskInput_hi[20591:20576]},
     {otherUnit_maskInput_hi[20575:20560]},
     {otherUnit_maskInput_hi[20559:20544]},
     {otherUnit_maskInput_hi[20543:20528]},
     {otherUnit_maskInput_hi[20527:20512]},
     {otherUnit_maskInput_hi[20511:20496]},
     {otherUnit_maskInput_hi[20495:20480]},
     {otherUnit_maskInput_hi[20479:20464]},
     {otherUnit_maskInput_hi[20463:20448]},
     {otherUnit_maskInput_hi[20447:20432]},
     {otherUnit_maskInput_hi[20431:20416]},
     {otherUnit_maskInput_hi[20415:20400]},
     {otherUnit_maskInput_hi[20399:20384]},
     {otherUnit_maskInput_hi[20383:20368]},
     {otherUnit_maskInput_hi[20367:20352]},
     {otherUnit_maskInput_hi[20351:20336]},
     {otherUnit_maskInput_hi[20335:20320]},
     {otherUnit_maskInput_hi[20319:20304]},
     {otherUnit_maskInput_hi[20303:20288]},
     {otherUnit_maskInput_hi[20287:20272]},
     {otherUnit_maskInput_hi[20271:20256]},
     {otherUnit_maskInput_hi[20255:20240]},
     {otherUnit_maskInput_hi[20239:20224]},
     {otherUnit_maskInput_hi[20223:20208]},
     {otherUnit_maskInput_hi[20207:20192]},
     {otherUnit_maskInput_hi[20191:20176]},
     {otherUnit_maskInput_hi[20175:20160]},
     {otherUnit_maskInput_hi[20159:20144]},
     {otherUnit_maskInput_hi[20143:20128]},
     {otherUnit_maskInput_hi[20127:20112]},
     {otherUnit_maskInput_hi[20111:20096]},
     {otherUnit_maskInput_hi[20095:20080]},
     {otherUnit_maskInput_hi[20079:20064]},
     {otherUnit_maskInput_hi[20063:20048]},
     {otherUnit_maskInput_hi[20047:20032]},
     {otherUnit_maskInput_hi[20031:20016]},
     {otherUnit_maskInput_hi[20015:20000]},
     {otherUnit_maskInput_hi[19999:19984]},
     {otherUnit_maskInput_hi[19983:19968]},
     {otherUnit_maskInput_hi[19967:19952]},
     {otherUnit_maskInput_hi[19951:19936]},
     {otherUnit_maskInput_hi[19935:19920]},
     {otherUnit_maskInput_hi[19919:19904]},
     {otherUnit_maskInput_hi[19903:19888]},
     {otherUnit_maskInput_hi[19887:19872]},
     {otherUnit_maskInput_hi[19871:19856]},
     {otherUnit_maskInput_hi[19855:19840]},
     {otherUnit_maskInput_hi[19839:19824]},
     {otherUnit_maskInput_hi[19823:19808]},
     {otherUnit_maskInput_hi[19807:19792]},
     {otherUnit_maskInput_hi[19791:19776]},
     {otherUnit_maskInput_hi[19775:19760]},
     {otherUnit_maskInput_hi[19759:19744]},
     {otherUnit_maskInput_hi[19743:19728]},
     {otherUnit_maskInput_hi[19727:19712]},
     {otherUnit_maskInput_hi[19711:19696]},
     {otherUnit_maskInput_hi[19695:19680]},
     {otherUnit_maskInput_hi[19679:19664]},
     {otherUnit_maskInput_hi[19663:19648]},
     {otherUnit_maskInput_hi[19647:19632]},
     {otherUnit_maskInput_hi[19631:19616]},
     {otherUnit_maskInput_hi[19615:19600]},
     {otherUnit_maskInput_hi[19599:19584]},
     {otherUnit_maskInput_hi[19583:19568]},
     {otherUnit_maskInput_hi[19567:19552]},
     {otherUnit_maskInput_hi[19551:19536]},
     {otherUnit_maskInput_hi[19535:19520]},
     {otherUnit_maskInput_hi[19519:19504]},
     {otherUnit_maskInput_hi[19503:19488]},
     {otherUnit_maskInput_hi[19487:19472]},
     {otherUnit_maskInput_hi[19471:19456]},
     {otherUnit_maskInput_hi[19455:19440]},
     {otherUnit_maskInput_hi[19439:19424]},
     {otherUnit_maskInput_hi[19423:19408]},
     {otherUnit_maskInput_hi[19407:19392]},
     {otherUnit_maskInput_hi[19391:19376]},
     {otherUnit_maskInput_hi[19375:19360]},
     {otherUnit_maskInput_hi[19359:19344]},
     {otherUnit_maskInput_hi[19343:19328]},
     {otherUnit_maskInput_hi[19327:19312]},
     {otherUnit_maskInput_hi[19311:19296]},
     {otherUnit_maskInput_hi[19295:19280]},
     {otherUnit_maskInput_hi[19279:19264]},
     {otherUnit_maskInput_hi[19263:19248]},
     {otherUnit_maskInput_hi[19247:19232]},
     {otherUnit_maskInput_hi[19231:19216]},
     {otherUnit_maskInput_hi[19215:19200]},
     {otherUnit_maskInput_hi[19199:19184]},
     {otherUnit_maskInput_hi[19183:19168]},
     {otherUnit_maskInput_hi[19167:19152]},
     {otherUnit_maskInput_hi[19151:19136]},
     {otherUnit_maskInput_hi[19135:19120]},
     {otherUnit_maskInput_hi[19119:19104]},
     {otherUnit_maskInput_hi[19103:19088]},
     {otherUnit_maskInput_hi[19087:19072]},
     {otherUnit_maskInput_hi[19071:19056]},
     {otherUnit_maskInput_hi[19055:19040]},
     {otherUnit_maskInput_hi[19039:19024]},
     {otherUnit_maskInput_hi[19023:19008]},
     {otherUnit_maskInput_hi[19007:18992]},
     {otherUnit_maskInput_hi[18991:18976]},
     {otherUnit_maskInput_hi[18975:18960]},
     {otherUnit_maskInput_hi[18959:18944]},
     {otherUnit_maskInput_hi[18943:18928]},
     {otherUnit_maskInput_hi[18927:18912]},
     {otherUnit_maskInput_hi[18911:18896]},
     {otherUnit_maskInput_hi[18895:18880]},
     {otherUnit_maskInput_hi[18879:18864]},
     {otherUnit_maskInput_hi[18863:18848]},
     {otherUnit_maskInput_hi[18847:18832]},
     {otherUnit_maskInput_hi[18831:18816]},
     {otherUnit_maskInput_hi[18815:18800]},
     {otherUnit_maskInput_hi[18799:18784]},
     {otherUnit_maskInput_hi[18783:18768]},
     {otherUnit_maskInput_hi[18767:18752]},
     {otherUnit_maskInput_hi[18751:18736]},
     {otherUnit_maskInput_hi[18735:18720]},
     {otherUnit_maskInput_hi[18719:18704]},
     {otherUnit_maskInput_hi[18703:18688]},
     {otherUnit_maskInput_hi[18687:18672]},
     {otherUnit_maskInput_hi[18671:18656]},
     {otherUnit_maskInput_hi[18655:18640]},
     {otherUnit_maskInput_hi[18639:18624]},
     {otherUnit_maskInput_hi[18623:18608]},
     {otherUnit_maskInput_hi[18607:18592]},
     {otherUnit_maskInput_hi[18591:18576]},
     {otherUnit_maskInput_hi[18575:18560]},
     {otherUnit_maskInput_hi[18559:18544]},
     {otherUnit_maskInput_hi[18543:18528]},
     {otherUnit_maskInput_hi[18527:18512]},
     {otherUnit_maskInput_hi[18511:18496]},
     {otherUnit_maskInput_hi[18495:18480]},
     {otherUnit_maskInput_hi[18479:18464]},
     {otherUnit_maskInput_hi[18463:18448]},
     {otherUnit_maskInput_hi[18447:18432]},
     {otherUnit_maskInput_hi[18431:18416]},
     {otherUnit_maskInput_hi[18415:18400]},
     {otherUnit_maskInput_hi[18399:18384]},
     {otherUnit_maskInput_hi[18383:18368]},
     {otherUnit_maskInput_hi[18367:18352]},
     {otherUnit_maskInput_hi[18351:18336]},
     {otherUnit_maskInput_hi[18335:18320]},
     {otherUnit_maskInput_hi[18319:18304]},
     {otherUnit_maskInput_hi[18303:18288]},
     {otherUnit_maskInput_hi[18287:18272]},
     {otherUnit_maskInput_hi[18271:18256]},
     {otherUnit_maskInput_hi[18255:18240]},
     {otherUnit_maskInput_hi[18239:18224]},
     {otherUnit_maskInput_hi[18223:18208]},
     {otherUnit_maskInput_hi[18207:18192]},
     {otherUnit_maskInput_hi[18191:18176]},
     {otherUnit_maskInput_hi[18175:18160]},
     {otherUnit_maskInput_hi[18159:18144]},
     {otherUnit_maskInput_hi[18143:18128]},
     {otherUnit_maskInput_hi[18127:18112]},
     {otherUnit_maskInput_hi[18111:18096]},
     {otherUnit_maskInput_hi[18095:18080]},
     {otherUnit_maskInput_hi[18079:18064]},
     {otherUnit_maskInput_hi[18063:18048]},
     {otherUnit_maskInput_hi[18047:18032]},
     {otherUnit_maskInput_hi[18031:18016]},
     {otherUnit_maskInput_hi[18015:18000]},
     {otherUnit_maskInput_hi[17999:17984]},
     {otherUnit_maskInput_hi[17983:17968]},
     {otherUnit_maskInput_hi[17967:17952]},
     {otherUnit_maskInput_hi[17951:17936]},
     {otherUnit_maskInput_hi[17935:17920]},
     {otherUnit_maskInput_hi[17919:17904]},
     {otherUnit_maskInput_hi[17903:17888]},
     {otherUnit_maskInput_hi[17887:17872]},
     {otherUnit_maskInput_hi[17871:17856]},
     {otherUnit_maskInput_hi[17855:17840]},
     {otherUnit_maskInput_hi[17839:17824]},
     {otherUnit_maskInput_hi[17823:17808]},
     {otherUnit_maskInput_hi[17807:17792]},
     {otherUnit_maskInput_hi[17791:17776]},
     {otherUnit_maskInput_hi[17775:17760]},
     {otherUnit_maskInput_hi[17759:17744]},
     {otherUnit_maskInput_hi[17743:17728]},
     {otherUnit_maskInput_hi[17727:17712]},
     {otherUnit_maskInput_hi[17711:17696]},
     {otherUnit_maskInput_hi[17695:17680]},
     {otherUnit_maskInput_hi[17679:17664]},
     {otherUnit_maskInput_hi[17663:17648]},
     {otherUnit_maskInput_hi[17647:17632]},
     {otherUnit_maskInput_hi[17631:17616]},
     {otherUnit_maskInput_hi[17615:17600]},
     {otherUnit_maskInput_hi[17599:17584]},
     {otherUnit_maskInput_hi[17583:17568]},
     {otherUnit_maskInput_hi[17567:17552]},
     {otherUnit_maskInput_hi[17551:17536]},
     {otherUnit_maskInput_hi[17535:17520]},
     {otherUnit_maskInput_hi[17519:17504]},
     {otherUnit_maskInput_hi[17503:17488]},
     {otherUnit_maskInput_hi[17487:17472]},
     {otherUnit_maskInput_hi[17471:17456]},
     {otherUnit_maskInput_hi[17455:17440]},
     {otherUnit_maskInput_hi[17439:17424]},
     {otherUnit_maskInput_hi[17423:17408]},
     {otherUnit_maskInput_hi[17407:17392]},
     {otherUnit_maskInput_hi[17391:17376]},
     {otherUnit_maskInput_hi[17375:17360]},
     {otherUnit_maskInput_hi[17359:17344]},
     {otherUnit_maskInput_hi[17343:17328]},
     {otherUnit_maskInput_hi[17327:17312]},
     {otherUnit_maskInput_hi[17311:17296]},
     {otherUnit_maskInput_hi[17295:17280]},
     {otherUnit_maskInput_hi[17279:17264]},
     {otherUnit_maskInput_hi[17263:17248]},
     {otherUnit_maskInput_hi[17247:17232]},
     {otherUnit_maskInput_hi[17231:17216]},
     {otherUnit_maskInput_hi[17215:17200]},
     {otherUnit_maskInput_hi[17199:17184]},
     {otherUnit_maskInput_hi[17183:17168]},
     {otherUnit_maskInput_hi[17167:17152]},
     {otherUnit_maskInput_hi[17151:17136]},
     {otherUnit_maskInput_hi[17135:17120]},
     {otherUnit_maskInput_hi[17119:17104]},
     {otherUnit_maskInput_hi[17103:17088]},
     {otherUnit_maskInput_hi[17087:17072]},
     {otherUnit_maskInput_hi[17071:17056]},
     {otherUnit_maskInput_hi[17055:17040]},
     {otherUnit_maskInput_hi[17039:17024]},
     {otherUnit_maskInput_hi[17023:17008]},
     {otherUnit_maskInput_hi[17007:16992]},
     {otherUnit_maskInput_hi[16991:16976]},
     {otherUnit_maskInput_hi[16975:16960]},
     {otherUnit_maskInput_hi[16959:16944]},
     {otherUnit_maskInput_hi[16943:16928]},
     {otherUnit_maskInput_hi[16927:16912]},
     {otherUnit_maskInput_hi[16911:16896]},
     {otherUnit_maskInput_hi[16895:16880]},
     {otherUnit_maskInput_hi[16879:16864]},
     {otherUnit_maskInput_hi[16863:16848]},
     {otherUnit_maskInput_hi[16847:16832]},
     {otherUnit_maskInput_hi[16831:16816]},
     {otherUnit_maskInput_hi[16815:16800]},
     {otherUnit_maskInput_hi[16799:16784]},
     {otherUnit_maskInput_hi[16783:16768]},
     {otherUnit_maskInput_hi[16767:16752]},
     {otherUnit_maskInput_hi[16751:16736]},
     {otherUnit_maskInput_hi[16735:16720]},
     {otherUnit_maskInput_hi[16719:16704]},
     {otherUnit_maskInput_hi[16703:16688]},
     {otherUnit_maskInput_hi[16687:16672]},
     {otherUnit_maskInput_hi[16671:16656]},
     {otherUnit_maskInput_hi[16655:16640]},
     {otherUnit_maskInput_hi[16639:16624]},
     {otherUnit_maskInput_hi[16623:16608]},
     {otherUnit_maskInput_hi[16607:16592]},
     {otherUnit_maskInput_hi[16591:16576]},
     {otherUnit_maskInput_hi[16575:16560]},
     {otherUnit_maskInput_hi[16559:16544]},
     {otherUnit_maskInput_hi[16543:16528]},
     {otherUnit_maskInput_hi[16527:16512]},
     {otherUnit_maskInput_hi[16511:16496]},
     {otherUnit_maskInput_hi[16495:16480]},
     {otherUnit_maskInput_hi[16479:16464]},
     {otherUnit_maskInput_hi[16463:16448]},
     {otherUnit_maskInput_hi[16447:16432]},
     {otherUnit_maskInput_hi[16431:16416]},
     {otherUnit_maskInput_hi[16415:16400]},
     {otherUnit_maskInput_hi[16399:16384]},
     {otherUnit_maskInput_hi[16383:16368]},
     {otherUnit_maskInput_hi[16367:16352]},
     {otherUnit_maskInput_hi[16351:16336]},
     {otherUnit_maskInput_hi[16335:16320]},
     {otherUnit_maskInput_hi[16319:16304]},
     {otherUnit_maskInput_hi[16303:16288]},
     {otherUnit_maskInput_hi[16287:16272]},
     {otherUnit_maskInput_hi[16271:16256]},
     {otherUnit_maskInput_hi[16255:16240]},
     {otherUnit_maskInput_hi[16239:16224]},
     {otherUnit_maskInput_hi[16223:16208]},
     {otherUnit_maskInput_hi[16207:16192]},
     {otherUnit_maskInput_hi[16191:16176]},
     {otherUnit_maskInput_hi[16175:16160]},
     {otherUnit_maskInput_hi[16159:16144]},
     {otherUnit_maskInput_hi[16143:16128]},
     {otherUnit_maskInput_hi[16127:16112]},
     {otherUnit_maskInput_hi[16111:16096]},
     {otherUnit_maskInput_hi[16095:16080]},
     {otherUnit_maskInput_hi[16079:16064]},
     {otherUnit_maskInput_hi[16063:16048]},
     {otherUnit_maskInput_hi[16047:16032]},
     {otherUnit_maskInput_hi[16031:16016]},
     {otherUnit_maskInput_hi[16015:16000]},
     {otherUnit_maskInput_hi[15999:15984]},
     {otherUnit_maskInput_hi[15983:15968]},
     {otherUnit_maskInput_hi[15967:15952]},
     {otherUnit_maskInput_hi[15951:15936]},
     {otherUnit_maskInput_hi[15935:15920]},
     {otherUnit_maskInput_hi[15919:15904]},
     {otherUnit_maskInput_hi[15903:15888]},
     {otherUnit_maskInput_hi[15887:15872]},
     {otherUnit_maskInput_hi[15871:15856]},
     {otherUnit_maskInput_hi[15855:15840]},
     {otherUnit_maskInput_hi[15839:15824]},
     {otherUnit_maskInput_hi[15823:15808]},
     {otherUnit_maskInput_hi[15807:15792]},
     {otherUnit_maskInput_hi[15791:15776]},
     {otherUnit_maskInput_hi[15775:15760]},
     {otherUnit_maskInput_hi[15759:15744]},
     {otherUnit_maskInput_hi[15743:15728]},
     {otherUnit_maskInput_hi[15727:15712]},
     {otherUnit_maskInput_hi[15711:15696]},
     {otherUnit_maskInput_hi[15695:15680]},
     {otherUnit_maskInput_hi[15679:15664]},
     {otherUnit_maskInput_hi[15663:15648]},
     {otherUnit_maskInput_hi[15647:15632]},
     {otherUnit_maskInput_hi[15631:15616]},
     {otherUnit_maskInput_hi[15615:15600]},
     {otherUnit_maskInput_hi[15599:15584]},
     {otherUnit_maskInput_hi[15583:15568]},
     {otherUnit_maskInput_hi[15567:15552]},
     {otherUnit_maskInput_hi[15551:15536]},
     {otherUnit_maskInput_hi[15535:15520]},
     {otherUnit_maskInput_hi[15519:15504]},
     {otherUnit_maskInput_hi[15503:15488]},
     {otherUnit_maskInput_hi[15487:15472]},
     {otherUnit_maskInput_hi[15471:15456]},
     {otherUnit_maskInput_hi[15455:15440]},
     {otherUnit_maskInput_hi[15439:15424]},
     {otherUnit_maskInput_hi[15423:15408]},
     {otherUnit_maskInput_hi[15407:15392]},
     {otherUnit_maskInput_hi[15391:15376]},
     {otherUnit_maskInput_hi[15375:15360]},
     {otherUnit_maskInput_hi[15359:15344]},
     {otherUnit_maskInput_hi[15343:15328]},
     {otherUnit_maskInput_hi[15327:15312]},
     {otherUnit_maskInput_hi[15311:15296]},
     {otherUnit_maskInput_hi[15295:15280]},
     {otherUnit_maskInput_hi[15279:15264]},
     {otherUnit_maskInput_hi[15263:15248]},
     {otherUnit_maskInput_hi[15247:15232]},
     {otherUnit_maskInput_hi[15231:15216]},
     {otherUnit_maskInput_hi[15215:15200]},
     {otherUnit_maskInput_hi[15199:15184]},
     {otherUnit_maskInput_hi[15183:15168]},
     {otherUnit_maskInput_hi[15167:15152]},
     {otherUnit_maskInput_hi[15151:15136]},
     {otherUnit_maskInput_hi[15135:15120]},
     {otherUnit_maskInput_hi[15119:15104]},
     {otherUnit_maskInput_hi[15103:15088]},
     {otherUnit_maskInput_hi[15087:15072]},
     {otherUnit_maskInput_hi[15071:15056]},
     {otherUnit_maskInput_hi[15055:15040]},
     {otherUnit_maskInput_hi[15039:15024]},
     {otherUnit_maskInput_hi[15023:15008]},
     {otherUnit_maskInput_hi[15007:14992]},
     {otherUnit_maskInput_hi[14991:14976]},
     {otherUnit_maskInput_hi[14975:14960]},
     {otherUnit_maskInput_hi[14959:14944]},
     {otherUnit_maskInput_hi[14943:14928]},
     {otherUnit_maskInput_hi[14927:14912]},
     {otherUnit_maskInput_hi[14911:14896]},
     {otherUnit_maskInput_hi[14895:14880]},
     {otherUnit_maskInput_hi[14879:14864]},
     {otherUnit_maskInput_hi[14863:14848]},
     {otherUnit_maskInput_hi[14847:14832]},
     {otherUnit_maskInput_hi[14831:14816]},
     {otherUnit_maskInput_hi[14815:14800]},
     {otherUnit_maskInput_hi[14799:14784]},
     {otherUnit_maskInput_hi[14783:14768]},
     {otherUnit_maskInput_hi[14767:14752]},
     {otherUnit_maskInput_hi[14751:14736]},
     {otherUnit_maskInput_hi[14735:14720]},
     {otherUnit_maskInput_hi[14719:14704]},
     {otherUnit_maskInput_hi[14703:14688]},
     {otherUnit_maskInput_hi[14687:14672]},
     {otherUnit_maskInput_hi[14671:14656]},
     {otherUnit_maskInput_hi[14655:14640]},
     {otherUnit_maskInput_hi[14639:14624]},
     {otherUnit_maskInput_hi[14623:14608]},
     {otherUnit_maskInput_hi[14607:14592]},
     {otherUnit_maskInput_hi[14591:14576]},
     {otherUnit_maskInput_hi[14575:14560]},
     {otherUnit_maskInput_hi[14559:14544]},
     {otherUnit_maskInput_hi[14543:14528]},
     {otherUnit_maskInput_hi[14527:14512]},
     {otherUnit_maskInput_hi[14511:14496]},
     {otherUnit_maskInput_hi[14495:14480]},
     {otherUnit_maskInput_hi[14479:14464]},
     {otherUnit_maskInput_hi[14463:14448]},
     {otherUnit_maskInput_hi[14447:14432]},
     {otherUnit_maskInput_hi[14431:14416]},
     {otherUnit_maskInput_hi[14415:14400]},
     {otherUnit_maskInput_hi[14399:14384]},
     {otherUnit_maskInput_hi[14383:14368]},
     {otherUnit_maskInput_hi[14367:14352]},
     {otherUnit_maskInput_hi[14351:14336]},
     {otherUnit_maskInput_hi[14335:14320]},
     {otherUnit_maskInput_hi[14319:14304]},
     {otherUnit_maskInput_hi[14303:14288]},
     {otherUnit_maskInput_hi[14287:14272]},
     {otherUnit_maskInput_hi[14271:14256]},
     {otherUnit_maskInput_hi[14255:14240]},
     {otherUnit_maskInput_hi[14239:14224]},
     {otherUnit_maskInput_hi[14223:14208]},
     {otherUnit_maskInput_hi[14207:14192]},
     {otherUnit_maskInput_hi[14191:14176]},
     {otherUnit_maskInput_hi[14175:14160]},
     {otherUnit_maskInput_hi[14159:14144]},
     {otherUnit_maskInput_hi[14143:14128]},
     {otherUnit_maskInput_hi[14127:14112]},
     {otherUnit_maskInput_hi[14111:14096]},
     {otherUnit_maskInput_hi[14095:14080]},
     {otherUnit_maskInput_hi[14079:14064]},
     {otherUnit_maskInput_hi[14063:14048]},
     {otherUnit_maskInput_hi[14047:14032]},
     {otherUnit_maskInput_hi[14031:14016]},
     {otherUnit_maskInput_hi[14015:14000]},
     {otherUnit_maskInput_hi[13999:13984]},
     {otherUnit_maskInput_hi[13983:13968]},
     {otherUnit_maskInput_hi[13967:13952]},
     {otherUnit_maskInput_hi[13951:13936]},
     {otherUnit_maskInput_hi[13935:13920]},
     {otherUnit_maskInput_hi[13919:13904]},
     {otherUnit_maskInput_hi[13903:13888]},
     {otherUnit_maskInput_hi[13887:13872]},
     {otherUnit_maskInput_hi[13871:13856]},
     {otherUnit_maskInput_hi[13855:13840]},
     {otherUnit_maskInput_hi[13839:13824]},
     {otherUnit_maskInput_hi[13823:13808]},
     {otherUnit_maskInput_hi[13807:13792]},
     {otherUnit_maskInput_hi[13791:13776]},
     {otherUnit_maskInput_hi[13775:13760]},
     {otherUnit_maskInput_hi[13759:13744]},
     {otherUnit_maskInput_hi[13743:13728]},
     {otherUnit_maskInput_hi[13727:13712]},
     {otherUnit_maskInput_hi[13711:13696]},
     {otherUnit_maskInput_hi[13695:13680]},
     {otherUnit_maskInput_hi[13679:13664]},
     {otherUnit_maskInput_hi[13663:13648]},
     {otherUnit_maskInput_hi[13647:13632]},
     {otherUnit_maskInput_hi[13631:13616]},
     {otherUnit_maskInput_hi[13615:13600]},
     {otherUnit_maskInput_hi[13599:13584]},
     {otherUnit_maskInput_hi[13583:13568]},
     {otherUnit_maskInput_hi[13567:13552]},
     {otherUnit_maskInput_hi[13551:13536]},
     {otherUnit_maskInput_hi[13535:13520]},
     {otherUnit_maskInput_hi[13519:13504]},
     {otherUnit_maskInput_hi[13503:13488]},
     {otherUnit_maskInput_hi[13487:13472]},
     {otherUnit_maskInput_hi[13471:13456]},
     {otherUnit_maskInput_hi[13455:13440]},
     {otherUnit_maskInput_hi[13439:13424]},
     {otherUnit_maskInput_hi[13423:13408]},
     {otherUnit_maskInput_hi[13407:13392]},
     {otherUnit_maskInput_hi[13391:13376]},
     {otherUnit_maskInput_hi[13375:13360]},
     {otherUnit_maskInput_hi[13359:13344]},
     {otherUnit_maskInput_hi[13343:13328]},
     {otherUnit_maskInput_hi[13327:13312]},
     {otherUnit_maskInput_hi[13311:13296]},
     {otherUnit_maskInput_hi[13295:13280]},
     {otherUnit_maskInput_hi[13279:13264]},
     {otherUnit_maskInput_hi[13263:13248]},
     {otherUnit_maskInput_hi[13247:13232]},
     {otherUnit_maskInput_hi[13231:13216]},
     {otherUnit_maskInput_hi[13215:13200]},
     {otherUnit_maskInput_hi[13199:13184]},
     {otherUnit_maskInput_hi[13183:13168]},
     {otherUnit_maskInput_hi[13167:13152]},
     {otherUnit_maskInput_hi[13151:13136]},
     {otherUnit_maskInput_hi[13135:13120]},
     {otherUnit_maskInput_hi[13119:13104]},
     {otherUnit_maskInput_hi[13103:13088]},
     {otherUnit_maskInput_hi[13087:13072]},
     {otherUnit_maskInput_hi[13071:13056]},
     {otherUnit_maskInput_hi[13055:13040]},
     {otherUnit_maskInput_hi[13039:13024]},
     {otherUnit_maskInput_hi[13023:13008]},
     {otherUnit_maskInput_hi[13007:12992]},
     {otherUnit_maskInput_hi[12991:12976]},
     {otherUnit_maskInput_hi[12975:12960]},
     {otherUnit_maskInput_hi[12959:12944]},
     {otherUnit_maskInput_hi[12943:12928]},
     {otherUnit_maskInput_hi[12927:12912]},
     {otherUnit_maskInput_hi[12911:12896]},
     {otherUnit_maskInput_hi[12895:12880]},
     {otherUnit_maskInput_hi[12879:12864]},
     {otherUnit_maskInput_hi[12863:12848]},
     {otherUnit_maskInput_hi[12847:12832]},
     {otherUnit_maskInput_hi[12831:12816]},
     {otherUnit_maskInput_hi[12815:12800]},
     {otherUnit_maskInput_hi[12799:12784]},
     {otherUnit_maskInput_hi[12783:12768]},
     {otherUnit_maskInput_hi[12767:12752]},
     {otherUnit_maskInput_hi[12751:12736]},
     {otherUnit_maskInput_hi[12735:12720]},
     {otherUnit_maskInput_hi[12719:12704]},
     {otherUnit_maskInput_hi[12703:12688]},
     {otherUnit_maskInput_hi[12687:12672]},
     {otherUnit_maskInput_hi[12671:12656]},
     {otherUnit_maskInput_hi[12655:12640]},
     {otherUnit_maskInput_hi[12639:12624]},
     {otherUnit_maskInput_hi[12623:12608]},
     {otherUnit_maskInput_hi[12607:12592]},
     {otherUnit_maskInput_hi[12591:12576]},
     {otherUnit_maskInput_hi[12575:12560]},
     {otherUnit_maskInput_hi[12559:12544]},
     {otherUnit_maskInput_hi[12543:12528]},
     {otherUnit_maskInput_hi[12527:12512]},
     {otherUnit_maskInput_hi[12511:12496]},
     {otherUnit_maskInput_hi[12495:12480]},
     {otherUnit_maskInput_hi[12479:12464]},
     {otherUnit_maskInput_hi[12463:12448]},
     {otherUnit_maskInput_hi[12447:12432]},
     {otherUnit_maskInput_hi[12431:12416]},
     {otherUnit_maskInput_hi[12415:12400]},
     {otherUnit_maskInput_hi[12399:12384]},
     {otherUnit_maskInput_hi[12383:12368]},
     {otherUnit_maskInput_hi[12367:12352]},
     {otherUnit_maskInput_hi[12351:12336]},
     {otherUnit_maskInput_hi[12335:12320]},
     {otherUnit_maskInput_hi[12319:12304]},
     {otherUnit_maskInput_hi[12303:12288]},
     {otherUnit_maskInput_hi[12287:12272]},
     {otherUnit_maskInput_hi[12271:12256]},
     {otherUnit_maskInput_hi[12255:12240]},
     {otherUnit_maskInput_hi[12239:12224]},
     {otherUnit_maskInput_hi[12223:12208]},
     {otherUnit_maskInput_hi[12207:12192]},
     {otherUnit_maskInput_hi[12191:12176]},
     {otherUnit_maskInput_hi[12175:12160]},
     {otherUnit_maskInput_hi[12159:12144]},
     {otherUnit_maskInput_hi[12143:12128]},
     {otherUnit_maskInput_hi[12127:12112]},
     {otherUnit_maskInput_hi[12111:12096]},
     {otherUnit_maskInput_hi[12095:12080]},
     {otherUnit_maskInput_hi[12079:12064]},
     {otherUnit_maskInput_hi[12063:12048]},
     {otherUnit_maskInput_hi[12047:12032]},
     {otherUnit_maskInput_hi[12031:12016]},
     {otherUnit_maskInput_hi[12015:12000]},
     {otherUnit_maskInput_hi[11999:11984]},
     {otherUnit_maskInput_hi[11983:11968]},
     {otherUnit_maskInput_hi[11967:11952]},
     {otherUnit_maskInput_hi[11951:11936]},
     {otherUnit_maskInput_hi[11935:11920]},
     {otherUnit_maskInput_hi[11919:11904]},
     {otherUnit_maskInput_hi[11903:11888]},
     {otherUnit_maskInput_hi[11887:11872]},
     {otherUnit_maskInput_hi[11871:11856]},
     {otherUnit_maskInput_hi[11855:11840]},
     {otherUnit_maskInput_hi[11839:11824]},
     {otherUnit_maskInput_hi[11823:11808]},
     {otherUnit_maskInput_hi[11807:11792]},
     {otherUnit_maskInput_hi[11791:11776]},
     {otherUnit_maskInput_hi[11775:11760]},
     {otherUnit_maskInput_hi[11759:11744]},
     {otherUnit_maskInput_hi[11743:11728]},
     {otherUnit_maskInput_hi[11727:11712]},
     {otherUnit_maskInput_hi[11711:11696]},
     {otherUnit_maskInput_hi[11695:11680]},
     {otherUnit_maskInput_hi[11679:11664]},
     {otherUnit_maskInput_hi[11663:11648]},
     {otherUnit_maskInput_hi[11647:11632]},
     {otherUnit_maskInput_hi[11631:11616]},
     {otherUnit_maskInput_hi[11615:11600]},
     {otherUnit_maskInput_hi[11599:11584]},
     {otherUnit_maskInput_hi[11583:11568]},
     {otherUnit_maskInput_hi[11567:11552]},
     {otherUnit_maskInput_hi[11551:11536]},
     {otherUnit_maskInput_hi[11535:11520]},
     {otherUnit_maskInput_hi[11519:11504]},
     {otherUnit_maskInput_hi[11503:11488]},
     {otherUnit_maskInput_hi[11487:11472]},
     {otherUnit_maskInput_hi[11471:11456]},
     {otherUnit_maskInput_hi[11455:11440]},
     {otherUnit_maskInput_hi[11439:11424]},
     {otherUnit_maskInput_hi[11423:11408]},
     {otherUnit_maskInput_hi[11407:11392]},
     {otherUnit_maskInput_hi[11391:11376]},
     {otherUnit_maskInput_hi[11375:11360]},
     {otherUnit_maskInput_hi[11359:11344]},
     {otherUnit_maskInput_hi[11343:11328]},
     {otherUnit_maskInput_hi[11327:11312]},
     {otherUnit_maskInput_hi[11311:11296]},
     {otherUnit_maskInput_hi[11295:11280]},
     {otherUnit_maskInput_hi[11279:11264]},
     {otherUnit_maskInput_hi[11263:11248]},
     {otherUnit_maskInput_hi[11247:11232]},
     {otherUnit_maskInput_hi[11231:11216]},
     {otherUnit_maskInput_hi[11215:11200]},
     {otherUnit_maskInput_hi[11199:11184]},
     {otherUnit_maskInput_hi[11183:11168]},
     {otherUnit_maskInput_hi[11167:11152]},
     {otherUnit_maskInput_hi[11151:11136]},
     {otherUnit_maskInput_hi[11135:11120]},
     {otherUnit_maskInput_hi[11119:11104]},
     {otherUnit_maskInput_hi[11103:11088]},
     {otherUnit_maskInput_hi[11087:11072]},
     {otherUnit_maskInput_hi[11071:11056]},
     {otherUnit_maskInput_hi[11055:11040]},
     {otherUnit_maskInput_hi[11039:11024]},
     {otherUnit_maskInput_hi[11023:11008]},
     {otherUnit_maskInput_hi[11007:10992]},
     {otherUnit_maskInput_hi[10991:10976]},
     {otherUnit_maskInput_hi[10975:10960]},
     {otherUnit_maskInput_hi[10959:10944]},
     {otherUnit_maskInput_hi[10943:10928]},
     {otherUnit_maskInput_hi[10927:10912]},
     {otherUnit_maskInput_hi[10911:10896]},
     {otherUnit_maskInput_hi[10895:10880]},
     {otherUnit_maskInput_hi[10879:10864]},
     {otherUnit_maskInput_hi[10863:10848]},
     {otherUnit_maskInput_hi[10847:10832]},
     {otherUnit_maskInput_hi[10831:10816]},
     {otherUnit_maskInput_hi[10815:10800]},
     {otherUnit_maskInput_hi[10799:10784]},
     {otherUnit_maskInput_hi[10783:10768]},
     {otherUnit_maskInput_hi[10767:10752]},
     {otherUnit_maskInput_hi[10751:10736]},
     {otherUnit_maskInput_hi[10735:10720]},
     {otherUnit_maskInput_hi[10719:10704]},
     {otherUnit_maskInput_hi[10703:10688]},
     {otherUnit_maskInput_hi[10687:10672]},
     {otherUnit_maskInput_hi[10671:10656]},
     {otherUnit_maskInput_hi[10655:10640]},
     {otherUnit_maskInput_hi[10639:10624]},
     {otherUnit_maskInput_hi[10623:10608]},
     {otherUnit_maskInput_hi[10607:10592]},
     {otherUnit_maskInput_hi[10591:10576]},
     {otherUnit_maskInput_hi[10575:10560]},
     {otherUnit_maskInput_hi[10559:10544]},
     {otherUnit_maskInput_hi[10543:10528]},
     {otherUnit_maskInput_hi[10527:10512]},
     {otherUnit_maskInput_hi[10511:10496]},
     {otherUnit_maskInput_hi[10495:10480]},
     {otherUnit_maskInput_hi[10479:10464]},
     {otherUnit_maskInput_hi[10463:10448]},
     {otherUnit_maskInput_hi[10447:10432]},
     {otherUnit_maskInput_hi[10431:10416]},
     {otherUnit_maskInput_hi[10415:10400]},
     {otherUnit_maskInput_hi[10399:10384]},
     {otherUnit_maskInput_hi[10383:10368]},
     {otherUnit_maskInput_hi[10367:10352]},
     {otherUnit_maskInput_hi[10351:10336]},
     {otherUnit_maskInput_hi[10335:10320]},
     {otherUnit_maskInput_hi[10319:10304]},
     {otherUnit_maskInput_hi[10303:10288]},
     {otherUnit_maskInput_hi[10287:10272]},
     {otherUnit_maskInput_hi[10271:10256]},
     {otherUnit_maskInput_hi[10255:10240]},
     {otherUnit_maskInput_hi[10239:10224]},
     {otherUnit_maskInput_hi[10223:10208]},
     {otherUnit_maskInput_hi[10207:10192]},
     {otherUnit_maskInput_hi[10191:10176]},
     {otherUnit_maskInput_hi[10175:10160]},
     {otherUnit_maskInput_hi[10159:10144]},
     {otherUnit_maskInput_hi[10143:10128]},
     {otherUnit_maskInput_hi[10127:10112]},
     {otherUnit_maskInput_hi[10111:10096]},
     {otherUnit_maskInput_hi[10095:10080]},
     {otherUnit_maskInput_hi[10079:10064]},
     {otherUnit_maskInput_hi[10063:10048]},
     {otherUnit_maskInput_hi[10047:10032]},
     {otherUnit_maskInput_hi[10031:10016]},
     {otherUnit_maskInput_hi[10015:10000]},
     {otherUnit_maskInput_hi[9999:9984]},
     {otherUnit_maskInput_hi[9983:9968]},
     {otherUnit_maskInput_hi[9967:9952]},
     {otherUnit_maskInput_hi[9951:9936]},
     {otherUnit_maskInput_hi[9935:9920]},
     {otherUnit_maskInput_hi[9919:9904]},
     {otherUnit_maskInput_hi[9903:9888]},
     {otherUnit_maskInput_hi[9887:9872]},
     {otherUnit_maskInput_hi[9871:9856]},
     {otherUnit_maskInput_hi[9855:9840]},
     {otherUnit_maskInput_hi[9839:9824]},
     {otherUnit_maskInput_hi[9823:9808]},
     {otherUnit_maskInput_hi[9807:9792]},
     {otherUnit_maskInput_hi[9791:9776]},
     {otherUnit_maskInput_hi[9775:9760]},
     {otherUnit_maskInput_hi[9759:9744]},
     {otherUnit_maskInput_hi[9743:9728]},
     {otherUnit_maskInput_hi[9727:9712]},
     {otherUnit_maskInput_hi[9711:9696]},
     {otherUnit_maskInput_hi[9695:9680]},
     {otherUnit_maskInput_hi[9679:9664]},
     {otherUnit_maskInput_hi[9663:9648]},
     {otherUnit_maskInput_hi[9647:9632]},
     {otherUnit_maskInput_hi[9631:9616]},
     {otherUnit_maskInput_hi[9615:9600]},
     {otherUnit_maskInput_hi[9599:9584]},
     {otherUnit_maskInput_hi[9583:9568]},
     {otherUnit_maskInput_hi[9567:9552]},
     {otherUnit_maskInput_hi[9551:9536]},
     {otherUnit_maskInput_hi[9535:9520]},
     {otherUnit_maskInput_hi[9519:9504]},
     {otherUnit_maskInput_hi[9503:9488]},
     {otherUnit_maskInput_hi[9487:9472]},
     {otherUnit_maskInput_hi[9471:9456]},
     {otherUnit_maskInput_hi[9455:9440]},
     {otherUnit_maskInput_hi[9439:9424]},
     {otherUnit_maskInput_hi[9423:9408]},
     {otherUnit_maskInput_hi[9407:9392]},
     {otherUnit_maskInput_hi[9391:9376]},
     {otherUnit_maskInput_hi[9375:9360]},
     {otherUnit_maskInput_hi[9359:9344]},
     {otherUnit_maskInput_hi[9343:9328]},
     {otherUnit_maskInput_hi[9327:9312]},
     {otherUnit_maskInput_hi[9311:9296]},
     {otherUnit_maskInput_hi[9295:9280]},
     {otherUnit_maskInput_hi[9279:9264]},
     {otherUnit_maskInput_hi[9263:9248]},
     {otherUnit_maskInput_hi[9247:9232]},
     {otherUnit_maskInput_hi[9231:9216]},
     {otherUnit_maskInput_hi[9215:9200]},
     {otherUnit_maskInput_hi[9199:9184]},
     {otherUnit_maskInput_hi[9183:9168]},
     {otherUnit_maskInput_hi[9167:9152]},
     {otherUnit_maskInput_hi[9151:9136]},
     {otherUnit_maskInput_hi[9135:9120]},
     {otherUnit_maskInput_hi[9119:9104]},
     {otherUnit_maskInput_hi[9103:9088]},
     {otherUnit_maskInput_hi[9087:9072]},
     {otherUnit_maskInput_hi[9071:9056]},
     {otherUnit_maskInput_hi[9055:9040]},
     {otherUnit_maskInput_hi[9039:9024]},
     {otherUnit_maskInput_hi[9023:9008]},
     {otherUnit_maskInput_hi[9007:8992]},
     {otherUnit_maskInput_hi[8991:8976]},
     {otherUnit_maskInput_hi[8975:8960]},
     {otherUnit_maskInput_hi[8959:8944]},
     {otherUnit_maskInput_hi[8943:8928]},
     {otherUnit_maskInput_hi[8927:8912]},
     {otherUnit_maskInput_hi[8911:8896]},
     {otherUnit_maskInput_hi[8895:8880]},
     {otherUnit_maskInput_hi[8879:8864]},
     {otherUnit_maskInput_hi[8863:8848]},
     {otherUnit_maskInput_hi[8847:8832]},
     {otherUnit_maskInput_hi[8831:8816]},
     {otherUnit_maskInput_hi[8815:8800]},
     {otherUnit_maskInput_hi[8799:8784]},
     {otherUnit_maskInput_hi[8783:8768]},
     {otherUnit_maskInput_hi[8767:8752]},
     {otherUnit_maskInput_hi[8751:8736]},
     {otherUnit_maskInput_hi[8735:8720]},
     {otherUnit_maskInput_hi[8719:8704]},
     {otherUnit_maskInput_hi[8703:8688]},
     {otherUnit_maskInput_hi[8687:8672]},
     {otherUnit_maskInput_hi[8671:8656]},
     {otherUnit_maskInput_hi[8655:8640]},
     {otherUnit_maskInput_hi[8639:8624]},
     {otherUnit_maskInput_hi[8623:8608]},
     {otherUnit_maskInput_hi[8607:8592]},
     {otherUnit_maskInput_hi[8591:8576]},
     {otherUnit_maskInput_hi[8575:8560]},
     {otherUnit_maskInput_hi[8559:8544]},
     {otherUnit_maskInput_hi[8543:8528]},
     {otherUnit_maskInput_hi[8527:8512]},
     {otherUnit_maskInput_hi[8511:8496]},
     {otherUnit_maskInput_hi[8495:8480]},
     {otherUnit_maskInput_hi[8479:8464]},
     {otherUnit_maskInput_hi[8463:8448]},
     {otherUnit_maskInput_hi[8447:8432]},
     {otherUnit_maskInput_hi[8431:8416]},
     {otherUnit_maskInput_hi[8415:8400]},
     {otherUnit_maskInput_hi[8399:8384]},
     {otherUnit_maskInput_hi[8383:8368]},
     {otherUnit_maskInput_hi[8367:8352]},
     {otherUnit_maskInput_hi[8351:8336]},
     {otherUnit_maskInput_hi[8335:8320]},
     {otherUnit_maskInput_hi[8319:8304]},
     {otherUnit_maskInput_hi[8303:8288]},
     {otherUnit_maskInput_hi[8287:8272]},
     {otherUnit_maskInput_hi[8271:8256]},
     {otherUnit_maskInput_hi[8255:8240]},
     {otherUnit_maskInput_hi[8239:8224]},
     {otherUnit_maskInput_hi[8223:8208]},
     {otherUnit_maskInput_hi[8207:8192]},
     {otherUnit_maskInput_hi[8191:8176]},
     {otherUnit_maskInput_hi[8175:8160]},
     {otherUnit_maskInput_hi[8159:8144]},
     {otherUnit_maskInput_hi[8143:8128]},
     {otherUnit_maskInput_hi[8127:8112]},
     {otherUnit_maskInput_hi[8111:8096]},
     {otherUnit_maskInput_hi[8095:8080]},
     {otherUnit_maskInput_hi[8079:8064]},
     {otherUnit_maskInput_hi[8063:8048]},
     {otherUnit_maskInput_hi[8047:8032]},
     {otherUnit_maskInput_hi[8031:8016]},
     {otherUnit_maskInput_hi[8015:8000]},
     {otherUnit_maskInput_hi[7999:7984]},
     {otherUnit_maskInput_hi[7983:7968]},
     {otherUnit_maskInput_hi[7967:7952]},
     {otherUnit_maskInput_hi[7951:7936]},
     {otherUnit_maskInput_hi[7935:7920]},
     {otherUnit_maskInput_hi[7919:7904]},
     {otherUnit_maskInput_hi[7903:7888]},
     {otherUnit_maskInput_hi[7887:7872]},
     {otherUnit_maskInput_hi[7871:7856]},
     {otherUnit_maskInput_hi[7855:7840]},
     {otherUnit_maskInput_hi[7839:7824]},
     {otherUnit_maskInput_hi[7823:7808]},
     {otherUnit_maskInput_hi[7807:7792]},
     {otherUnit_maskInput_hi[7791:7776]},
     {otherUnit_maskInput_hi[7775:7760]},
     {otherUnit_maskInput_hi[7759:7744]},
     {otherUnit_maskInput_hi[7743:7728]},
     {otherUnit_maskInput_hi[7727:7712]},
     {otherUnit_maskInput_hi[7711:7696]},
     {otherUnit_maskInput_hi[7695:7680]},
     {otherUnit_maskInput_hi[7679:7664]},
     {otherUnit_maskInput_hi[7663:7648]},
     {otherUnit_maskInput_hi[7647:7632]},
     {otherUnit_maskInput_hi[7631:7616]},
     {otherUnit_maskInput_hi[7615:7600]},
     {otherUnit_maskInput_hi[7599:7584]},
     {otherUnit_maskInput_hi[7583:7568]},
     {otherUnit_maskInput_hi[7567:7552]},
     {otherUnit_maskInput_hi[7551:7536]},
     {otherUnit_maskInput_hi[7535:7520]},
     {otherUnit_maskInput_hi[7519:7504]},
     {otherUnit_maskInput_hi[7503:7488]},
     {otherUnit_maskInput_hi[7487:7472]},
     {otherUnit_maskInput_hi[7471:7456]},
     {otherUnit_maskInput_hi[7455:7440]},
     {otherUnit_maskInput_hi[7439:7424]},
     {otherUnit_maskInput_hi[7423:7408]},
     {otherUnit_maskInput_hi[7407:7392]},
     {otherUnit_maskInput_hi[7391:7376]},
     {otherUnit_maskInput_hi[7375:7360]},
     {otherUnit_maskInput_hi[7359:7344]},
     {otherUnit_maskInput_hi[7343:7328]},
     {otherUnit_maskInput_hi[7327:7312]},
     {otherUnit_maskInput_hi[7311:7296]},
     {otherUnit_maskInput_hi[7295:7280]},
     {otherUnit_maskInput_hi[7279:7264]},
     {otherUnit_maskInput_hi[7263:7248]},
     {otherUnit_maskInput_hi[7247:7232]},
     {otherUnit_maskInput_hi[7231:7216]},
     {otherUnit_maskInput_hi[7215:7200]},
     {otherUnit_maskInput_hi[7199:7184]},
     {otherUnit_maskInput_hi[7183:7168]},
     {otherUnit_maskInput_hi[7167:7152]},
     {otherUnit_maskInput_hi[7151:7136]},
     {otherUnit_maskInput_hi[7135:7120]},
     {otherUnit_maskInput_hi[7119:7104]},
     {otherUnit_maskInput_hi[7103:7088]},
     {otherUnit_maskInput_hi[7087:7072]},
     {otherUnit_maskInput_hi[7071:7056]},
     {otherUnit_maskInput_hi[7055:7040]},
     {otherUnit_maskInput_hi[7039:7024]},
     {otherUnit_maskInput_hi[7023:7008]},
     {otherUnit_maskInput_hi[7007:6992]},
     {otherUnit_maskInput_hi[6991:6976]},
     {otherUnit_maskInput_hi[6975:6960]},
     {otherUnit_maskInput_hi[6959:6944]},
     {otherUnit_maskInput_hi[6943:6928]},
     {otherUnit_maskInput_hi[6927:6912]},
     {otherUnit_maskInput_hi[6911:6896]},
     {otherUnit_maskInput_hi[6895:6880]},
     {otherUnit_maskInput_hi[6879:6864]},
     {otherUnit_maskInput_hi[6863:6848]},
     {otherUnit_maskInput_hi[6847:6832]},
     {otherUnit_maskInput_hi[6831:6816]},
     {otherUnit_maskInput_hi[6815:6800]},
     {otherUnit_maskInput_hi[6799:6784]},
     {otherUnit_maskInput_hi[6783:6768]},
     {otherUnit_maskInput_hi[6767:6752]},
     {otherUnit_maskInput_hi[6751:6736]},
     {otherUnit_maskInput_hi[6735:6720]},
     {otherUnit_maskInput_hi[6719:6704]},
     {otherUnit_maskInput_hi[6703:6688]},
     {otherUnit_maskInput_hi[6687:6672]},
     {otherUnit_maskInput_hi[6671:6656]},
     {otherUnit_maskInput_hi[6655:6640]},
     {otherUnit_maskInput_hi[6639:6624]},
     {otherUnit_maskInput_hi[6623:6608]},
     {otherUnit_maskInput_hi[6607:6592]},
     {otherUnit_maskInput_hi[6591:6576]},
     {otherUnit_maskInput_hi[6575:6560]},
     {otherUnit_maskInput_hi[6559:6544]},
     {otherUnit_maskInput_hi[6543:6528]},
     {otherUnit_maskInput_hi[6527:6512]},
     {otherUnit_maskInput_hi[6511:6496]},
     {otherUnit_maskInput_hi[6495:6480]},
     {otherUnit_maskInput_hi[6479:6464]},
     {otherUnit_maskInput_hi[6463:6448]},
     {otherUnit_maskInput_hi[6447:6432]},
     {otherUnit_maskInput_hi[6431:6416]},
     {otherUnit_maskInput_hi[6415:6400]},
     {otherUnit_maskInput_hi[6399:6384]},
     {otherUnit_maskInput_hi[6383:6368]},
     {otherUnit_maskInput_hi[6367:6352]},
     {otherUnit_maskInput_hi[6351:6336]},
     {otherUnit_maskInput_hi[6335:6320]},
     {otherUnit_maskInput_hi[6319:6304]},
     {otherUnit_maskInput_hi[6303:6288]},
     {otherUnit_maskInput_hi[6287:6272]},
     {otherUnit_maskInput_hi[6271:6256]},
     {otherUnit_maskInput_hi[6255:6240]},
     {otherUnit_maskInput_hi[6239:6224]},
     {otherUnit_maskInput_hi[6223:6208]},
     {otherUnit_maskInput_hi[6207:6192]},
     {otherUnit_maskInput_hi[6191:6176]},
     {otherUnit_maskInput_hi[6175:6160]},
     {otherUnit_maskInput_hi[6159:6144]},
     {otherUnit_maskInput_hi[6143:6128]},
     {otherUnit_maskInput_hi[6127:6112]},
     {otherUnit_maskInput_hi[6111:6096]},
     {otherUnit_maskInput_hi[6095:6080]},
     {otherUnit_maskInput_hi[6079:6064]},
     {otherUnit_maskInput_hi[6063:6048]},
     {otherUnit_maskInput_hi[6047:6032]},
     {otherUnit_maskInput_hi[6031:6016]},
     {otherUnit_maskInput_hi[6015:6000]},
     {otherUnit_maskInput_hi[5999:5984]},
     {otherUnit_maskInput_hi[5983:5968]},
     {otherUnit_maskInput_hi[5967:5952]},
     {otherUnit_maskInput_hi[5951:5936]},
     {otherUnit_maskInput_hi[5935:5920]},
     {otherUnit_maskInput_hi[5919:5904]},
     {otherUnit_maskInput_hi[5903:5888]},
     {otherUnit_maskInput_hi[5887:5872]},
     {otherUnit_maskInput_hi[5871:5856]},
     {otherUnit_maskInput_hi[5855:5840]},
     {otherUnit_maskInput_hi[5839:5824]},
     {otherUnit_maskInput_hi[5823:5808]},
     {otherUnit_maskInput_hi[5807:5792]},
     {otherUnit_maskInput_hi[5791:5776]},
     {otherUnit_maskInput_hi[5775:5760]},
     {otherUnit_maskInput_hi[5759:5744]},
     {otherUnit_maskInput_hi[5743:5728]},
     {otherUnit_maskInput_hi[5727:5712]},
     {otherUnit_maskInput_hi[5711:5696]},
     {otherUnit_maskInput_hi[5695:5680]},
     {otherUnit_maskInput_hi[5679:5664]},
     {otherUnit_maskInput_hi[5663:5648]},
     {otherUnit_maskInput_hi[5647:5632]},
     {otherUnit_maskInput_hi[5631:5616]},
     {otherUnit_maskInput_hi[5615:5600]},
     {otherUnit_maskInput_hi[5599:5584]},
     {otherUnit_maskInput_hi[5583:5568]},
     {otherUnit_maskInput_hi[5567:5552]},
     {otherUnit_maskInput_hi[5551:5536]},
     {otherUnit_maskInput_hi[5535:5520]},
     {otherUnit_maskInput_hi[5519:5504]},
     {otherUnit_maskInput_hi[5503:5488]},
     {otherUnit_maskInput_hi[5487:5472]},
     {otherUnit_maskInput_hi[5471:5456]},
     {otherUnit_maskInput_hi[5455:5440]},
     {otherUnit_maskInput_hi[5439:5424]},
     {otherUnit_maskInput_hi[5423:5408]},
     {otherUnit_maskInput_hi[5407:5392]},
     {otherUnit_maskInput_hi[5391:5376]},
     {otherUnit_maskInput_hi[5375:5360]},
     {otherUnit_maskInput_hi[5359:5344]},
     {otherUnit_maskInput_hi[5343:5328]},
     {otherUnit_maskInput_hi[5327:5312]},
     {otherUnit_maskInput_hi[5311:5296]},
     {otherUnit_maskInput_hi[5295:5280]},
     {otherUnit_maskInput_hi[5279:5264]},
     {otherUnit_maskInput_hi[5263:5248]},
     {otherUnit_maskInput_hi[5247:5232]},
     {otherUnit_maskInput_hi[5231:5216]},
     {otherUnit_maskInput_hi[5215:5200]},
     {otherUnit_maskInput_hi[5199:5184]},
     {otherUnit_maskInput_hi[5183:5168]},
     {otherUnit_maskInput_hi[5167:5152]},
     {otherUnit_maskInput_hi[5151:5136]},
     {otherUnit_maskInput_hi[5135:5120]},
     {otherUnit_maskInput_hi[5119:5104]},
     {otherUnit_maskInput_hi[5103:5088]},
     {otherUnit_maskInput_hi[5087:5072]},
     {otherUnit_maskInput_hi[5071:5056]},
     {otherUnit_maskInput_hi[5055:5040]},
     {otherUnit_maskInput_hi[5039:5024]},
     {otherUnit_maskInput_hi[5023:5008]},
     {otherUnit_maskInput_hi[5007:4992]},
     {otherUnit_maskInput_hi[4991:4976]},
     {otherUnit_maskInput_hi[4975:4960]},
     {otherUnit_maskInput_hi[4959:4944]},
     {otherUnit_maskInput_hi[4943:4928]},
     {otherUnit_maskInput_hi[4927:4912]},
     {otherUnit_maskInput_hi[4911:4896]},
     {otherUnit_maskInput_hi[4895:4880]},
     {otherUnit_maskInput_hi[4879:4864]},
     {otherUnit_maskInput_hi[4863:4848]},
     {otherUnit_maskInput_hi[4847:4832]},
     {otherUnit_maskInput_hi[4831:4816]},
     {otherUnit_maskInput_hi[4815:4800]},
     {otherUnit_maskInput_hi[4799:4784]},
     {otherUnit_maskInput_hi[4783:4768]},
     {otherUnit_maskInput_hi[4767:4752]},
     {otherUnit_maskInput_hi[4751:4736]},
     {otherUnit_maskInput_hi[4735:4720]},
     {otherUnit_maskInput_hi[4719:4704]},
     {otherUnit_maskInput_hi[4703:4688]},
     {otherUnit_maskInput_hi[4687:4672]},
     {otherUnit_maskInput_hi[4671:4656]},
     {otherUnit_maskInput_hi[4655:4640]},
     {otherUnit_maskInput_hi[4639:4624]},
     {otherUnit_maskInput_hi[4623:4608]},
     {otherUnit_maskInput_hi[4607:4592]},
     {otherUnit_maskInput_hi[4591:4576]},
     {otherUnit_maskInput_hi[4575:4560]},
     {otherUnit_maskInput_hi[4559:4544]},
     {otherUnit_maskInput_hi[4543:4528]},
     {otherUnit_maskInput_hi[4527:4512]},
     {otherUnit_maskInput_hi[4511:4496]},
     {otherUnit_maskInput_hi[4495:4480]},
     {otherUnit_maskInput_hi[4479:4464]},
     {otherUnit_maskInput_hi[4463:4448]},
     {otherUnit_maskInput_hi[4447:4432]},
     {otherUnit_maskInput_hi[4431:4416]},
     {otherUnit_maskInput_hi[4415:4400]},
     {otherUnit_maskInput_hi[4399:4384]},
     {otherUnit_maskInput_hi[4383:4368]},
     {otherUnit_maskInput_hi[4367:4352]},
     {otherUnit_maskInput_hi[4351:4336]},
     {otherUnit_maskInput_hi[4335:4320]},
     {otherUnit_maskInput_hi[4319:4304]},
     {otherUnit_maskInput_hi[4303:4288]},
     {otherUnit_maskInput_hi[4287:4272]},
     {otherUnit_maskInput_hi[4271:4256]},
     {otherUnit_maskInput_hi[4255:4240]},
     {otherUnit_maskInput_hi[4239:4224]},
     {otherUnit_maskInput_hi[4223:4208]},
     {otherUnit_maskInput_hi[4207:4192]},
     {otherUnit_maskInput_hi[4191:4176]},
     {otherUnit_maskInput_hi[4175:4160]},
     {otherUnit_maskInput_hi[4159:4144]},
     {otherUnit_maskInput_hi[4143:4128]},
     {otherUnit_maskInput_hi[4127:4112]},
     {otherUnit_maskInput_hi[4111:4096]},
     {otherUnit_maskInput_hi[4095:4080]},
     {otherUnit_maskInput_hi[4079:4064]},
     {otherUnit_maskInput_hi[4063:4048]},
     {otherUnit_maskInput_hi[4047:4032]},
     {otherUnit_maskInput_hi[4031:4016]},
     {otherUnit_maskInput_hi[4015:4000]},
     {otherUnit_maskInput_hi[3999:3984]},
     {otherUnit_maskInput_hi[3983:3968]},
     {otherUnit_maskInput_hi[3967:3952]},
     {otherUnit_maskInput_hi[3951:3936]},
     {otherUnit_maskInput_hi[3935:3920]},
     {otherUnit_maskInput_hi[3919:3904]},
     {otherUnit_maskInput_hi[3903:3888]},
     {otherUnit_maskInput_hi[3887:3872]},
     {otherUnit_maskInput_hi[3871:3856]},
     {otherUnit_maskInput_hi[3855:3840]},
     {otherUnit_maskInput_hi[3839:3824]},
     {otherUnit_maskInput_hi[3823:3808]},
     {otherUnit_maskInput_hi[3807:3792]},
     {otherUnit_maskInput_hi[3791:3776]},
     {otherUnit_maskInput_hi[3775:3760]},
     {otherUnit_maskInput_hi[3759:3744]},
     {otherUnit_maskInput_hi[3743:3728]},
     {otherUnit_maskInput_hi[3727:3712]},
     {otherUnit_maskInput_hi[3711:3696]},
     {otherUnit_maskInput_hi[3695:3680]},
     {otherUnit_maskInput_hi[3679:3664]},
     {otherUnit_maskInput_hi[3663:3648]},
     {otherUnit_maskInput_hi[3647:3632]},
     {otherUnit_maskInput_hi[3631:3616]},
     {otherUnit_maskInput_hi[3615:3600]},
     {otherUnit_maskInput_hi[3599:3584]},
     {otherUnit_maskInput_hi[3583:3568]},
     {otherUnit_maskInput_hi[3567:3552]},
     {otherUnit_maskInput_hi[3551:3536]},
     {otherUnit_maskInput_hi[3535:3520]},
     {otherUnit_maskInput_hi[3519:3504]},
     {otherUnit_maskInput_hi[3503:3488]},
     {otherUnit_maskInput_hi[3487:3472]},
     {otherUnit_maskInput_hi[3471:3456]},
     {otherUnit_maskInput_hi[3455:3440]},
     {otherUnit_maskInput_hi[3439:3424]},
     {otherUnit_maskInput_hi[3423:3408]},
     {otherUnit_maskInput_hi[3407:3392]},
     {otherUnit_maskInput_hi[3391:3376]},
     {otherUnit_maskInput_hi[3375:3360]},
     {otherUnit_maskInput_hi[3359:3344]},
     {otherUnit_maskInput_hi[3343:3328]},
     {otherUnit_maskInput_hi[3327:3312]},
     {otherUnit_maskInput_hi[3311:3296]},
     {otherUnit_maskInput_hi[3295:3280]},
     {otherUnit_maskInput_hi[3279:3264]},
     {otherUnit_maskInput_hi[3263:3248]},
     {otherUnit_maskInput_hi[3247:3232]},
     {otherUnit_maskInput_hi[3231:3216]},
     {otherUnit_maskInput_hi[3215:3200]},
     {otherUnit_maskInput_hi[3199:3184]},
     {otherUnit_maskInput_hi[3183:3168]},
     {otherUnit_maskInput_hi[3167:3152]},
     {otherUnit_maskInput_hi[3151:3136]},
     {otherUnit_maskInput_hi[3135:3120]},
     {otherUnit_maskInput_hi[3119:3104]},
     {otherUnit_maskInput_hi[3103:3088]},
     {otherUnit_maskInput_hi[3087:3072]},
     {otherUnit_maskInput_hi[3071:3056]},
     {otherUnit_maskInput_hi[3055:3040]},
     {otherUnit_maskInput_hi[3039:3024]},
     {otherUnit_maskInput_hi[3023:3008]},
     {otherUnit_maskInput_hi[3007:2992]},
     {otherUnit_maskInput_hi[2991:2976]},
     {otherUnit_maskInput_hi[2975:2960]},
     {otherUnit_maskInput_hi[2959:2944]},
     {otherUnit_maskInput_hi[2943:2928]},
     {otherUnit_maskInput_hi[2927:2912]},
     {otherUnit_maskInput_hi[2911:2896]},
     {otherUnit_maskInput_hi[2895:2880]},
     {otherUnit_maskInput_hi[2879:2864]},
     {otherUnit_maskInput_hi[2863:2848]},
     {otherUnit_maskInput_hi[2847:2832]},
     {otherUnit_maskInput_hi[2831:2816]},
     {otherUnit_maskInput_hi[2815:2800]},
     {otherUnit_maskInput_hi[2799:2784]},
     {otherUnit_maskInput_hi[2783:2768]},
     {otherUnit_maskInput_hi[2767:2752]},
     {otherUnit_maskInput_hi[2751:2736]},
     {otherUnit_maskInput_hi[2735:2720]},
     {otherUnit_maskInput_hi[2719:2704]},
     {otherUnit_maskInput_hi[2703:2688]},
     {otherUnit_maskInput_hi[2687:2672]},
     {otherUnit_maskInput_hi[2671:2656]},
     {otherUnit_maskInput_hi[2655:2640]},
     {otherUnit_maskInput_hi[2639:2624]},
     {otherUnit_maskInput_hi[2623:2608]},
     {otherUnit_maskInput_hi[2607:2592]},
     {otherUnit_maskInput_hi[2591:2576]},
     {otherUnit_maskInput_hi[2575:2560]},
     {otherUnit_maskInput_hi[2559:2544]},
     {otherUnit_maskInput_hi[2543:2528]},
     {otherUnit_maskInput_hi[2527:2512]},
     {otherUnit_maskInput_hi[2511:2496]},
     {otherUnit_maskInput_hi[2495:2480]},
     {otherUnit_maskInput_hi[2479:2464]},
     {otherUnit_maskInput_hi[2463:2448]},
     {otherUnit_maskInput_hi[2447:2432]},
     {otherUnit_maskInput_hi[2431:2416]},
     {otherUnit_maskInput_hi[2415:2400]},
     {otherUnit_maskInput_hi[2399:2384]},
     {otherUnit_maskInput_hi[2383:2368]},
     {otherUnit_maskInput_hi[2367:2352]},
     {otherUnit_maskInput_hi[2351:2336]},
     {otherUnit_maskInput_hi[2335:2320]},
     {otherUnit_maskInput_hi[2319:2304]},
     {otherUnit_maskInput_hi[2303:2288]},
     {otherUnit_maskInput_hi[2287:2272]},
     {otherUnit_maskInput_hi[2271:2256]},
     {otherUnit_maskInput_hi[2255:2240]},
     {otherUnit_maskInput_hi[2239:2224]},
     {otherUnit_maskInput_hi[2223:2208]},
     {otherUnit_maskInput_hi[2207:2192]},
     {otherUnit_maskInput_hi[2191:2176]},
     {otherUnit_maskInput_hi[2175:2160]},
     {otherUnit_maskInput_hi[2159:2144]},
     {otherUnit_maskInput_hi[2143:2128]},
     {otherUnit_maskInput_hi[2127:2112]},
     {otherUnit_maskInput_hi[2111:2096]},
     {otherUnit_maskInput_hi[2095:2080]},
     {otherUnit_maskInput_hi[2079:2064]},
     {otherUnit_maskInput_hi[2063:2048]},
     {otherUnit_maskInput_hi[2047:2032]},
     {otherUnit_maskInput_hi[2031:2016]},
     {otherUnit_maskInput_hi[2015:2000]},
     {otherUnit_maskInput_hi[1999:1984]},
     {otherUnit_maskInput_hi[1983:1968]},
     {otherUnit_maskInput_hi[1967:1952]},
     {otherUnit_maskInput_hi[1951:1936]},
     {otherUnit_maskInput_hi[1935:1920]},
     {otherUnit_maskInput_hi[1919:1904]},
     {otherUnit_maskInput_hi[1903:1888]},
     {otherUnit_maskInput_hi[1887:1872]},
     {otherUnit_maskInput_hi[1871:1856]},
     {otherUnit_maskInput_hi[1855:1840]},
     {otherUnit_maskInput_hi[1839:1824]},
     {otherUnit_maskInput_hi[1823:1808]},
     {otherUnit_maskInput_hi[1807:1792]},
     {otherUnit_maskInput_hi[1791:1776]},
     {otherUnit_maskInput_hi[1775:1760]},
     {otherUnit_maskInput_hi[1759:1744]},
     {otherUnit_maskInput_hi[1743:1728]},
     {otherUnit_maskInput_hi[1727:1712]},
     {otherUnit_maskInput_hi[1711:1696]},
     {otherUnit_maskInput_hi[1695:1680]},
     {otherUnit_maskInput_hi[1679:1664]},
     {otherUnit_maskInput_hi[1663:1648]},
     {otherUnit_maskInput_hi[1647:1632]},
     {otherUnit_maskInput_hi[1631:1616]},
     {otherUnit_maskInput_hi[1615:1600]},
     {otherUnit_maskInput_hi[1599:1584]},
     {otherUnit_maskInput_hi[1583:1568]},
     {otherUnit_maskInput_hi[1567:1552]},
     {otherUnit_maskInput_hi[1551:1536]},
     {otherUnit_maskInput_hi[1535:1520]},
     {otherUnit_maskInput_hi[1519:1504]},
     {otherUnit_maskInput_hi[1503:1488]},
     {otherUnit_maskInput_hi[1487:1472]},
     {otherUnit_maskInput_hi[1471:1456]},
     {otherUnit_maskInput_hi[1455:1440]},
     {otherUnit_maskInput_hi[1439:1424]},
     {otherUnit_maskInput_hi[1423:1408]},
     {otherUnit_maskInput_hi[1407:1392]},
     {otherUnit_maskInput_hi[1391:1376]},
     {otherUnit_maskInput_hi[1375:1360]},
     {otherUnit_maskInput_hi[1359:1344]},
     {otherUnit_maskInput_hi[1343:1328]},
     {otherUnit_maskInput_hi[1327:1312]},
     {otherUnit_maskInput_hi[1311:1296]},
     {otherUnit_maskInput_hi[1295:1280]},
     {otherUnit_maskInput_hi[1279:1264]},
     {otherUnit_maskInput_hi[1263:1248]},
     {otherUnit_maskInput_hi[1247:1232]},
     {otherUnit_maskInput_hi[1231:1216]},
     {otherUnit_maskInput_hi[1215:1200]},
     {otherUnit_maskInput_hi[1199:1184]},
     {otherUnit_maskInput_hi[1183:1168]},
     {otherUnit_maskInput_hi[1167:1152]},
     {otherUnit_maskInput_hi[1151:1136]},
     {otherUnit_maskInput_hi[1135:1120]},
     {otherUnit_maskInput_hi[1119:1104]},
     {otherUnit_maskInput_hi[1103:1088]},
     {otherUnit_maskInput_hi[1087:1072]},
     {otherUnit_maskInput_hi[1071:1056]},
     {otherUnit_maskInput_hi[1055:1040]},
     {otherUnit_maskInput_hi[1039:1024]},
     {otherUnit_maskInput_hi[1023:1008]},
     {otherUnit_maskInput_hi[1007:992]},
     {otherUnit_maskInput_hi[991:976]},
     {otherUnit_maskInput_hi[975:960]},
     {otherUnit_maskInput_hi[959:944]},
     {otherUnit_maskInput_hi[943:928]},
     {otherUnit_maskInput_hi[927:912]},
     {otherUnit_maskInput_hi[911:896]},
     {otherUnit_maskInput_hi[895:880]},
     {otherUnit_maskInput_hi[879:864]},
     {otherUnit_maskInput_hi[863:848]},
     {otherUnit_maskInput_hi[847:832]},
     {otherUnit_maskInput_hi[831:816]},
     {otherUnit_maskInput_hi[815:800]},
     {otherUnit_maskInput_hi[799:784]},
     {otherUnit_maskInput_hi[783:768]},
     {otherUnit_maskInput_hi[767:752]},
     {otherUnit_maskInput_hi[751:736]},
     {otherUnit_maskInput_hi[735:720]},
     {otherUnit_maskInput_hi[719:704]},
     {otherUnit_maskInput_hi[703:688]},
     {otherUnit_maskInput_hi[687:672]},
     {otherUnit_maskInput_hi[671:656]},
     {otherUnit_maskInput_hi[655:640]},
     {otherUnit_maskInput_hi[639:624]},
     {otherUnit_maskInput_hi[623:608]},
     {otherUnit_maskInput_hi[607:592]},
     {otherUnit_maskInput_hi[591:576]},
     {otherUnit_maskInput_hi[575:560]},
     {otherUnit_maskInput_hi[559:544]},
     {otherUnit_maskInput_hi[543:528]},
     {otherUnit_maskInput_hi[527:512]},
     {otherUnit_maskInput_hi[511:496]},
     {otherUnit_maskInput_hi[495:480]},
     {otherUnit_maskInput_hi[479:464]},
     {otherUnit_maskInput_hi[463:448]},
     {otherUnit_maskInput_hi[447:432]},
     {otherUnit_maskInput_hi[431:416]},
     {otherUnit_maskInput_hi[415:400]},
     {otherUnit_maskInput_hi[399:384]},
     {otherUnit_maskInput_hi[383:368]},
     {otherUnit_maskInput_hi[367:352]},
     {otherUnit_maskInput_hi[351:336]},
     {otherUnit_maskInput_hi[335:320]},
     {otherUnit_maskInput_hi[319:304]},
     {otherUnit_maskInput_hi[303:288]},
     {otherUnit_maskInput_hi[287:272]},
     {otherUnit_maskInput_hi[271:256]},
     {otherUnit_maskInput_hi[255:240]},
     {otherUnit_maskInput_hi[239:224]},
     {otherUnit_maskInput_hi[223:208]},
     {otherUnit_maskInput_hi[207:192]},
     {otherUnit_maskInput_hi[191:176]},
     {otherUnit_maskInput_hi[175:160]},
     {otherUnit_maskInput_hi[159:144]},
     {otherUnit_maskInput_hi[143:128]},
     {otherUnit_maskInput_hi[127:112]},
     {otherUnit_maskInput_hi[111:96]},
     {otherUnit_maskInput_hi[95:80]},
     {otherUnit_maskInput_hi[79:64]},
     {otherUnit_maskInput_hi[63:48]},
     {otherUnit_maskInput_hi[47:32]},
     {otherUnit_maskInput_hi[31:16]},
     {otherUnit_maskInput_hi[15:0]},
     {otherUnit_maskInput_lo[32767:32752]},
     {otherUnit_maskInput_lo[32751:32736]},
     {otherUnit_maskInput_lo[32735:32720]},
     {otherUnit_maskInput_lo[32719:32704]},
     {otherUnit_maskInput_lo[32703:32688]},
     {otherUnit_maskInput_lo[32687:32672]},
     {otherUnit_maskInput_lo[32671:32656]},
     {otherUnit_maskInput_lo[32655:32640]},
     {otherUnit_maskInput_lo[32639:32624]},
     {otherUnit_maskInput_lo[32623:32608]},
     {otherUnit_maskInput_lo[32607:32592]},
     {otherUnit_maskInput_lo[32591:32576]},
     {otherUnit_maskInput_lo[32575:32560]},
     {otherUnit_maskInput_lo[32559:32544]},
     {otherUnit_maskInput_lo[32543:32528]},
     {otherUnit_maskInput_lo[32527:32512]},
     {otherUnit_maskInput_lo[32511:32496]},
     {otherUnit_maskInput_lo[32495:32480]},
     {otherUnit_maskInput_lo[32479:32464]},
     {otherUnit_maskInput_lo[32463:32448]},
     {otherUnit_maskInput_lo[32447:32432]},
     {otherUnit_maskInput_lo[32431:32416]},
     {otherUnit_maskInput_lo[32415:32400]},
     {otherUnit_maskInput_lo[32399:32384]},
     {otherUnit_maskInput_lo[32383:32368]},
     {otherUnit_maskInput_lo[32367:32352]},
     {otherUnit_maskInput_lo[32351:32336]},
     {otherUnit_maskInput_lo[32335:32320]},
     {otherUnit_maskInput_lo[32319:32304]},
     {otherUnit_maskInput_lo[32303:32288]},
     {otherUnit_maskInput_lo[32287:32272]},
     {otherUnit_maskInput_lo[32271:32256]},
     {otherUnit_maskInput_lo[32255:32240]},
     {otherUnit_maskInput_lo[32239:32224]},
     {otherUnit_maskInput_lo[32223:32208]},
     {otherUnit_maskInput_lo[32207:32192]},
     {otherUnit_maskInput_lo[32191:32176]},
     {otherUnit_maskInput_lo[32175:32160]},
     {otherUnit_maskInput_lo[32159:32144]},
     {otherUnit_maskInput_lo[32143:32128]},
     {otherUnit_maskInput_lo[32127:32112]},
     {otherUnit_maskInput_lo[32111:32096]},
     {otherUnit_maskInput_lo[32095:32080]},
     {otherUnit_maskInput_lo[32079:32064]},
     {otherUnit_maskInput_lo[32063:32048]},
     {otherUnit_maskInput_lo[32047:32032]},
     {otherUnit_maskInput_lo[32031:32016]},
     {otherUnit_maskInput_lo[32015:32000]},
     {otherUnit_maskInput_lo[31999:31984]},
     {otherUnit_maskInput_lo[31983:31968]},
     {otherUnit_maskInput_lo[31967:31952]},
     {otherUnit_maskInput_lo[31951:31936]},
     {otherUnit_maskInput_lo[31935:31920]},
     {otherUnit_maskInput_lo[31919:31904]},
     {otherUnit_maskInput_lo[31903:31888]},
     {otherUnit_maskInput_lo[31887:31872]},
     {otherUnit_maskInput_lo[31871:31856]},
     {otherUnit_maskInput_lo[31855:31840]},
     {otherUnit_maskInput_lo[31839:31824]},
     {otherUnit_maskInput_lo[31823:31808]},
     {otherUnit_maskInput_lo[31807:31792]},
     {otherUnit_maskInput_lo[31791:31776]},
     {otherUnit_maskInput_lo[31775:31760]},
     {otherUnit_maskInput_lo[31759:31744]},
     {otherUnit_maskInput_lo[31743:31728]},
     {otherUnit_maskInput_lo[31727:31712]},
     {otherUnit_maskInput_lo[31711:31696]},
     {otherUnit_maskInput_lo[31695:31680]},
     {otherUnit_maskInput_lo[31679:31664]},
     {otherUnit_maskInput_lo[31663:31648]},
     {otherUnit_maskInput_lo[31647:31632]},
     {otherUnit_maskInput_lo[31631:31616]},
     {otherUnit_maskInput_lo[31615:31600]},
     {otherUnit_maskInput_lo[31599:31584]},
     {otherUnit_maskInput_lo[31583:31568]},
     {otherUnit_maskInput_lo[31567:31552]},
     {otherUnit_maskInput_lo[31551:31536]},
     {otherUnit_maskInput_lo[31535:31520]},
     {otherUnit_maskInput_lo[31519:31504]},
     {otherUnit_maskInput_lo[31503:31488]},
     {otherUnit_maskInput_lo[31487:31472]},
     {otherUnit_maskInput_lo[31471:31456]},
     {otherUnit_maskInput_lo[31455:31440]},
     {otherUnit_maskInput_lo[31439:31424]},
     {otherUnit_maskInput_lo[31423:31408]},
     {otherUnit_maskInput_lo[31407:31392]},
     {otherUnit_maskInput_lo[31391:31376]},
     {otherUnit_maskInput_lo[31375:31360]},
     {otherUnit_maskInput_lo[31359:31344]},
     {otherUnit_maskInput_lo[31343:31328]},
     {otherUnit_maskInput_lo[31327:31312]},
     {otherUnit_maskInput_lo[31311:31296]},
     {otherUnit_maskInput_lo[31295:31280]},
     {otherUnit_maskInput_lo[31279:31264]},
     {otherUnit_maskInput_lo[31263:31248]},
     {otherUnit_maskInput_lo[31247:31232]},
     {otherUnit_maskInput_lo[31231:31216]},
     {otherUnit_maskInput_lo[31215:31200]},
     {otherUnit_maskInput_lo[31199:31184]},
     {otherUnit_maskInput_lo[31183:31168]},
     {otherUnit_maskInput_lo[31167:31152]},
     {otherUnit_maskInput_lo[31151:31136]},
     {otherUnit_maskInput_lo[31135:31120]},
     {otherUnit_maskInput_lo[31119:31104]},
     {otherUnit_maskInput_lo[31103:31088]},
     {otherUnit_maskInput_lo[31087:31072]},
     {otherUnit_maskInput_lo[31071:31056]},
     {otherUnit_maskInput_lo[31055:31040]},
     {otherUnit_maskInput_lo[31039:31024]},
     {otherUnit_maskInput_lo[31023:31008]},
     {otherUnit_maskInput_lo[31007:30992]},
     {otherUnit_maskInput_lo[30991:30976]},
     {otherUnit_maskInput_lo[30975:30960]},
     {otherUnit_maskInput_lo[30959:30944]},
     {otherUnit_maskInput_lo[30943:30928]},
     {otherUnit_maskInput_lo[30927:30912]},
     {otherUnit_maskInput_lo[30911:30896]},
     {otherUnit_maskInput_lo[30895:30880]},
     {otherUnit_maskInput_lo[30879:30864]},
     {otherUnit_maskInput_lo[30863:30848]},
     {otherUnit_maskInput_lo[30847:30832]},
     {otherUnit_maskInput_lo[30831:30816]},
     {otherUnit_maskInput_lo[30815:30800]},
     {otherUnit_maskInput_lo[30799:30784]},
     {otherUnit_maskInput_lo[30783:30768]},
     {otherUnit_maskInput_lo[30767:30752]},
     {otherUnit_maskInput_lo[30751:30736]},
     {otherUnit_maskInput_lo[30735:30720]},
     {otherUnit_maskInput_lo[30719:30704]},
     {otherUnit_maskInput_lo[30703:30688]},
     {otherUnit_maskInput_lo[30687:30672]},
     {otherUnit_maskInput_lo[30671:30656]},
     {otherUnit_maskInput_lo[30655:30640]},
     {otherUnit_maskInput_lo[30639:30624]},
     {otherUnit_maskInput_lo[30623:30608]},
     {otherUnit_maskInput_lo[30607:30592]},
     {otherUnit_maskInput_lo[30591:30576]},
     {otherUnit_maskInput_lo[30575:30560]},
     {otherUnit_maskInput_lo[30559:30544]},
     {otherUnit_maskInput_lo[30543:30528]},
     {otherUnit_maskInput_lo[30527:30512]},
     {otherUnit_maskInput_lo[30511:30496]},
     {otherUnit_maskInput_lo[30495:30480]},
     {otherUnit_maskInput_lo[30479:30464]},
     {otherUnit_maskInput_lo[30463:30448]},
     {otherUnit_maskInput_lo[30447:30432]},
     {otherUnit_maskInput_lo[30431:30416]},
     {otherUnit_maskInput_lo[30415:30400]},
     {otherUnit_maskInput_lo[30399:30384]},
     {otherUnit_maskInput_lo[30383:30368]},
     {otherUnit_maskInput_lo[30367:30352]},
     {otherUnit_maskInput_lo[30351:30336]},
     {otherUnit_maskInput_lo[30335:30320]},
     {otherUnit_maskInput_lo[30319:30304]},
     {otherUnit_maskInput_lo[30303:30288]},
     {otherUnit_maskInput_lo[30287:30272]},
     {otherUnit_maskInput_lo[30271:30256]},
     {otherUnit_maskInput_lo[30255:30240]},
     {otherUnit_maskInput_lo[30239:30224]},
     {otherUnit_maskInput_lo[30223:30208]},
     {otherUnit_maskInput_lo[30207:30192]},
     {otherUnit_maskInput_lo[30191:30176]},
     {otherUnit_maskInput_lo[30175:30160]},
     {otherUnit_maskInput_lo[30159:30144]},
     {otherUnit_maskInput_lo[30143:30128]},
     {otherUnit_maskInput_lo[30127:30112]},
     {otherUnit_maskInput_lo[30111:30096]},
     {otherUnit_maskInput_lo[30095:30080]},
     {otherUnit_maskInput_lo[30079:30064]},
     {otherUnit_maskInput_lo[30063:30048]},
     {otherUnit_maskInput_lo[30047:30032]},
     {otherUnit_maskInput_lo[30031:30016]},
     {otherUnit_maskInput_lo[30015:30000]},
     {otherUnit_maskInput_lo[29999:29984]},
     {otherUnit_maskInput_lo[29983:29968]},
     {otherUnit_maskInput_lo[29967:29952]},
     {otherUnit_maskInput_lo[29951:29936]},
     {otherUnit_maskInput_lo[29935:29920]},
     {otherUnit_maskInput_lo[29919:29904]},
     {otherUnit_maskInput_lo[29903:29888]},
     {otherUnit_maskInput_lo[29887:29872]},
     {otherUnit_maskInput_lo[29871:29856]},
     {otherUnit_maskInput_lo[29855:29840]},
     {otherUnit_maskInput_lo[29839:29824]},
     {otherUnit_maskInput_lo[29823:29808]},
     {otherUnit_maskInput_lo[29807:29792]},
     {otherUnit_maskInput_lo[29791:29776]},
     {otherUnit_maskInput_lo[29775:29760]},
     {otherUnit_maskInput_lo[29759:29744]},
     {otherUnit_maskInput_lo[29743:29728]},
     {otherUnit_maskInput_lo[29727:29712]},
     {otherUnit_maskInput_lo[29711:29696]},
     {otherUnit_maskInput_lo[29695:29680]},
     {otherUnit_maskInput_lo[29679:29664]},
     {otherUnit_maskInput_lo[29663:29648]},
     {otherUnit_maskInput_lo[29647:29632]},
     {otherUnit_maskInput_lo[29631:29616]},
     {otherUnit_maskInput_lo[29615:29600]},
     {otherUnit_maskInput_lo[29599:29584]},
     {otherUnit_maskInput_lo[29583:29568]},
     {otherUnit_maskInput_lo[29567:29552]},
     {otherUnit_maskInput_lo[29551:29536]},
     {otherUnit_maskInput_lo[29535:29520]},
     {otherUnit_maskInput_lo[29519:29504]},
     {otherUnit_maskInput_lo[29503:29488]},
     {otherUnit_maskInput_lo[29487:29472]},
     {otherUnit_maskInput_lo[29471:29456]},
     {otherUnit_maskInput_lo[29455:29440]},
     {otherUnit_maskInput_lo[29439:29424]},
     {otherUnit_maskInput_lo[29423:29408]},
     {otherUnit_maskInput_lo[29407:29392]},
     {otherUnit_maskInput_lo[29391:29376]},
     {otherUnit_maskInput_lo[29375:29360]},
     {otherUnit_maskInput_lo[29359:29344]},
     {otherUnit_maskInput_lo[29343:29328]},
     {otherUnit_maskInput_lo[29327:29312]},
     {otherUnit_maskInput_lo[29311:29296]},
     {otherUnit_maskInput_lo[29295:29280]},
     {otherUnit_maskInput_lo[29279:29264]},
     {otherUnit_maskInput_lo[29263:29248]},
     {otherUnit_maskInput_lo[29247:29232]},
     {otherUnit_maskInput_lo[29231:29216]},
     {otherUnit_maskInput_lo[29215:29200]},
     {otherUnit_maskInput_lo[29199:29184]},
     {otherUnit_maskInput_lo[29183:29168]},
     {otherUnit_maskInput_lo[29167:29152]},
     {otherUnit_maskInput_lo[29151:29136]},
     {otherUnit_maskInput_lo[29135:29120]},
     {otherUnit_maskInput_lo[29119:29104]},
     {otherUnit_maskInput_lo[29103:29088]},
     {otherUnit_maskInput_lo[29087:29072]},
     {otherUnit_maskInput_lo[29071:29056]},
     {otherUnit_maskInput_lo[29055:29040]},
     {otherUnit_maskInput_lo[29039:29024]},
     {otherUnit_maskInput_lo[29023:29008]},
     {otherUnit_maskInput_lo[29007:28992]},
     {otherUnit_maskInput_lo[28991:28976]},
     {otherUnit_maskInput_lo[28975:28960]},
     {otherUnit_maskInput_lo[28959:28944]},
     {otherUnit_maskInput_lo[28943:28928]},
     {otherUnit_maskInput_lo[28927:28912]},
     {otherUnit_maskInput_lo[28911:28896]},
     {otherUnit_maskInput_lo[28895:28880]},
     {otherUnit_maskInput_lo[28879:28864]},
     {otherUnit_maskInput_lo[28863:28848]},
     {otherUnit_maskInput_lo[28847:28832]},
     {otherUnit_maskInput_lo[28831:28816]},
     {otherUnit_maskInput_lo[28815:28800]},
     {otherUnit_maskInput_lo[28799:28784]},
     {otherUnit_maskInput_lo[28783:28768]},
     {otherUnit_maskInput_lo[28767:28752]},
     {otherUnit_maskInput_lo[28751:28736]},
     {otherUnit_maskInput_lo[28735:28720]},
     {otherUnit_maskInput_lo[28719:28704]},
     {otherUnit_maskInput_lo[28703:28688]},
     {otherUnit_maskInput_lo[28687:28672]},
     {otherUnit_maskInput_lo[28671:28656]},
     {otherUnit_maskInput_lo[28655:28640]},
     {otherUnit_maskInput_lo[28639:28624]},
     {otherUnit_maskInput_lo[28623:28608]},
     {otherUnit_maskInput_lo[28607:28592]},
     {otherUnit_maskInput_lo[28591:28576]},
     {otherUnit_maskInput_lo[28575:28560]},
     {otherUnit_maskInput_lo[28559:28544]},
     {otherUnit_maskInput_lo[28543:28528]},
     {otherUnit_maskInput_lo[28527:28512]},
     {otherUnit_maskInput_lo[28511:28496]},
     {otherUnit_maskInput_lo[28495:28480]},
     {otherUnit_maskInput_lo[28479:28464]},
     {otherUnit_maskInput_lo[28463:28448]},
     {otherUnit_maskInput_lo[28447:28432]},
     {otherUnit_maskInput_lo[28431:28416]},
     {otherUnit_maskInput_lo[28415:28400]},
     {otherUnit_maskInput_lo[28399:28384]},
     {otherUnit_maskInput_lo[28383:28368]},
     {otherUnit_maskInput_lo[28367:28352]},
     {otherUnit_maskInput_lo[28351:28336]},
     {otherUnit_maskInput_lo[28335:28320]},
     {otherUnit_maskInput_lo[28319:28304]},
     {otherUnit_maskInput_lo[28303:28288]},
     {otherUnit_maskInput_lo[28287:28272]},
     {otherUnit_maskInput_lo[28271:28256]},
     {otherUnit_maskInput_lo[28255:28240]},
     {otherUnit_maskInput_lo[28239:28224]},
     {otherUnit_maskInput_lo[28223:28208]},
     {otherUnit_maskInput_lo[28207:28192]},
     {otherUnit_maskInput_lo[28191:28176]},
     {otherUnit_maskInput_lo[28175:28160]},
     {otherUnit_maskInput_lo[28159:28144]},
     {otherUnit_maskInput_lo[28143:28128]},
     {otherUnit_maskInput_lo[28127:28112]},
     {otherUnit_maskInput_lo[28111:28096]},
     {otherUnit_maskInput_lo[28095:28080]},
     {otherUnit_maskInput_lo[28079:28064]},
     {otherUnit_maskInput_lo[28063:28048]},
     {otherUnit_maskInput_lo[28047:28032]},
     {otherUnit_maskInput_lo[28031:28016]},
     {otherUnit_maskInput_lo[28015:28000]},
     {otherUnit_maskInput_lo[27999:27984]},
     {otherUnit_maskInput_lo[27983:27968]},
     {otherUnit_maskInput_lo[27967:27952]},
     {otherUnit_maskInput_lo[27951:27936]},
     {otherUnit_maskInput_lo[27935:27920]},
     {otherUnit_maskInput_lo[27919:27904]},
     {otherUnit_maskInput_lo[27903:27888]},
     {otherUnit_maskInput_lo[27887:27872]},
     {otherUnit_maskInput_lo[27871:27856]},
     {otherUnit_maskInput_lo[27855:27840]},
     {otherUnit_maskInput_lo[27839:27824]},
     {otherUnit_maskInput_lo[27823:27808]},
     {otherUnit_maskInput_lo[27807:27792]},
     {otherUnit_maskInput_lo[27791:27776]},
     {otherUnit_maskInput_lo[27775:27760]},
     {otherUnit_maskInput_lo[27759:27744]},
     {otherUnit_maskInput_lo[27743:27728]},
     {otherUnit_maskInput_lo[27727:27712]},
     {otherUnit_maskInput_lo[27711:27696]},
     {otherUnit_maskInput_lo[27695:27680]},
     {otherUnit_maskInput_lo[27679:27664]},
     {otherUnit_maskInput_lo[27663:27648]},
     {otherUnit_maskInput_lo[27647:27632]},
     {otherUnit_maskInput_lo[27631:27616]},
     {otherUnit_maskInput_lo[27615:27600]},
     {otherUnit_maskInput_lo[27599:27584]},
     {otherUnit_maskInput_lo[27583:27568]},
     {otherUnit_maskInput_lo[27567:27552]},
     {otherUnit_maskInput_lo[27551:27536]},
     {otherUnit_maskInput_lo[27535:27520]},
     {otherUnit_maskInput_lo[27519:27504]},
     {otherUnit_maskInput_lo[27503:27488]},
     {otherUnit_maskInput_lo[27487:27472]},
     {otherUnit_maskInput_lo[27471:27456]},
     {otherUnit_maskInput_lo[27455:27440]},
     {otherUnit_maskInput_lo[27439:27424]},
     {otherUnit_maskInput_lo[27423:27408]},
     {otherUnit_maskInput_lo[27407:27392]},
     {otherUnit_maskInput_lo[27391:27376]},
     {otherUnit_maskInput_lo[27375:27360]},
     {otherUnit_maskInput_lo[27359:27344]},
     {otherUnit_maskInput_lo[27343:27328]},
     {otherUnit_maskInput_lo[27327:27312]},
     {otherUnit_maskInput_lo[27311:27296]},
     {otherUnit_maskInput_lo[27295:27280]},
     {otherUnit_maskInput_lo[27279:27264]},
     {otherUnit_maskInput_lo[27263:27248]},
     {otherUnit_maskInput_lo[27247:27232]},
     {otherUnit_maskInput_lo[27231:27216]},
     {otherUnit_maskInput_lo[27215:27200]},
     {otherUnit_maskInput_lo[27199:27184]},
     {otherUnit_maskInput_lo[27183:27168]},
     {otherUnit_maskInput_lo[27167:27152]},
     {otherUnit_maskInput_lo[27151:27136]},
     {otherUnit_maskInput_lo[27135:27120]},
     {otherUnit_maskInput_lo[27119:27104]},
     {otherUnit_maskInput_lo[27103:27088]},
     {otherUnit_maskInput_lo[27087:27072]},
     {otherUnit_maskInput_lo[27071:27056]},
     {otherUnit_maskInput_lo[27055:27040]},
     {otherUnit_maskInput_lo[27039:27024]},
     {otherUnit_maskInput_lo[27023:27008]},
     {otherUnit_maskInput_lo[27007:26992]},
     {otherUnit_maskInput_lo[26991:26976]},
     {otherUnit_maskInput_lo[26975:26960]},
     {otherUnit_maskInput_lo[26959:26944]},
     {otherUnit_maskInput_lo[26943:26928]},
     {otherUnit_maskInput_lo[26927:26912]},
     {otherUnit_maskInput_lo[26911:26896]},
     {otherUnit_maskInput_lo[26895:26880]},
     {otherUnit_maskInput_lo[26879:26864]},
     {otherUnit_maskInput_lo[26863:26848]},
     {otherUnit_maskInput_lo[26847:26832]},
     {otherUnit_maskInput_lo[26831:26816]},
     {otherUnit_maskInput_lo[26815:26800]},
     {otherUnit_maskInput_lo[26799:26784]},
     {otherUnit_maskInput_lo[26783:26768]},
     {otherUnit_maskInput_lo[26767:26752]},
     {otherUnit_maskInput_lo[26751:26736]},
     {otherUnit_maskInput_lo[26735:26720]},
     {otherUnit_maskInput_lo[26719:26704]},
     {otherUnit_maskInput_lo[26703:26688]},
     {otherUnit_maskInput_lo[26687:26672]},
     {otherUnit_maskInput_lo[26671:26656]},
     {otherUnit_maskInput_lo[26655:26640]},
     {otherUnit_maskInput_lo[26639:26624]},
     {otherUnit_maskInput_lo[26623:26608]},
     {otherUnit_maskInput_lo[26607:26592]},
     {otherUnit_maskInput_lo[26591:26576]},
     {otherUnit_maskInput_lo[26575:26560]},
     {otherUnit_maskInput_lo[26559:26544]},
     {otherUnit_maskInput_lo[26543:26528]},
     {otherUnit_maskInput_lo[26527:26512]},
     {otherUnit_maskInput_lo[26511:26496]},
     {otherUnit_maskInput_lo[26495:26480]},
     {otherUnit_maskInput_lo[26479:26464]},
     {otherUnit_maskInput_lo[26463:26448]},
     {otherUnit_maskInput_lo[26447:26432]},
     {otherUnit_maskInput_lo[26431:26416]},
     {otherUnit_maskInput_lo[26415:26400]},
     {otherUnit_maskInput_lo[26399:26384]},
     {otherUnit_maskInput_lo[26383:26368]},
     {otherUnit_maskInput_lo[26367:26352]},
     {otherUnit_maskInput_lo[26351:26336]},
     {otherUnit_maskInput_lo[26335:26320]},
     {otherUnit_maskInput_lo[26319:26304]},
     {otherUnit_maskInput_lo[26303:26288]},
     {otherUnit_maskInput_lo[26287:26272]},
     {otherUnit_maskInput_lo[26271:26256]},
     {otherUnit_maskInput_lo[26255:26240]},
     {otherUnit_maskInput_lo[26239:26224]},
     {otherUnit_maskInput_lo[26223:26208]},
     {otherUnit_maskInput_lo[26207:26192]},
     {otherUnit_maskInput_lo[26191:26176]},
     {otherUnit_maskInput_lo[26175:26160]},
     {otherUnit_maskInput_lo[26159:26144]},
     {otherUnit_maskInput_lo[26143:26128]},
     {otherUnit_maskInput_lo[26127:26112]},
     {otherUnit_maskInput_lo[26111:26096]},
     {otherUnit_maskInput_lo[26095:26080]},
     {otherUnit_maskInput_lo[26079:26064]},
     {otherUnit_maskInput_lo[26063:26048]},
     {otherUnit_maskInput_lo[26047:26032]},
     {otherUnit_maskInput_lo[26031:26016]},
     {otherUnit_maskInput_lo[26015:26000]},
     {otherUnit_maskInput_lo[25999:25984]},
     {otherUnit_maskInput_lo[25983:25968]},
     {otherUnit_maskInput_lo[25967:25952]},
     {otherUnit_maskInput_lo[25951:25936]},
     {otherUnit_maskInput_lo[25935:25920]},
     {otherUnit_maskInput_lo[25919:25904]},
     {otherUnit_maskInput_lo[25903:25888]},
     {otherUnit_maskInput_lo[25887:25872]},
     {otherUnit_maskInput_lo[25871:25856]},
     {otherUnit_maskInput_lo[25855:25840]},
     {otherUnit_maskInput_lo[25839:25824]},
     {otherUnit_maskInput_lo[25823:25808]},
     {otherUnit_maskInput_lo[25807:25792]},
     {otherUnit_maskInput_lo[25791:25776]},
     {otherUnit_maskInput_lo[25775:25760]},
     {otherUnit_maskInput_lo[25759:25744]},
     {otherUnit_maskInput_lo[25743:25728]},
     {otherUnit_maskInput_lo[25727:25712]},
     {otherUnit_maskInput_lo[25711:25696]},
     {otherUnit_maskInput_lo[25695:25680]},
     {otherUnit_maskInput_lo[25679:25664]},
     {otherUnit_maskInput_lo[25663:25648]},
     {otherUnit_maskInput_lo[25647:25632]},
     {otherUnit_maskInput_lo[25631:25616]},
     {otherUnit_maskInput_lo[25615:25600]},
     {otherUnit_maskInput_lo[25599:25584]},
     {otherUnit_maskInput_lo[25583:25568]},
     {otherUnit_maskInput_lo[25567:25552]},
     {otherUnit_maskInput_lo[25551:25536]},
     {otherUnit_maskInput_lo[25535:25520]},
     {otherUnit_maskInput_lo[25519:25504]},
     {otherUnit_maskInput_lo[25503:25488]},
     {otherUnit_maskInput_lo[25487:25472]},
     {otherUnit_maskInput_lo[25471:25456]},
     {otherUnit_maskInput_lo[25455:25440]},
     {otherUnit_maskInput_lo[25439:25424]},
     {otherUnit_maskInput_lo[25423:25408]},
     {otherUnit_maskInput_lo[25407:25392]},
     {otherUnit_maskInput_lo[25391:25376]},
     {otherUnit_maskInput_lo[25375:25360]},
     {otherUnit_maskInput_lo[25359:25344]},
     {otherUnit_maskInput_lo[25343:25328]},
     {otherUnit_maskInput_lo[25327:25312]},
     {otherUnit_maskInput_lo[25311:25296]},
     {otherUnit_maskInput_lo[25295:25280]},
     {otherUnit_maskInput_lo[25279:25264]},
     {otherUnit_maskInput_lo[25263:25248]},
     {otherUnit_maskInput_lo[25247:25232]},
     {otherUnit_maskInput_lo[25231:25216]},
     {otherUnit_maskInput_lo[25215:25200]},
     {otherUnit_maskInput_lo[25199:25184]},
     {otherUnit_maskInput_lo[25183:25168]},
     {otherUnit_maskInput_lo[25167:25152]},
     {otherUnit_maskInput_lo[25151:25136]},
     {otherUnit_maskInput_lo[25135:25120]},
     {otherUnit_maskInput_lo[25119:25104]},
     {otherUnit_maskInput_lo[25103:25088]},
     {otherUnit_maskInput_lo[25087:25072]},
     {otherUnit_maskInput_lo[25071:25056]},
     {otherUnit_maskInput_lo[25055:25040]},
     {otherUnit_maskInput_lo[25039:25024]},
     {otherUnit_maskInput_lo[25023:25008]},
     {otherUnit_maskInput_lo[25007:24992]},
     {otherUnit_maskInput_lo[24991:24976]},
     {otherUnit_maskInput_lo[24975:24960]},
     {otherUnit_maskInput_lo[24959:24944]},
     {otherUnit_maskInput_lo[24943:24928]},
     {otherUnit_maskInput_lo[24927:24912]},
     {otherUnit_maskInput_lo[24911:24896]},
     {otherUnit_maskInput_lo[24895:24880]},
     {otherUnit_maskInput_lo[24879:24864]},
     {otherUnit_maskInput_lo[24863:24848]},
     {otherUnit_maskInput_lo[24847:24832]},
     {otherUnit_maskInput_lo[24831:24816]},
     {otherUnit_maskInput_lo[24815:24800]},
     {otherUnit_maskInput_lo[24799:24784]},
     {otherUnit_maskInput_lo[24783:24768]},
     {otherUnit_maskInput_lo[24767:24752]},
     {otherUnit_maskInput_lo[24751:24736]},
     {otherUnit_maskInput_lo[24735:24720]},
     {otherUnit_maskInput_lo[24719:24704]},
     {otherUnit_maskInput_lo[24703:24688]},
     {otherUnit_maskInput_lo[24687:24672]},
     {otherUnit_maskInput_lo[24671:24656]},
     {otherUnit_maskInput_lo[24655:24640]},
     {otherUnit_maskInput_lo[24639:24624]},
     {otherUnit_maskInput_lo[24623:24608]},
     {otherUnit_maskInput_lo[24607:24592]},
     {otherUnit_maskInput_lo[24591:24576]},
     {otherUnit_maskInput_lo[24575:24560]},
     {otherUnit_maskInput_lo[24559:24544]},
     {otherUnit_maskInput_lo[24543:24528]},
     {otherUnit_maskInput_lo[24527:24512]},
     {otherUnit_maskInput_lo[24511:24496]},
     {otherUnit_maskInput_lo[24495:24480]},
     {otherUnit_maskInput_lo[24479:24464]},
     {otherUnit_maskInput_lo[24463:24448]},
     {otherUnit_maskInput_lo[24447:24432]},
     {otherUnit_maskInput_lo[24431:24416]},
     {otherUnit_maskInput_lo[24415:24400]},
     {otherUnit_maskInput_lo[24399:24384]},
     {otherUnit_maskInput_lo[24383:24368]},
     {otherUnit_maskInput_lo[24367:24352]},
     {otherUnit_maskInput_lo[24351:24336]},
     {otherUnit_maskInput_lo[24335:24320]},
     {otherUnit_maskInput_lo[24319:24304]},
     {otherUnit_maskInput_lo[24303:24288]},
     {otherUnit_maskInput_lo[24287:24272]},
     {otherUnit_maskInput_lo[24271:24256]},
     {otherUnit_maskInput_lo[24255:24240]},
     {otherUnit_maskInput_lo[24239:24224]},
     {otherUnit_maskInput_lo[24223:24208]},
     {otherUnit_maskInput_lo[24207:24192]},
     {otherUnit_maskInput_lo[24191:24176]},
     {otherUnit_maskInput_lo[24175:24160]},
     {otherUnit_maskInput_lo[24159:24144]},
     {otherUnit_maskInput_lo[24143:24128]},
     {otherUnit_maskInput_lo[24127:24112]},
     {otherUnit_maskInput_lo[24111:24096]},
     {otherUnit_maskInput_lo[24095:24080]},
     {otherUnit_maskInput_lo[24079:24064]},
     {otherUnit_maskInput_lo[24063:24048]},
     {otherUnit_maskInput_lo[24047:24032]},
     {otherUnit_maskInput_lo[24031:24016]},
     {otherUnit_maskInput_lo[24015:24000]},
     {otherUnit_maskInput_lo[23999:23984]},
     {otherUnit_maskInput_lo[23983:23968]},
     {otherUnit_maskInput_lo[23967:23952]},
     {otherUnit_maskInput_lo[23951:23936]},
     {otherUnit_maskInput_lo[23935:23920]},
     {otherUnit_maskInput_lo[23919:23904]},
     {otherUnit_maskInput_lo[23903:23888]},
     {otherUnit_maskInput_lo[23887:23872]},
     {otherUnit_maskInput_lo[23871:23856]},
     {otherUnit_maskInput_lo[23855:23840]},
     {otherUnit_maskInput_lo[23839:23824]},
     {otherUnit_maskInput_lo[23823:23808]},
     {otherUnit_maskInput_lo[23807:23792]},
     {otherUnit_maskInput_lo[23791:23776]},
     {otherUnit_maskInput_lo[23775:23760]},
     {otherUnit_maskInput_lo[23759:23744]},
     {otherUnit_maskInput_lo[23743:23728]},
     {otherUnit_maskInput_lo[23727:23712]},
     {otherUnit_maskInput_lo[23711:23696]},
     {otherUnit_maskInput_lo[23695:23680]},
     {otherUnit_maskInput_lo[23679:23664]},
     {otherUnit_maskInput_lo[23663:23648]},
     {otherUnit_maskInput_lo[23647:23632]},
     {otherUnit_maskInput_lo[23631:23616]},
     {otherUnit_maskInput_lo[23615:23600]},
     {otherUnit_maskInput_lo[23599:23584]},
     {otherUnit_maskInput_lo[23583:23568]},
     {otherUnit_maskInput_lo[23567:23552]},
     {otherUnit_maskInput_lo[23551:23536]},
     {otherUnit_maskInput_lo[23535:23520]},
     {otherUnit_maskInput_lo[23519:23504]},
     {otherUnit_maskInput_lo[23503:23488]},
     {otherUnit_maskInput_lo[23487:23472]},
     {otherUnit_maskInput_lo[23471:23456]},
     {otherUnit_maskInput_lo[23455:23440]},
     {otherUnit_maskInput_lo[23439:23424]},
     {otherUnit_maskInput_lo[23423:23408]},
     {otherUnit_maskInput_lo[23407:23392]},
     {otherUnit_maskInput_lo[23391:23376]},
     {otherUnit_maskInput_lo[23375:23360]},
     {otherUnit_maskInput_lo[23359:23344]},
     {otherUnit_maskInput_lo[23343:23328]},
     {otherUnit_maskInput_lo[23327:23312]},
     {otherUnit_maskInput_lo[23311:23296]},
     {otherUnit_maskInput_lo[23295:23280]},
     {otherUnit_maskInput_lo[23279:23264]},
     {otherUnit_maskInput_lo[23263:23248]},
     {otherUnit_maskInput_lo[23247:23232]},
     {otherUnit_maskInput_lo[23231:23216]},
     {otherUnit_maskInput_lo[23215:23200]},
     {otherUnit_maskInput_lo[23199:23184]},
     {otherUnit_maskInput_lo[23183:23168]},
     {otherUnit_maskInput_lo[23167:23152]},
     {otherUnit_maskInput_lo[23151:23136]},
     {otherUnit_maskInput_lo[23135:23120]},
     {otherUnit_maskInput_lo[23119:23104]},
     {otherUnit_maskInput_lo[23103:23088]},
     {otherUnit_maskInput_lo[23087:23072]},
     {otherUnit_maskInput_lo[23071:23056]},
     {otherUnit_maskInput_lo[23055:23040]},
     {otherUnit_maskInput_lo[23039:23024]},
     {otherUnit_maskInput_lo[23023:23008]},
     {otherUnit_maskInput_lo[23007:22992]},
     {otherUnit_maskInput_lo[22991:22976]},
     {otherUnit_maskInput_lo[22975:22960]},
     {otherUnit_maskInput_lo[22959:22944]},
     {otherUnit_maskInput_lo[22943:22928]},
     {otherUnit_maskInput_lo[22927:22912]},
     {otherUnit_maskInput_lo[22911:22896]},
     {otherUnit_maskInput_lo[22895:22880]},
     {otherUnit_maskInput_lo[22879:22864]},
     {otherUnit_maskInput_lo[22863:22848]},
     {otherUnit_maskInput_lo[22847:22832]},
     {otherUnit_maskInput_lo[22831:22816]},
     {otherUnit_maskInput_lo[22815:22800]},
     {otherUnit_maskInput_lo[22799:22784]},
     {otherUnit_maskInput_lo[22783:22768]},
     {otherUnit_maskInput_lo[22767:22752]},
     {otherUnit_maskInput_lo[22751:22736]},
     {otherUnit_maskInput_lo[22735:22720]},
     {otherUnit_maskInput_lo[22719:22704]},
     {otherUnit_maskInput_lo[22703:22688]},
     {otherUnit_maskInput_lo[22687:22672]},
     {otherUnit_maskInput_lo[22671:22656]},
     {otherUnit_maskInput_lo[22655:22640]},
     {otherUnit_maskInput_lo[22639:22624]},
     {otherUnit_maskInput_lo[22623:22608]},
     {otherUnit_maskInput_lo[22607:22592]},
     {otherUnit_maskInput_lo[22591:22576]},
     {otherUnit_maskInput_lo[22575:22560]},
     {otherUnit_maskInput_lo[22559:22544]},
     {otherUnit_maskInput_lo[22543:22528]},
     {otherUnit_maskInput_lo[22527:22512]},
     {otherUnit_maskInput_lo[22511:22496]},
     {otherUnit_maskInput_lo[22495:22480]},
     {otherUnit_maskInput_lo[22479:22464]},
     {otherUnit_maskInput_lo[22463:22448]},
     {otherUnit_maskInput_lo[22447:22432]},
     {otherUnit_maskInput_lo[22431:22416]},
     {otherUnit_maskInput_lo[22415:22400]},
     {otherUnit_maskInput_lo[22399:22384]},
     {otherUnit_maskInput_lo[22383:22368]},
     {otherUnit_maskInput_lo[22367:22352]},
     {otherUnit_maskInput_lo[22351:22336]},
     {otherUnit_maskInput_lo[22335:22320]},
     {otherUnit_maskInput_lo[22319:22304]},
     {otherUnit_maskInput_lo[22303:22288]},
     {otherUnit_maskInput_lo[22287:22272]},
     {otherUnit_maskInput_lo[22271:22256]},
     {otherUnit_maskInput_lo[22255:22240]},
     {otherUnit_maskInput_lo[22239:22224]},
     {otherUnit_maskInput_lo[22223:22208]},
     {otherUnit_maskInput_lo[22207:22192]},
     {otherUnit_maskInput_lo[22191:22176]},
     {otherUnit_maskInput_lo[22175:22160]},
     {otherUnit_maskInput_lo[22159:22144]},
     {otherUnit_maskInput_lo[22143:22128]},
     {otherUnit_maskInput_lo[22127:22112]},
     {otherUnit_maskInput_lo[22111:22096]},
     {otherUnit_maskInput_lo[22095:22080]},
     {otherUnit_maskInput_lo[22079:22064]},
     {otherUnit_maskInput_lo[22063:22048]},
     {otherUnit_maskInput_lo[22047:22032]},
     {otherUnit_maskInput_lo[22031:22016]},
     {otherUnit_maskInput_lo[22015:22000]},
     {otherUnit_maskInput_lo[21999:21984]},
     {otherUnit_maskInput_lo[21983:21968]},
     {otherUnit_maskInput_lo[21967:21952]},
     {otherUnit_maskInput_lo[21951:21936]},
     {otherUnit_maskInput_lo[21935:21920]},
     {otherUnit_maskInput_lo[21919:21904]},
     {otherUnit_maskInput_lo[21903:21888]},
     {otherUnit_maskInput_lo[21887:21872]},
     {otherUnit_maskInput_lo[21871:21856]},
     {otherUnit_maskInput_lo[21855:21840]},
     {otherUnit_maskInput_lo[21839:21824]},
     {otherUnit_maskInput_lo[21823:21808]},
     {otherUnit_maskInput_lo[21807:21792]},
     {otherUnit_maskInput_lo[21791:21776]},
     {otherUnit_maskInput_lo[21775:21760]},
     {otherUnit_maskInput_lo[21759:21744]},
     {otherUnit_maskInput_lo[21743:21728]},
     {otherUnit_maskInput_lo[21727:21712]},
     {otherUnit_maskInput_lo[21711:21696]},
     {otherUnit_maskInput_lo[21695:21680]},
     {otherUnit_maskInput_lo[21679:21664]},
     {otherUnit_maskInput_lo[21663:21648]},
     {otherUnit_maskInput_lo[21647:21632]},
     {otherUnit_maskInput_lo[21631:21616]},
     {otherUnit_maskInput_lo[21615:21600]},
     {otherUnit_maskInput_lo[21599:21584]},
     {otherUnit_maskInput_lo[21583:21568]},
     {otherUnit_maskInput_lo[21567:21552]},
     {otherUnit_maskInput_lo[21551:21536]},
     {otherUnit_maskInput_lo[21535:21520]},
     {otherUnit_maskInput_lo[21519:21504]},
     {otherUnit_maskInput_lo[21503:21488]},
     {otherUnit_maskInput_lo[21487:21472]},
     {otherUnit_maskInput_lo[21471:21456]},
     {otherUnit_maskInput_lo[21455:21440]},
     {otherUnit_maskInput_lo[21439:21424]},
     {otherUnit_maskInput_lo[21423:21408]},
     {otherUnit_maskInput_lo[21407:21392]},
     {otherUnit_maskInput_lo[21391:21376]},
     {otherUnit_maskInput_lo[21375:21360]},
     {otherUnit_maskInput_lo[21359:21344]},
     {otherUnit_maskInput_lo[21343:21328]},
     {otherUnit_maskInput_lo[21327:21312]},
     {otherUnit_maskInput_lo[21311:21296]},
     {otherUnit_maskInput_lo[21295:21280]},
     {otherUnit_maskInput_lo[21279:21264]},
     {otherUnit_maskInput_lo[21263:21248]},
     {otherUnit_maskInput_lo[21247:21232]},
     {otherUnit_maskInput_lo[21231:21216]},
     {otherUnit_maskInput_lo[21215:21200]},
     {otherUnit_maskInput_lo[21199:21184]},
     {otherUnit_maskInput_lo[21183:21168]},
     {otherUnit_maskInput_lo[21167:21152]},
     {otherUnit_maskInput_lo[21151:21136]},
     {otherUnit_maskInput_lo[21135:21120]},
     {otherUnit_maskInput_lo[21119:21104]},
     {otherUnit_maskInput_lo[21103:21088]},
     {otherUnit_maskInput_lo[21087:21072]},
     {otherUnit_maskInput_lo[21071:21056]},
     {otherUnit_maskInput_lo[21055:21040]},
     {otherUnit_maskInput_lo[21039:21024]},
     {otherUnit_maskInput_lo[21023:21008]},
     {otherUnit_maskInput_lo[21007:20992]},
     {otherUnit_maskInput_lo[20991:20976]},
     {otherUnit_maskInput_lo[20975:20960]},
     {otherUnit_maskInput_lo[20959:20944]},
     {otherUnit_maskInput_lo[20943:20928]},
     {otherUnit_maskInput_lo[20927:20912]},
     {otherUnit_maskInput_lo[20911:20896]},
     {otherUnit_maskInput_lo[20895:20880]},
     {otherUnit_maskInput_lo[20879:20864]},
     {otherUnit_maskInput_lo[20863:20848]},
     {otherUnit_maskInput_lo[20847:20832]},
     {otherUnit_maskInput_lo[20831:20816]},
     {otherUnit_maskInput_lo[20815:20800]},
     {otherUnit_maskInput_lo[20799:20784]},
     {otherUnit_maskInput_lo[20783:20768]},
     {otherUnit_maskInput_lo[20767:20752]},
     {otherUnit_maskInput_lo[20751:20736]},
     {otherUnit_maskInput_lo[20735:20720]},
     {otherUnit_maskInput_lo[20719:20704]},
     {otherUnit_maskInput_lo[20703:20688]},
     {otherUnit_maskInput_lo[20687:20672]},
     {otherUnit_maskInput_lo[20671:20656]},
     {otherUnit_maskInput_lo[20655:20640]},
     {otherUnit_maskInput_lo[20639:20624]},
     {otherUnit_maskInput_lo[20623:20608]},
     {otherUnit_maskInput_lo[20607:20592]},
     {otherUnit_maskInput_lo[20591:20576]},
     {otherUnit_maskInput_lo[20575:20560]},
     {otherUnit_maskInput_lo[20559:20544]},
     {otherUnit_maskInput_lo[20543:20528]},
     {otherUnit_maskInput_lo[20527:20512]},
     {otherUnit_maskInput_lo[20511:20496]},
     {otherUnit_maskInput_lo[20495:20480]},
     {otherUnit_maskInput_lo[20479:20464]},
     {otherUnit_maskInput_lo[20463:20448]},
     {otherUnit_maskInput_lo[20447:20432]},
     {otherUnit_maskInput_lo[20431:20416]},
     {otherUnit_maskInput_lo[20415:20400]},
     {otherUnit_maskInput_lo[20399:20384]},
     {otherUnit_maskInput_lo[20383:20368]},
     {otherUnit_maskInput_lo[20367:20352]},
     {otherUnit_maskInput_lo[20351:20336]},
     {otherUnit_maskInput_lo[20335:20320]},
     {otherUnit_maskInput_lo[20319:20304]},
     {otherUnit_maskInput_lo[20303:20288]},
     {otherUnit_maskInput_lo[20287:20272]},
     {otherUnit_maskInput_lo[20271:20256]},
     {otherUnit_maskInput_lo[20255:20240]},
     {otherUnit_maskInput_lo[20239:20224]},
     {otherUnit_maskInput_lo[20223:20208]},
     {otherUnit_maskInput_lo[20207:20192]},
     {otherUnit_maskInput_lo[20191:20176]},
     {otherUnit_maskInput_lo[20175:20160]},
     {otherUnit_maskInput_lo[20159:20144]},
     {otherUnit_maskInput_lo[20143:20128]},
     {otherUnit_maskInput_lo[20127:20112]},
     {otherUnit_maskInput_lo[20111:20096]},
     {otherUnit_maskInput_lo[20095:20080]},
     {otherUnit_maskInput_lo[20079:20064]},
     {otherUnit_maskInput_lo[20063:20048]},
     {otherUnit_maskInput_lo[20047:20032]},
     {otherUnit_maskInput_lo[20031:20016]},
     {otherUnit_maskInput_lo[20015:20000]},
     {otherUnit_maskInput_lo[19999:19984]},
     {otherUnit_maskInput_lo[19983:19968]},
     {otherUnit_maskInput_lo[19967:19952]},
     {otherUnit_maskInput_lo[19951:19936]},
     {otherUnit_maskInput_lo[19935:19920]},
     {otherUnit_maskInput_lo[19919:19904]},
     {otherUnit_maskInput_lo[19903:19888]},
     {otherUnit_maskInput_lo[19887:19872]},
     {otherUnit_maskInput_lo[19871:19856]},
     {otherUnit_maskInput_lo[19855:19840]},
     {otherUnit_maskInput_lo[19839:19824]},
     {otherUnit_maskInput_lo[19823:19808]},
     {otherUnit_maskInput_lo[19807:19792]},
     {otherUnit_maskInput_lo[19791:19776]},
     {otherUnit_maskInput_lo[19775:19760]},
     {otherUnit_maskInput_lo[19759:19744]},
     {otherUnit_maskInput_lo[19743:19728]},
     {otherUnit_maskInput_lo[19727:19712]},
     {otherUnit_maskInput_lo[19711:19696]},
     {otherUnit_maskInput_lo[19695:19680]},
     {otherUnit_maskInput_lo[19679:19664]},
     {otherUnit_maskInput_lo[19663:19648]},
     {otherUnit_maskInput_lo[19647:19632]},
     {otherUnit_maskInput_lo[19631:19616]},
     {otherUnit_maskInput_lo[19615:19600]},
     {otherUnit_maskInput_lo[19599:19584]},
     {otherUnit_maskInput_lo[19583:19568]},
     {otherUnit_maskInput_lo[19567:19552]},
     {otherUnit_maskInput_lo[19551:19536]},
     {otherUnit_maskInput_lo[19535:19520]},
     {otherUnit_maskInput_lo[19519:19504]},
     {otherUnit_maskInput_lo[19503:19488]},
     {otherUnit_maskInput_lo[19487:19472]},
     {otherUnit_maskInput_lo[19471:19456]},
     {otherUnit_maskInput_lo[19455:19440]},
     {otherUnit_maskInput_lo[19439:19424]},
     {otherUnit_maskInput_lo[19423:19408]},
     {otherUnit_maskInput_lo[19407:19392]},
     {otherUnit_maskInput_lo[19391:19376]},
     {otherUnit_maskInput_lo[19375:19360]},
     {otherUnit_maskInput_lo[19359:19344]},
     {otherUnit_maskInput_lo[19343:19328]},
     {otherUnit_maskInput_lo[19327:19312]},
     {otherUnit_maskInput_lo[19311:19296]},
     {otherUnit_maskInput_lo[19295:19280]},
     {otherUnit_maskInput_lo[19279:19264]},
     {otherUnit_maskInput_lo[19263:19248]},
     {otherUnit_maskInput_lo[19247:19232]},
     {otherUnit_maskInput_lo[19231:19216]},
     {otherUnit_maskInput_lo[19215:19200]},
     {otherUnit_maskInput_lo[19199:19184]},
     {otherUnit_maskInput_lo[19183:19168]},
     {otherUnit_maskInput_lo[19167:19152]},
     {otherUnit_maskInput_lo[19151:19136]},
     {otherUnit_maskInput_lo[19135:19120]},
     {otherUnit_maskInput_lo[19119:19104]},
     {otherUnit_maskInput_lo[19103:19088]},
     {otherUnit_maskInput_lo[19087:19072]},
     {otherUnit_maskInput_lo[19071:19056]},
     {otherUnit_maskInput_lo[19055:19040]},
     {otherUnit_maskInput_lo[19039:19024]},
     {otherUnit_maskInput_lo[19023:19008]},
     {otherUnit_maskInput_lo[19007:18992]},
     {otherUnit_maskInput_lo[18991:18976]},
     {otherUnit_maskInput_lo[18975:18960]},
     {otherUnit_maskInput_lo[18959:18944]},
     {otherUnit_maskInput_lo[18943:18928]},
     {otherUnit_maskInput_lo[18927:18912]},
     {otherUnit_maskInput_lo[18911:18896]},
     {otherUnit_maskInput_lo[18895:18880]},
     {otherUnit_maskInput_lo[18879:18864]},
     {otherUnit_maskInput_lo[18863:18848]},
     {otherUnit_maskInput_lo[18847:18832]},
     {otherUnit_maskInput_lo[18831:18816]},
     {otherUnit_maskInput_lo[18815:18800]},
     {otherUnit_maskInput_lo[18799:18784]},
     {otherUnit_maskInput_lo[18783:18768]},
     {otherUnit_maskInput_lo[18767:18752]},
     {otherUnit_maskInput_lo[18751:18736]},
     {otherUnit_maskInput_lo[18735:18720]},
     {otherUnit_maskInput_lo[18719:18704]},
     {otherUnit_maskInput_lo[18703:18688]},
     {otherUnit_maskInput_lo[18687:18672]},
     {otherUnit_maskInput_lo[18671:18656]},
     {otherUnit_maskInput_lo[18655:18640]},
     {otherUnit_maskInput_lo[18639:18624]},
     {otherUnit_maskInput_lo[18623:18608]},
     {otherUnit_maskInput_lo[18607:18592]},
     {otherUnit_maskInput_lo[18591:18576]},
     {otherUnit_maskInput_lo[18575:18560]},
     {otherUnit_maskInput_lo[18559:18544]},
     {otherUnit_maskInput_lo[18543:18528]},
     {otherUnit_maskInput_lo[18527:18512]},
     {otherUnit_maskInput_lo[18511:18496]},
     {otherUnit_maskInput_lo[18495:18480]},
     {otherUnit_maskInput_lo[18479:18464]},
     {otherUnit_maskInput_lo[18463:18448]},
     {otherUnit_maskInput_lo[18447:18432]},
     {otherUnit_maskInput_lo[18431:18416]},
     {otherUnit_maskInput_lo[18415:18400]},
     {otherUnit_maskInput_lo[18399:18384]},
     {otherUnit_maskInput_lo[18383:18368]},
     {otherUnit_maskInput_lo[18367:18352]},
     {otherUnit_maskInput_lo[18351:18336]},
     {otherUnit_maskInput_lo[18335:18320]},
     {otherUnit_maskInput_lo[18319:18304]},
     {otherUnit_maskInput_lo[18303:18288]},
     {otherUnit_maskInput_lo[18287:18272]},
     {otherUnit_maskInput_lo[18271:18256]},
     {otherUnit_maskInput_lo[18255:18240]},
     {otherUnit_maskInput_lo[18239:18224]},
     {otherUnit_maskInput_lo[18223:18208]},
     {otherUnit_maskInput_lo[18207:18192]},
     {otherUnit_maskInput_lo[18191:18176]},
     {otherUnit_maskInput_lo[18175:18160]},
     {otherUnit_maskInput_lo[18159:18144]},
     {otherUnit_maskInput_lo[18143:18128]},
     {otherUnit_maskInput_lo[18127:18112]},
     {otherUnit_maskInput_lo[18111:18096]},
     {otherUnit_maskInput_lo[18095:18080]},
     {otherUnit_maskInput_lo[18079:18064]},
     {otherUnit_maskInput_lo[18063:18048]},
     {otherUnit_maskInput_lo[18047:18032]},
     {otherUnit_maskInput_lo[18031:18016]},
     {otherUnit_maskInput_lo[18015:18000]},
     {otherUnit_maskInput_lo[17999:17984]},
     {otherUnit_maskInput_lo[17983:17968]},
     {otherUnit_maskInput_lo[17967:17952]},
     {otherUnit_maskInput_lo[17951:17936]},
     {otherUnit_maskInput_lo[17935:17920]},
     {otherUnit_maskInput_lo[17919:17904]},
     {otherUnit_maskInput_lo[17903:17888]},
     {otherUnit_maskInput_lo[17887:17872]},
     {otherUnit_maskInput_lo[17871:17856]},
     {otherUnit_maskInput_lo[17855:17840]},
     {otherUnit_maskInput_lo[17839:17824]},
     {otherUnit_maskInput_lo[17823:17808]},
     {otherUnit_maskInput_lo[17807:17792]},
     {otherUnit_maskInput_lo[17791:17776]},
     {otherUnit_maskInput_lo[17775:17760]},
     {otherUnit_maskInput_lo[17759:17744]},
     {otherUnit_maskInput_lo[17743:17728]},
     {otherUnit_maskInput_lo[17727:17712]},
     {otherUnit_maskInput_lo[17711:17696]},
     {otherUnit_maskInput_lo[17695:17680]},
     {otherUnit_maskInput_lo[17679:17664]},
     {otherUnit_maskInput_lo[17663:17648]},
     {otherUnit_maskInput_lo[17647:17632]},
     {otherUnit_maskInput_lo[17631:17616]},
     {otherUnit_maskInput_lo[17615:17600]},
     {otherUnit_maskInput_lo[17599:17584]},
     {otherUnit_maskInput_lo[17583:17568]},
     {otherUnit_maskInput_lo[17567:17552]},
     {otherUnit_maskInput_lo[17551:17536]},
     {otherUnit_maskInput_lo[17535:17520]},
     {otherUnit_maskInput_lo[17519:17504]},
     {otherUnit_maskInput_lo[17503:17488]},
     {otherUnit_maskInput_lo[17487:17472]},
     {otherUnit_maskInput_lo[17471:17456]},
     {otherUnit_maskInput_lo[17455:17440]},
     {otherUnit_maskInput_lo[17439:17424]},
     {otherUnit_maskInput_lo[17423:17408]},
     {otherUnit_maskInput_lo[17407:17392]},
     {otherUnit_maskInput_lo[17391:17376]},
     {otherUnit_maskInput_lo[17375:17360]},
     {otherUnit_maskInput_lo[17359:17344]},
     {otherUnit_maskInput_lo[17343:17328]},
     {otherUnit_maskInput_lo[17327:17312]},
     {otherUnit_maskInput_lo[17311:17296]},
     {otherUnit_maskInput_lo[17295:17280]},
     {otherUnit_maskInput_lo[17279:17264]},
     {otherUnit_maskInput_lo[17263:17248]},
     {otherUnit_maskInput_lo[17247:17232]},
     {otherUnit_maskInput_lo[17231:17216]},
     {otherUnit_maskInput_lo[17215:17200]},
     {otherUnit_maskInput_lo[17199:17184]},
     {otherUnit_maskInput_lo[17183:17168]},
     {otherUnit_maskInput_lo[17167:17152]},
     {otherUnit_maskInput_lo[17151:17136]},
     {otherUnit_maskInput_lo[17135:17120]},
     {otherUnit_maskInput_lo[17119:17104]},
     {otherUnit_maskInput_lo[17103:17088]},
     {otherUnit_maskInput_lo[17087:17072]},
     {otherUnit_maskInput_lo[17071:17056]},
     {otherUnit_maskInput_lo[17055:17040]},
     {otherUnit_maskInput_lo[17039:17024]},
     {otherUnit_maskInput_lo[17023:17008]},
     {otherUnit_maskInput_lo[17007:16992]},
     {otherUnit_maskInput_lo[16991:16976]},
     {otherUnit_maskInput_lo[16975:16960]},
     {otherUnit_maskInput_lo[16959:16944]},
     {otherUnit_maskInput_lo[16943:16928]},
     {otherUnit_maskInput_lo[16927:16912]},
     {otherUnit_maskInput_lo[16911:16896]},
     {otherUnit_maskInput_lo[16895:16880]},
     {otherUnit_maskInput_lo[16879:16864]},
     {otherUnit_maskInput_lo[16863:16848]},
     {otherUnit_maskInput_lo[16847:16832]},
     {otherUnit_maskInput_lo[16831:16816]},
     {otherUnit_maskInput_lo[16815:16800]},
     {otherUnit_maskInput_lo[16799:16784]},
     {otherUnit_maskInput_lo[16783:16768]},
     {otherUnit_maskInput_lo[16767:16752]},
     {otherUnit_maskInput_lo[16751:16736]},
     {otherUnit_maskInput_lo[16735:16720]},
     {otherUnit_maskInput_lo[16719:16704]},
     {otherUnit_maskInput_lo[16703:16688]},
     {otherUnit_maskInput_lo[16687:16672]},
     {otherUnit_maskInput_lo[16671:16656]},
     {otherUnit_maskInput_lo[16655:16640]},
     {otherUnit_maskInput_lo[16639:16624]},
     {otherUnit_maskInput_lo[16623:16608]},
     {otherUnit_maskInput_lo[16607:16592]},
     {otherUnit_maskInput_lo[16591:16576]},
     {otherUnit_maskInput_lo[16575:16560]},
     {otherUnit_maskInput_lo[16559:16544]},
     {otherUnit_maskInput_lo[16543:16528]},
     {otherUnit_maskInput_lo[16527:16512]},
     {otherUnit_maskInput_lo[16511:16496]},
     {otherUnit_maskInput_lo[16495:16480]},
     {otherUnit_maskInput_lo[16479:16464]},
     {otherUnit_maskInput_lo[16463:16448]},
     {otherUnit_maskInput_lo[16447:16432]},
     {otherUnit_maskInput_lo[16431:16416]},
     {otherUnit_maskInput_lo[16415:16400]},
     {otherUnit_maskInput_lo[16399:16384]},
     {otherUnit_maskInput_lo[16383:16368]},
     {otherUnit_maskInput_lo[16367:16352]},
     {otherUnit_maskInput_lo[16351:16336]},
     {otherUnit_maskInput_lo[16335:16320]},
     {otherUnit_maskInput_lo[16319:16304]},
     {otherUnit_maskInput_lo[16303:16288]},
     {otherUnit_maskInput_lo[16287:16272]},
     {otherUnit_maskInput_lo[16271:16256]},
     {otherUnit_maskInput_lo[16255:16240]},
     {otherUnit_maskInput_lo[16239:16224]},
     {otherUnit_maskInput_lo[16223:16208]},
     {otherUnit_maskInput_lo[16207:16192]},
     {otherUnit_maskInput_lo[16191:16176]},
     {otherUnit_maskInput_lo[16175:16160]},
     {otherUnit_maskInput_lo[16159:16144]},
     {otherUnit_maskInput_lo[16143:16128]},
     {otherUnit_maskInput_lo[16127:16112]},
     {otherUnit_maskInput_lo[16111:16096]},
     {otherUnit_maskInput_lo[16095:16080]},
     {otherUnit_maskInput_lo[16079:16064]},
     {otherUnit_maskInput_lo[16063:16048]},
     {otherUnit_maskInput_lo[16047:16032]},
     {otherUnit_maskInput_lo[16031:16016]},
     {otherUnit_maskInput_lo[16015:16000]},
     {otherUnit_maskInput_lo[15999:15984]},
     {otherUnit_maskInput_lo[15983:15968]},
     {otherUnit_maskInput_lo[15967:15952]},
     {otherUnit_maskInput_lo[15951:15936]},
     {otherUnit_maskInput_lo[15935:15920]},
     {otherUnit_maskInput_lo[15919:15904]},
     {otherUnit_maskInput_lo[15903:15888]},
     {otherUnit_maskInput_lo[15887:15872]},
     {otherUnit_maskInput_lo[15871:15856]},
     {otherUnit_maskInput_lo[15855:15840]},
     {otherUnit_maskInput_lo[15839:15824]},
     {otherUnit_maskInput_lo[15823:15808]},
     {otherUnit_maskInput_lo[15807:15792]},
     {otherUnit_maskInput_lo[15791:15776]},
     {otherUnit_maskInput_lo[15775:15760]},
     {otherUnit_maskInput_lo[15759:15744]},
     {otherUnit_maskInput_lo[15743:15728]},
     {otherUnit_maskInput_lo[15727:15712]},
     {otherUnit_maskInput_lo[15711:15696]},
     {otherUnit_maskInput_lo[15695:15680]},
     {otherUnit_maskInput_lo[15679:15664]},
     {otherUnit_maskInput_lo[15663:15648]},
     {otherUnit_maskInput_lo[15647:15632]},
     {otherUnit_maskInput_lo[15631:15616]},
     {otherUnit_maskInput_lo[15615:15600]},
     {otherUnit_maskInput_lo[15599:15584]},
     {otherUnit_maskInput_lo[15583:15568]},
     {otherUnit_maskInput_lo[15567:15552]},
     {otherUnit_maskInput_lo[15551:15536]},
     {otherUnit_maskInput_lo[15535:15520]},
     {otherUnit_maskInput_lo[15519:15504]},
     {otherUnit_maskInput_lo[15503:15488]},
     {otherUnit_maskInput_lo[15487:15472]},
     {otherUnit_maskInput_lo[15471:15456]},
     {otherUnit_maskInput_lo[15455:15440]},
     {otherUnit_maskInput_lo[15439:15424]},
     {otherUnit_maskInput_lo[15423:15408]},
     {otherUnit_maskInput_lo[15407:15392]},
     {otherUnit_maskInput_lo[15391:15376]},
     {otherUnit_maskInput_lo[15375:15360]},
     {otherUnit_maskInput_lo[15359:15344]},
     {otherUnit_maskInput_lo[15343:15328]},
     {otherUnit_maskInput_lo[15327:15312]},
     {otherUnit_maskInput_lo[15311:15296]},
     {otherUnit_maskInput_lo[15295:15280]},
     {otherUnit_maskInput_lo[15279:15264]},
     {otherUnit_maskInput_lo[15263:15248]},
     {otherUnit_maskInput_lo[15247:15232]},
     {otherUnit_maskInput_lo[15231:15216]},
     {otherUnit_maskInput_lo[15215:15200]},
     {otherUnit_maskInput_lo[15199:15184]},
     {otherUnit_maskInput_lo[15183:15168]},
     {otherUnit_maskInput_lo[15167:15152]},
     {otherUnit_maskInput_lo[15151:15136]},
     {otherUnit_maskInput_lo[15135:15120]},
     {otherUnit_maskInput_lo[15119:15104]},
     {otherUnit_maskInput_lo[15103:15088]},
     {otherUnit_maskInput_lo[15087:15072]},
     {otherUnit_maskInput_lo[15071:15056]},
     {otherUnit_maskInput_lo[15055:15040]},
     {otherUnit_maskInput_lo[15039:15024]},
     {otherUnit_maskInput_lo[15023:15008]},
     {otherUnit_maskInput_lo[15007:14992]},
     {otherUnit_maskInput_lo[14991:14976]},
     {otherUnit_maskInput_lo[14975:14960]},
     {otherUnit_maskInput_lo[14959:14944]},
     {otherUnit_maskInput_lo[14943:14928]},
     {otherUnit_maskInput_lo[14927:14912]},
     {otherUnit_maskInput_lo[14911:14896]},
     {otherUnit_maskInput_lo[14895:14880]},
     {otherUnit_maskInput_lo[14879:14864]},
     {otherUnit_maskInput_lo[14863:14848]},
     {otherUnit_maskInput_lo[14847:14832]},
     {otherUnit_maskInput_lo[14831:14816]},
     {otherUnit_maskInput_lo[14815:14800]},
     {otherUnit_maskInput_lo[14799:14784]},
     {otherUnit_maskInput_lo[14783:14768]},
     {otherUnit_maskInput_lo[14767:14752]},
     {otherUnit_maskInput_lo[14751:14736]},
     {otherUnit_maskInput_lo[14735:14720]},
     {otherUnit_maskInput_lo[14719:14704]},
     {otherUnit_maskInput_lo[14703:14688]},
     {otherUnit_maskInput_lo[14687:14672]},
     {otherUnit_maskInput_lo[14671:14656]},
     {otherUnit_maskInput_lo[14655:14640]},
     {otherUnit_maskInput_lo[14639:14624]},
     {otherUnit_maskInput_lo[14623:14608]},
     {otherUnit_maskInput_lo[14607:14592]},
     {otherUnit_maskInput_lo[14591:14576]},
     {otherUnit_maskInput_lo[14575:14560]},
     {otherUnit_maskInput_lo[14559:14544]},
     {otherUnit_maskInput_lo[14543:14528]},
     {otherUnit_maskInput_lo[14527:14512]},
     {otherUnit_maskInput_lo[14511:14496]},
     {otherUnit_maskInput_lo[14495:14480]},
     {otherUnit_maskInput_lo[14479:14464]},
     {otherUnit_maskInput_lo[14463:14448]},
     {otherUnit_maskInput_lo[14447:14432]},
     {otherUnit_maskInput_lo[14431:14416]},
     {otherUnit_maskInput_lo[14415:14400]},
     {otherUnit_maskInput_lo[14399:14384]},
     {otherUnit_maskInput_lo[14383:14368]},
     {otherUnit_maskInput_lo[14367:14352]},
     {otherUnit_maskInput_lo[14351:14336]},
     {otherUnit_maskInput_lo[14335:14320]},
     {otherUnit_maskInput_lo[14319:14304]},
     {otherUnit_maskInput_lo[14303:14288]},
     {otherUnit_maskInput_lo[14287:14272]},
     {otherUnit_maskInput_lo[14271:14256]},
     {otherUnit_maskInput_lo[14255:14240]},
     {otherUnit_maskInput_lo[14239:14224]},
     {otherUnit_maskInput_lo[14223:14208]},
     {otherUnit_maskInput_lo[14207:14192]},
     {otherUnit_maskInput_lo[14191:14176]},
     {otherUnit_maskInput_lo[14175:14160]},
     {otherUnit_maskInput_lo[14159:14144]},
     {otherUnit_maskInput_lo[14143:14128]},
     {otherUnit_maskInput_lo[14127:14112]},
     {otherUnit_maskInput_lo[14111:14096]},
     {otherUnit_maskInput_lo[14095:14080]},
     {otherUnit_maskInput_lo[14079:14064]},
     {otherUnit_maskInput_lo[14063:14048]},
     {otherUnit_maskInput_lo[14047:14032]},
     {otherUnit_maskInput_lo[14031:14016]},
     {otherUnit_maskInput_lo[14015:14000]},
     {otherUnit_maskInput_lo[13999:13984]},
     {otherUnit_maskInput_lo[13983:13968]},
     {otherUnit_maskInput_lo[13967:13952]},
     {otherUnit_maskInput_lo[13951:13936]},
     {otherUnit_maskInput_lo[13935:13920]},
     {otherUnit_maskInput_lo[13919:13904]},
     {otherUnit_maskInput_lo[13903:13888]},
     {otherUnit_maskInput_lo[13887:13872]},
     {otherUnit_maskInput_lo[13871:13856]},
     {otherUnit_maskInput_lo[13855:13840]},
     {otherUnit_maskInput_lo[13839:13824]},
     {otherUnit_maskInput_lo[13823:13808]},
     {otherUnit_maskInput_lo[13807:13792]},
     {otherUnit_maskInput_lo[13791:13776]},
     {otherUnit_maskInput_lo[13775:13760]},
     {otherUnit_maskInput_lo[13759:13744]},
     {otherUnit_maskInput_lo[13743:13728]},
     {otherUnit_maskInput_lo[13727:13712]},
     {otherUnit_maskInput_lo[13711:13696]},
     {otherUnit_maskInput_lo[13695:13680]},
     {otherUnit_maskInput_lo[13679:13664]},
     {otherUnit_maskInput_lo[13663:13648]},
     {otherUnit_maskInput_lo[13647:13632]},
     {otherUnit_maskInput_lo[13631:13616]},
     {otherUnit_maskInput_lo[13615:13600]},
     {otherUnit_maskInput_lo[13599:13584]},
     {otherUnit_maskInput_lo[13583:13568]},
     {otherUnit_maskInput_lo[13567:13552]},
     {otherUnit_maskInput_lo[13551:13536]},
     {otherUnit_maskInput_lo[13535:13520]},
     {otherUnit_maskInput_lo[13519:13504]},
     {otherUnit_maskInput_lo[13503:13488]},
     {otherUnit_maskInput_lo[13487:13472]},
     {otherUnit_maskInput_lo[13471:13456]},
     {otherUnit_maskInput_lo[13455:13440]},
     {otherUnit_maskInput_lo[13439:13424]},
     {otherUnit_maskInput_lo[13423:13408]},
     {otherUnit_maskInput_lo[13407:13392]},
     {otherUnit_maskInput_lo[13391:13376]},
     {otherUnit_maskInput_lo[13375:13360]},
     {otherUnit_maskInput_lo[13359:13344]},
     {otherUnit_maskInput_lo[13343:13328]},
     {otherUnit_maskInput_lo[13327:13312]},
     {otherUnit_maskInput_lo[13311:13296]},
     {otherUnit_maskInput_lo[13295:13280]},
     {otherUnit_maskInput_lo[13279:13264]},
     {otherUnit_maskInput_lo[13263:13248]},
     {otherUnit_maskInput_lo[13247:13232]},
     {otherUnit_maskInput_lo[13231:13216]},
     {otherUnit_maskInput_lo[13215:13200]},
     {otherUnit_maskInput_lo[13199:13184]},
     {otherUnit_maskInput_lo[13183:13168]},
     {otherUnit_maskInput_lo[13167:13152]},
     {otherUnit_maskInput_lo[13151:13136]},
     {otherUnit_maskInput_lo[13135:13120]},
     {otherUnit_maskInput_lo[13119:13104]},
     {otherUnit_maskInput_lo[13103:13088]},
     {otherUnit_maskInput_lo[13087:13072]},
     {otherUnit_maskInput_lo[13071:13056]},
     {otherUnit_maskInput_lo[13055:13040]},
     {otherUnit_maskInput_lo[13039:13024]},
     {otherUnit_maskInput_lo[13023:13008]},
     {otherUnit_maskInput_lo[13007:12992]},
     {otherUnit_maskInput_lo[12991:12976]},
     {otherUnit_maskInput_lo[12975:12960]},
     {otherUnit_maskInput_lo[12959:12944]},
     {otherUnit_maskInput_lo[12943:12928]},
     {otherUnit_maskInput_lo[12927:12912]},
     {otherUnit_maskInput_lo[12911:12896]},
     {otherUnit_maskInput_lo[12895:12880]},
     {otherUnit_maskInput_lo[12879:12864]},
     {otherUnit_maskInput_lo[12863:12848]},
     {otherUnit_maskInput_lo[12847:12832]},
     {otherUnit_maskInput_lo[12831:12816]},
     {otherUnit_maskInput_lo[12815:12800]},
     {otherUnit_maskInput_lo[12799:12784]},
     {otherUnit_maskInput_lo[12783:12768]},
     {otherUnit_maskInput_lo[12767:12752]},
     {otherUnit_maskInput_lo[12751:12736]},
     {otherUnit_maskInput_lo[12735:12720]},
     {otherUnit_maskInput_lo[12719:12704]},
     {otherUnit_maskInput_lo[12703:12688]},
     {otherUnit_maskInput_lo[12687:12672]},
     {otherUnit_maskInput_lo[12671:12656]},
     {otherUnit_maskInput_lo[12655:12640]},
     {otherUnit_maskInput_lo[12639:12624]},
     {otherUnit_maskInput_lo[12623:12608]},
     {otherUnit_maskInput_lo[12607:12592]},
     {otherUnit_maskInput_lo[12591:12576]},
     {otherUnit_maskInput_lo[12575:12560]},
     {otherUnit_maskInput_lo[12559:12544]},
     {otherUnit_maskInput_lo[12543:12528]},
     {otherUnit_maskInput_lo[12527:12512]},
     {otherUnit_maskInput_lo[12511:12496]},
     {otherUnit_maskInput_lo[12495:12480]},
     {otherUnit_maskInput_lo[12479:12464]},
     {otherUnit_maskInput_lo[12463:12448]},
     {otherUnit_maskInput_lo[12447:12432]},
     {otherUnit_maskInput_lo[12431:12416]},
     {otherUnit_maskInput_lo[12415:12400]},
     {otherUnit_maskInput_lo[12399:12384]},
     {otherUnit_maskInput_lo[12383:12368]},
     {otherUnit_maskInput_lo[12367:12352]},
     {otherUnit_maskInput_lo[12351:12336]},
     {otherUnit_maskInput_lo[12335:12320]},
     {otherUnit_maskInput_lo[12319:12304]},
     {otherUnit_maskInput_lo[12303:12288]},
     {otherUnit_maskInput_lo[12287:12272]},
     {otherUnit_maskInput_lo[12271:12256]},
     {otherUnit_maskInput_lo[12255:12240]},
     {otherUnit_maskInput_lo[12239:12224]},
     {otherUnit_maskInput_lo[12223:12208]},
     {otherUnit_maskInput_lo[12207:12192]},
     {otherUnit_maskInput_lo[12191:12176]},
     {otherUnit_maskInput_lo[12175:12160]},
     {otherUnit_maskInput_lo[12159:12144]},
     {otherUnit_maskInput_lo[12143:12128]},
     {otherUnit_maskInput_lo[12127:12112]},
     {otherUnit_maskInput_lo[12111:12096]},
     {otherUnit_maskInput_lo[12095:12080]},
     {otherUnit_maskInput_lo[12079:12064]},
     {otherUnit_maskInput_lo[12063:12048]},
     {otherUnit_maskInput_lo[12047:12032]},
     {otherUnit_maskInput_lo[12031:12016]},
     {otherUnit_maskInput_lo[12015:12000]},
     {otherUnit_maskInput_lo[11999:11984]},
     {otherUnit_maskInput_lo[11983:11968]},
     {otherUnit_maskInput_lo[11967:11952]},
     {otherUnit_maskInput_lo[11951:11936]},
     {otherUnit_maskInput_lo[11935:11920]},
     {otherUnit_maskInput_lo[11919:11904]},
     {otherUnit_maskInput_lo[11903:11888]},
     {otherUnit_maskInput_lo[11887:11872]},
     {otherUnit_maskInput_lo[11871:11856]},
     {otherUnit_maskInput_lo[11855:11840]},
     {otherUnit_maskInput_lo[11839:11824]},
     {otherUnit_maskInput_lo[11823:11808]},
     {otherUnit_maskInput_lo[11807:11792]},
     {otherUnit_maskInput_lo[11791:11776]},
     {otherUnit_maskInput_lo[11775:11760]},
     {otherUnit_maskInput_lo[11759:11744]},
     {otherUnit_maskInput_lo[11743:11728]},
     {otherUnit_maskInput_lo[11727:11712]},
     {otherUnit_maskInput_lo[11711:11696]},
     {otherUnit_maskInput_lo[11695:11680]},
     {otherUnit_maskInput_lo[11679:11664]},
     {otherUnit_maskInput_lo[11663:11648]},
     {otherUnit_maskInput_lo[11647:11632]},
     {otherUnit_maskInput_lo[11631:11616]},
     {otherUnit_maskInput_lo[11615:11600]},
     {otherUnit_maskInput_lo[11599:11584]},
     {otherUnit_maskInput_lo[11583:11568]},
     {otherUnit_maskInput_lo[11567:11552]},
     {otherUnit_maskInput_lo[11551:11536]},
     {otherUnit_maskInput_lo[11535:11520]},
     {otherUnit_maskInput_lo[11519:11504]},
     {otherUnit_maskInput_lo[11503:11488]},
     {otherUnit_maskInput_lo[11487:11472]},
     {otherUnit_maskInput_lo[11471:11456]},
     {otherUnit_maskInput_lo[11455:11440]},
     {otherUnit_maskInput_lo[11439:11424]},
     {otherUnit_maskInput_lo[11423:11408]},
     {otherUnit_maskInput_lo[11407:11392]},
     {otherUnit_maskInput_lo[11391:11376]},
     {otherUnit_maskInput_lo[11375:11360]},
     {otherUnit_maskInput_lo[11359:11344]},
     {otherUnit_maskInput_lo[11343:11328]},
     {otherUnit_maskInput_lo[11327:11312]},
     {otherUnit_maskInput_lo[11311:11296]},
     {otherUnit_maskInput_lo[11295:11280]},
     {otherUnit_maskInput_lo[11279:11264]},
     {otherUnit_maskInput_lo[11263:11248]},
     {otherUnit_maskInput_lo[11247:11232]},
     {otherUnit_maskInput_lo[11231:11216]},
     {otherUnit_maskInput_lo[11215:11200]},
     {otherUnit_maskInput_lo[11199:11184]},
     {otherUnit_maskInput_lo[11183:11168]},
     {otherUnit_maskInput_lo[11167:11152]},
     {otherUnit_maskInput_lo[11151:11136]},
     {otherUnit_maskInput_lo[11135:11120]},
     {otherUnit_maskInput_lo[11119:11104]},
     {otherUnit_maskInput_lo[11103:11088]},
     {otherUnit_maskInput_lo[11087:11072]},
     {otherUnit_maskInput_lo[11071:11056]},
     {otherUnit_maskInput_lo[11055:11040]},
     {otherUnit_maskInput_lo[11039:11024]},
     {otherUnit_maskInput_lo[11023:11008]},
     {otherUnit_maskInput_lo[11007:10992]},
     {otherUnit_maskInput_lo[10991:10976]},
     {otherUnit_maskInput_lo[10975:10960]},
     {otherUnit_maskInput_lo[10959:10944]},
     {otherUnit_maskInput_lo[10943:10928]},
     {otherUnit_maskInput_lo[10927:10912]},
     {otherUnit_maskInput_lo[10911:10896]},
     {otherUnit_maskInput_lo[10895:10880]},
     {otherUnit_maskInput_lo[10879:10864]},
     {otherUnit_maskInput_lo[10863:10848]},
     {otherUnit_maskInput_lo[10847:10832]},
     {otherUnit_maskInput_lo[10831:10816]},
     {otherUnit_maskInput_lo[10815:10800]},
     {otherUnit_maskInput_lo[10799:10784]},
     {otherUnit_maskInput_lo[10783:10768]},
     {otherUnit_maskInput_lo[10767:10752]},
     {otherUnit_maskInput_lo[10751:10736]},
     {otherUnit_maskInput_lo[10735:10720]},
     {otherUnit_maskInput_lo[10719:10704]},
     {otherUnit_maskInput_lo[10703:10688]},
     {otherUnit_maskInput_lo[10687:10672]},
     {otherUnit_maskInput_lo[10671:10656]},
     {otherUnit_maskInput_lo[10655:10640]},
     {otherUnit_maskInput_lo[10639:10624]},
     {otherUnit_maskInput_lo[10623:10608]},
     {otherUnit_maskInput_lo[10607:10592]},
     {otherUnit_maskInput_lo[10591:10576]},
     {otherUnit_maskInput_lo[10575:10560]},
     {otherUnit_maskInput_lo[10559:10544]},
     {otherUnit_maskInput_lo[10543:10528]},
     {otherUnit_maskInput_lo[10527:10512]},
     {otherUnit_maskInput_lo[10511:10496]},
     {otherUnit_maskInput_lo[10495:10480]},
     {otherUnit_maskInput_lo[10479:10464]},
     {otherUnit_maskInput_lo[10463:10448]},
     {otherUnit_maskInput_lo[10447:10432]},
     {otherUnit_maskInput_lo[10431:10416]},
     {otherUnit_maskInput_lo[10415:10400]},
     {otherUnit_maskInput_lo[10399:10384]},
     {otherUnit_maskInput_lo[10383:10368]},
     {otherUnit_maskInput_lo[10367:10352]},
     {otherUnit_maskInput_lo[10351:10336]},
     {otherUnit_maskInput_lo[10335:10320]},
     {otherUnit_maskInput_lo[10319:10304]},
     {otherUnit_maskInput_lo[10303:10288]},
     {otherUnit_maskInput_lo[10287:10272]},
     {otherUnit_maskInput_lo[10271:10256]},
     {otherUnit_maskInput_lo[10255:10240]},
     {otherUnit_maskInput_lo[10239:10224]},
     {otherUnit_maskInput_lo[10223:10208]},
     {otherUnit_maskInput_lo[10207:10192]},
     {otherUnit_maskInput_lo[10191:10176]},
     {otherUnit_maskInput_lo[10175:10160]},
     {otherUnit_maskInput_lo[10159:10144]},
     {otherUnit_maskInput_lo[10143:10128]},
     {otherUnit_maskInput_lo[10127:10112]},
     {otherUnit_maskInput_lo[10111:10096]},
     {otherUnit_maskInput_lo[10095:10080]},
     {otherUnit_maskInput_lo[10079:10064]},
     {otherUnit_maskInput_lo[10063:10048]},
     {otherUnit_maskInput_lo[10047:10032]},
     {otherUnit_maskInput_lo[10031:10016]},
     {otherUnit_maskInput_lo[10015:10000]},
     {otherUnit_maskInput_lo[9999:9984]},
     {otherUnit_maskInput_lo[9983:9968]},
     {otherUnit_maskInput_lo[9967:9952]},
     {otherUnit_maskInput_lo[9951:9936]},
     {otherUnit_maskInput_lo[9935:9920]},
     {otherUnit_maskInput_lo[9919:9904]},
     {otherUnit_maskInput_lo[9903:9888]},
     {otherUnit_maskInput_lo[9887:9872]},
     {otherUnit_maskInput_lo[9871:9856]},
     {otherUnit_maskInput_lo[9855:9840]},
     {otherUnit_maskInput_lo[9839:9824]},
     {otherUnit_maskInput_lo[9823:9808]},
     {otherUnit_maskInput_lo[9807:9792]},
     {otherUnit_maskInput_lo[9791:9776]},
     {otherUnit_maskInput_lo[9775:9760]},
     {otherUnit_maskInput_lo[9759:9744]},
     {otherUnit_maskInput_lo[9743:9728]},
     {otherUnit_maskInput_lo[9727:9712]},
     {otherUnit_maskInput_lo[9711:9696]},
     {otherUnit_maskInput_lo[9695:9680]},
     {otherUnit_maskInput_lo[9679:9664]},
     {otherUnit_maskInput_lo[9663:9648]},
     {otherUnit_maskInput_lo[9647:9632]},
     {otherUnit_maskInput_lo[9631:9616]},
     {otherUnit_maskInput_lo[9615:9600]},
     {otherUnit_maskInput_lo[9599:9584]},
     {otherUnit_maskInput_lo[9583:9568]},
     {otherUnit_maskInput_lo[9567:9552]},
     {otherUnit_maskInput_lo[9551:9536]},
     {otherUnit_maskInput_lo[9535:9520]},
     {otherUnit_maskInput_lo[9519:9504]},
     {otherUnit_maskInput_lo[9503:9488]},
     {otherUnit_maskInput_lo[9487:9472]},
     {otherUnit_maskInput_lo[9471:9456]},
     {otherUnit_maskInput_lo[9455:9440]},
     {otherUnit_maskInput_lo[9439:9424]},
     {otherUnit_maskInput_lo[9423:9408]},
     {otherUnit_maskInput_lo[9407:9392]},
     {otherUnit_maskInput_lo[9391:9376]},
     {otherUnit_maskInput_lo[9375:9360]},
     {otherUnit_maskInput_lo[9359:9344]},
     {otherUnit_maskInput_lo[9343:9328]},
     {otherUnit_maskInput_lo[9327:9312]},
     {otherUnit_maskInput_lo[9311:9296]},
     {otherUnit_maskInput_lo[9295:9280]},
     {otherUnit_maskInput_lo[9279:9264]},
     {otherUnit_maskInput_lo[9263:9248]},
     {otherUnit_maskInput_lo[9247:9232]},
     {otherUnit_maskInput_lo[9231:9216]},
     {otherUnit_maskInput_lo[9215:9200]},
     {otherUnit_maskInput_lo[9199:9184]},
     {otherUnit_maskInput_lo[9183:9168]},
     {otherUnit_maskInput_lo[9167:9152]},
     {otherUnit_maskInput_lo[9151:9136]},
     {otherUnit_maskInput_lo[9135:9120]},
     {otherUnit_maskInput_lo[9119:9104]},
     {otherUnit_maskInput_lo[9103:9088]},
     {otherUnit_maskInput_lo[9087:9072]},
     {otherUnit_maskInput_lo[9071:9056]},
     {otherUnit_maskInput_lo[9055:9040]},
     {otherUnit_maskInput_lo[9039:9024]},
     {otherUnit_maskInput_lo[9023:9008]},
     {otherUnit_maskInput_lo[9007:8992]},
     {otherUnit_maskInput_lo[8991:8976]},
     {otherUnit_maskInput_lo[8975:8960]},
     {otherUnit_maskInput_lo[8959:8944]},
     {otherUnit_maskInput_lo[8943:8928]},
     {otherUnit_maskInput_lo[8927:8912]},
     {otherUnit_maskInput_lo[8911:8896]},
     {otherUnit_maskInput_lo[8895:8880]},
     {otherUnit_maskInput_lo[8879:8864]},
     {otherUnit_maskInput_lo[8863:8848]},
     {otherUnit_maskInput_lo[8847:8832]},
     {otherUnit_maskInput_lo[8831:8816]},
     {otherUnit_maskInput_lo[8815:8800]},
     {otherUnit_maskInput_lo[8799:8784]},
     {otherUnit_maskInput_lo[8783:8768]},
     {otherUnit_maskInput_lo[8767:8752]},
     {otherUnit_maskInput_lo[8751:8736]},
     {otherUnit_maskInput_lo[8735:8720]},
     {otherUnit_maskInput_lo[8719:8704]},
     {otherUnit_maskInput_lo[8703:8688]},
     {otherUnit_maskInput_lo[8687:8672]},
     {otherUnit_maskInput_lo[8671:8656]},
     {otherUnit_maskInput_lo[8655:8640]},
     {otherUnit_maskInput_lo[8639:8624]},
     {otherUnit_maskInput_lo[8623:8608]},
     {otherUnit_maskInput_lo[8607:8592]},
     {otherUnit_maskInput_lo[8591:8576]},
     {otherUnit_maskInput_lo[8575:8560]},
     {otherUnit_maskInput_lo[8559:8544]},
     {otherUnit_maskInput_lo[8543:8528]},
     {otherUnit_maskInput_lo[8527:8512]},
     {otherUnit_maskInput_lo[8511:8496]},
     {otherUnit_maskInput_lo[8495:8480]},
     {otherUnit_maskInput_lo[8479:8464]},
     {otherUnit_maskInput_lo[8463:8448]},
     {otherUnit_maskInput_lo[8447:8432]},
     {otherUnit_maskInput_lo[8431:8416]},
     {otherUnit_maskInput_lo[8415:8400]},
     {otherUnit_maskInput_lo[8399:8384]},
     {otherUnit_maskInput_lo[8383:8368]},
     {otherUnit_maskInput_lo[8367:8352]},
     {otherUnit_maskInput_lo[8351:8336]},
     {otherUnit_maskInput_lo[8335:8320]},
     {otherUnit_maskInput_lo[8319:8304]},
     {otherUnit_maskInput_lo[8303:8288]},
     {otherUnit_maskInput_lo[8287:8272]},
     {otherUnit_maskInput_lo[8271:8256]},
     {otherUnit_maskInput_lo[8255:8240]},
     {otherUnit_maskInput_lo[8239:8224]},
     {otherUnit_maskInput_lo[8223:8208]},
     {otherUnit_maskInput_lo[8207:8192]},
     {otherUnit_maskInput_lo[8191:8176]},
     {otherUnit_maskInput_lo[8175:8160]},
     {otherUnit_maskInput_lo[8159:8144]},
     {otherUnit_maskInput_lo[8143:8128]},
     {otherUnit_maskInput_lo[8127:8112]},
     {otherUnit_maskInput_lo[8111:8096]},
     {otherUnit_maskInput_lo[8095:8080]},
     {otherUnit_maskInput_lo[8079:8064]},
     {otherUnit_maskInput_lo[8063:8048]},
     {otherUnit_maskInput_lo[8047:8032]},
     {otherUnit_maskInput_lo[8031:8016]},
     {otherUnit_maskInput_lo[8015:8000]},
     {otherUnit_maskInput_lo[7999:7984]},
     {otherUnit_maskInput_lo[7983:7968]},
     {otherUnit_maskInput_lo[7967:7952]},
     {otherUnit_maskInput_lo[7951:7936]},
     {otherUnit_maskInput_lo[7935:7920]},
     {otherUnit_maskInput_lo[7919:7904]},
     {otherUnit_maskInput_lo[7903:7888]},
     {otherUnit_maskInput_lo[7887:7872]},
     {otherUnit_maskInput_lo[7871:7856]},
     {otherUnit_maskInput_lo[7855:7840]},
     {otherUnit_maskInput_lo[7839:7824]},
     {otherUnit_maskInput_lo[7823:7808]},
     {otherUnit_maskInput_lo[7807:7792]},
     {otherUnit_maskInput_lo[7791:7776]},
     {otherUnit_maskInput_lo[7775:7760]},
     {otherUnit_maskInput_lo[7759:7744]},
     {otherUnit_maskInput_lo[7743:7728]},
     {otherUnit_maskInput_lo[7727:7712]},
     {otherUnit_maskInput_lo[7711:7696]},
     {otherUnit_maskInput_lo[7695:7680]},
     {otherUnit_maskInput_lo[7679:7664]},
     {otherUnit_maskInput_lo[7663:7648]},
     {otherUnit_maskInput_lo[7647:7632]},
     {otherUnit_maskInput_lo[7631:7616]},
     {otherUnit_maskInput_lo[7615:7600]},
     {otherUnit_maskInput_lo[7599:7584]},
     {otherUnit_maskInput_lo[7583:7568]},
     {otherUnit_maskInput_lo[7567:7552]},
     {otherUnit_maskInput_lo[7551:7536]},
     {otherUnit_maskInput_lo[7535:7520]},
     {otherUnit_maskInput_lo[7519:7504]},
     {otherUnit_maskInput_lo[7503:7488]},
     {otherUnit_maskInput_lo[7487:7472]},
     {otherUnit_maskInput_lo[7471:7456]},
     {otherUnit_maskInput_lo[7455:7440]},
     {otherUnit_maskInput_lo[7439:7424]},
     {otherUnit_maskInput_lo[7423:7408]},
     {otherUnit_maskInput_lo[7407:7392]},
     {otherUnit_maskInput_lo[7391:7376]},
     {otherUnit_maskInput_lo[7375:7360]},
     {otherUnit_maskInput_lo[7359:7344]},
     {otherUnit_maskInput_lo[7343:7328]},
     {otherUnit_maskInput_lo[7327:7312]},
     {otherUnit_maskInput_lo[7311:7296]},
     {otherUnit_maskInput_lo[7295:7280]},
     {otherUnit_maskInput_lo[7279:7264]},
     {otherUnit_maskInput_lo[7263:7248]},
     {otherUnit_maskInput_lo[7247:7232]},
     {otherUnit_maskInput_lo[7231:7216]},
     {otherUnit_maskInput_lo[7215:7200]},
     {otherUnit_maskInput_lo[7199:7184]},
     {otherUnit_maskInput_lo[7183:7168]},
     {otherUnit_maskInput_lo[7167:7152]},
     {otherUnit_maskInput_lo[7151:7136]},
     {otherUnit_maskInput_lo[7135:7120]},
     {otherUnit_maskInput_lo[7119:7104]},
     {otherUnit_maskInput_lo[7103:7088]},
     {otherUnit_maskInput_lo[7087:7072]},
     {otherUnit_maskInput_lo[7071:7056]},
     {otherUnit_maskInput_lo[7055:7040]},
     {otherUnit_maskInput_lo[7039:7024]},
     {otherUnit_maskInput_lo[7023:7008]},
     {otherUnit_maskInput_lo[7007:6992]},
     {otherUnit_maskInput_lo[6991:6976]},
     {otherUnit_maskInput_lo[6975:6960]},
     {otherUnit_maskInput_lo[6959:6944]},
     {otherUnit_maskInput_lo[6943:6928]},
     {otherUnit_maskInput_lo[6927:6912]},
     {otherUnit_maskInput_lo[6911:6896]},
     {otherUnit_maskInput_lo[6895:6880]},
     {otherUnit_maskInput_lo[6879:6864]},
     {otherUnit_maskInput_lo[6863:6848]},
     {otherUnit_maskInput_lo[6847:6832]},
     {otherUnit_maskInput_lo[6831:6816]},
     {otherUnit_maskInput_lo[6815:6800]},
     {otherUnit_maskInput_lo[6799:6784]},
     {otherUnit_maskInput_lo[6783:6768]},
     {otherUnit_maskInput_lo[6767:6752]},
     {otherUnit_maskInput_lo[6751:6736]},
     {otherUnit_maskInput_lo[6735:6720]},
     {otherUnit_maskInput_lo[6719:6704]},
     {otherUnit_maskInput_lo[6703:6688]},
     {otherUnit_maskInput_lo[6687:6672]},
     {otherUnit_maskInput_lo[6671:6656]},
     {otherUnit_maskInput_lo[6655:6640]},
     {otherUnit_maskInput_lo[6639:6624]},
     {otherUnit_maskInput_lo[6623:6608]},
     {otherUnit_maskInput_lo[6607:6592]},
     {otherUnit_maskInput_lo[6591:6576]},
     {otherUnit_maskInput_lo[6575:6560]},
     {otherUnit_maskInput_lo[6559:6544]},
     {otherUnit_maskInput_lo[6543:6528]},
     {otherUnit_maskInput_lo[6527:6512]},
     {otherUnit_maskInput_lo[6511:6496]},
     {otherUnit_maskInput_lo[6495:6480]},
     {otherUnit_maskInput_lo[6479:6464]},
     {otherUnit_maskInput_lo[6463:6448]},
     {otherUnit_maskInput_lo[6447:6432]},
     {otherUnit_maskInput_lo[6431:6416]},
     {otherUnit_maskInput_lo[6415:6400]},
     {otherUnit_maskInput_lo[6399:6384]},
     {otherUnit_maskInput_lo[6383:6368]},
     {otherUnit_maskInput_lo[6367:6352]},
     {otherUnit_maskInput_lo[6351:6336]},
     {otherUnit_maskInput_lo[6335:6320]},
     {otherUnit_maskInput_lo[6319:6304]},
     {otherUnit_maskInput_lo[6303:6288]},
     {otherUnit_maskInput_lo[6287:6272]},
     {otherUnit_maskInput_lo[6271:6256]},
     {otherUnit_maskInput_lo[6255:6240]},
     {otherUnit_maskInput_lo[6239:6224]},
     {otherUnit_maskInput_lo[6223:6208]},
     {otherUnit_maskInput_lo[6207:6192]},
     {otherUnit_maskInput_lo[6191:6176]},
     {otherUnit_maskInput_lo[6175:6160]},
     {otherUnit_maskInput_lo[6159:6144]},
     {otherUnit_maskInput_lo[6143:6128]},
     {otherUnit_maskInput_lo[6127:6112]},
     {otherUnit_maskInput_lo[6111:6096]},
     {otherUnit_maskInput_lo[6095:6080]},
     {otherUnit_maskInput_lo[6079:6064]},
     {otherUnit_maskInput_lo[6063:6048]},
     {otherUnit_maskInput_lo[6047:6032]},
     {otherUnit_maskInput_lo[6031:6016]},
     {otherUnit_maskInput_lo[6015:6000]},
     {otherUnit_maskInput_lo[5999:5984]},
     {otherUnit_maskInput_lo[5983:5968]},
     {otherUnit_maskInput_lo[5967:5952]},
     {otherUnit_maskInput_lo[5951:5936]},
     {otherUnit_maskInput_lo[5935:5920]},
     {otherUnit_maskInput_lo[5919:5904]},
     {otherUnit_maskInput_lo[5903:5888]},
     {otherUnit_maskInput_lo[5887:5872]},
     {otherUnit_maskInput_lo[5871:5856]},
     {otherUnit_maskInput_lo[5855:5840]},
     {otherUnit_maskInput_lo[5839:5824]},
     {otherUnit_maskInput_lo[5823:5808]},
     {otherUnit_maskInput_lo[5807:5792]},
     {otherUnit_maskInput_lo[5791:5776]},
     {otherUnit_maskInput_lo[5775:5760]},
     {otherUnit_maskInput_lo[5759:5744]},
     {otherUnit_maskInput_lo[5743:5728]},
     {otherUnit_maskInput_lo[5727:5712]},
     {otherUnit_maskInput_lo[5711:5696]},
     {otherUnit_maskInput_lo[5695:5680]},
     {otherUnit_maskInput_lo[5679:5664]},
     {otherUnit_maskInput_lo[5663:5648]},
     {otherUnit_maskInput_lo[5647:5632]},
     {otherUnit_maskInput_lo[5631:5616]},
     {otherUnit_maskInput_lo[5615:5600]},
     {otherUnit_maskInput_lo[5599:5584]},
     {otherUnit_maskInput_lo[5583:5568]},
     {otherUnit_maskInput_lo[5567:5552]},
     {otherUnit_maskInput_lo[5551:5536]},
     {otherUnit_maskInput_lo[5535:5520]},
     {otherUnit_maskInput_lo[5519:5504]},
     {otherUnit_maskInput_lo[5503:5488]},
     {otherUnit_maskInput_lo[5487:5472]},
     {otherUnit_maskInput_lo[5471:5456]},
     {otherUnit_maskInput_lo[5455:5440]},
     {otherUnit_maskInput_lo[5439:5424]},
     {otherUnit_maskInput_lo[5423:5408]},
     {otherUnit_maskInput_lo[5407:5392]},
     {otherUnit_maskInput_lo[5391:5376]},
     {otherUnit_maskInput_lo[5375:5360]},
     {otherUnit_maskInput_lo[5359:5344]},
     {otherUnit_maskInput_lo[5343:5328]},
     {otherUnit_maskInput_lo[5327:5312]},
     {otherUnit_maskInput_lo[5311:5296]},
     {otherUnit_maskInput_lo[5295:5280]},
     {otherUnit_maskInput_lo[5279:5264]},
     {otherUnit_maskInput_lo[5263:5248]},
     {otherUnit_maskInput_lo[5247:5232]},
     {otherUnit_maskInput_lo[5231:5216]},
     {otherUnit_maskInput_lo[5215:5200]},
     {otherUnit_maskInput_lo[5199:5184]},
     {otherUnit_maskInput_lo[5183:5168]},
     {otherUnit_maskInput_lo[5167:5152]},
     {otherUnit_maskInput_lo[5151:5136]},
     {otherUnit_maskInput_lo[5135:5120]},
     {otherUnit_maskInput_lo[5119:5104]},
     {otherUnit_maskInput_lo[5103:5088]},
     {otherUnit_maskInput_lo[5087:5072]},
     {otherUnit_maskInput_lo[5071:5056]},
     {otherUnit_maskInput_lo[5055:5040]},
     {otherUnit_maskInput_lo[5039:5024]},
     {otherUnit_maskInput_lo[5023:5008]},
     {otherUnit_maskInput_lo[5007:4992]},
     {otherUnit_maskInput_lo[4991:4976]},
     {otherUnit_maskInput_lo[4975:4960]},
     {otherUnit_maskInput_lo[4959:4944]},
     {otherUnit_maskInput_lo[4943:4928]},
     {otherUnit_maskInput_lo[4927:4912]},
     {otherUnit_maskInput_lo[4911:4896]},
     {otherUnit_maskInput_lo[4895:4880]},
     {otherUnit_maskInput_lo[4879:4864]},
     {otherUnit_maskInput_lo[4863:4848]},
     {otherUnit_maskInput_lo[4847:4832]},
     {otherUnit_maskInput_lo[4831:4816]},
     {otherUnit_maskInput_lo[4815:4800]},
     {otherUnit_maskInput_lo[4799:4784]},
     {otherUnit_maskInput_lo[4783:4768]},
     {otherUnit_maskInput_lo[4767:4752]},
     {otherUnit_maskInput_lo[4751:4736]},
     {otherUnit_maskInput_lo[4735:4720]},
     {otherUnit_maskInput_lo[4719:4704]},
     {otherUnit_maskInput_lo[4703:4688]},
     {otherUnit_maskInput_lo[4687:4672]},
     {otherUnit_maskInput_lo[4671:4656]},
     {otherUnit_maskInput_lo[4655:4640]},
     {otherUnit_maskInput_lo[4639:4624]},
     {otherUnit_maskInput_lo[4623:4608]},
     {otherUnit_maskInput_lo[4607:4592]},
     {otherUnit_maskInput_lo[4591:4576]},
     {otherUnit_maskInput_lo[4575:4560]},
     {otherUnit_maskInput_lo[4559:4544]},
     {otherUnit_maskInput_lo[4543:4528]},
     {otherUnit_maskInput_lo[4527:4512]},
     {otherUnit_maskInput_lo[4511:4496]},
     {otherUnit_maskInput_lo[4495:4480]},
     {otherUnit_maskInput_lo[4479:4464]},
     {otherUnit_maskInput_lo[4463:4448]},
     {otherUnit_maskInput_lo[4447:4432]},
     {otherUnit_maskInput_lo[4431:4416]},
     {otherUnit_maskInput_lo[4415:4400]},
     {otherUnit_maskInput_lo[4399:4384]},
     {otherUnit_maskInput_lo[4383:4368]},
     {otherUnit_maskInput_lo[4367:4352]},
     {otherUnit_maskInput_lo[4351:4336]},
     {otherUnit_maskInput_lo[4335:4320]},
     {otherUnit_maskInput_lo[4319:4304]},
     {otherUnit_maskInput_lo[4303:4288]},
     {otherUnit_maskInput_lo[4287:4272]},
     {otherUnit_maskInput_lo[4271:4256]},
     {otherUnit_maskInput_lo[4255:4240]},
     {otherUnit_maskInput_lo[4239:4224]},
     {otherUnit_maskInput_lo[4223:4208]},
     {otherUnit_maskInput_lo[4207:4192]},
     {otherUnit_maskInput_lo[4191:4176]},
     {otherUnit_maskInput_lo[4175:4160]},
     {otherUnit_maskInput_lo[4159:4144]},
     {otherUnit_maskInput_lo[4143:4128]},
     {otherUnit_maskInput_lo[4127:4112]},
     {otherUnit_maskInput_lo[4111:4096]},
     {otherUnit_maskInput_lo[4095:4080]},
     {otherUnit_maskInput_lo[4079:4064]},
     {otherUnit_maskInput_lo[4063:4048]},
     {otherUnit_maskInput_lo[4047:4032]},
     {otherUnit_maskInput_lo[4031:4016]},
     {otherUnit_maskInput_lo[4015:4000]},
     {otherUnit_maskInput_lo[3999:3984]},
     {otherUnit_maskInput_lo[3983:3968]},
     {otherUnit_maskInput_lo[3967:3952]},
     {otherUnit_maskInput_lo[3951:3936]},
     {otherUnit_maskInput_lo[3935:3920]},
     {otherUnit_maskInput_lo[3919:3904]},
     {otherUnit_maskInput_lo[3903:3888]},
     {otherUnit_maskInput_lo[3887:3872]},
     {otherUnit_maskInput_lo[3871:3856]},
     {otherUnit_maskInput_lo[3855:3840]},
     {otherUnit_maskInput_lo[3839:3824]},
     {otherUnit_maskInput_lo[3823:3808]},
     {otherUnit_maskInput_lo[3807:3792]},
     {otherUnit_maskInput_lo[3791:3776]},
     {otherUnit_maskInput_lo[3775:3760]},
     {otherUnit_maskInput_lo[3759:3744]},
     {otherUnit_maskInput_lo[3743:3728]},
     {otherUnit_maskInput_lo[3727:3712]},
     {otherUnit_maskInput_lo[3711:3696]},
     {otherUnit_maskInput_lo[3695:3680]},
     {otherUnit_maskInput_lo[3679:3664]},
     {otherUnit_maskInput_lo[3663:3648]},
     {otherUnit_maskInput_lo[3647:3632]},
     {otherUnit_maskInput_lo[3631:3616]},
     {otherUnit_maskInput_lo[3615:3600]},
     {otherUnit_maskInput_lo[3599:3584]},
     {otherUnit_maskInput_lo[3583:3568]},
     {otherUnit_maskInput_lo[3567:3552]},
     {otherUnit_maskInput_lo[3551:3536]},
     {otherUnit_maskInput_lo[3535:3520]},
     {otherUnit_maskInput_lo[3519:3504]},
     {otherUnit_maskInput_lo[3503:3488]},
     {otherUnit_maskInput_lo[3487:3472]},
     {otherUnit_maskInput_lo[3471:3456]},
     {otherUnit_maskInput_lo[3455:3440]},
     {otherUnit_maskInput_lo[3439:3424]},
     {otherUnit_maskInput_lo[3423:3408]},
     {otherUnit_maskInput_lo[3407:3392]},
     {otherUnit_maskInput_lo[3391:3376]},
     {otherUnit_maskInput_lo[3375:3360]},
     {otherUnit_maskInput_lo[3359:3344]},
     {otherUnit_maskInput_lo[3343:3328]},
     {otherUnit_maskInput_lo[3327:3312]},
     {otherUnit_maskInput_lo[3311:3296]},
     {otherUnit_maskInput_lo[3295:3280]},
     {otherUnit_maskInput_lo[3279:3264]},
     {otherUnit_maskInput_lo[3263:3248]},
     {otherUnit_maskInput_lo[3247:3232]},
     {otherUnit_maskInput_lo[3231:3216]},
     {otherUnit_maskInput_lo[3215:3200]},
     {otherUnit_maskInput_lo[3199:3184]},
     {otherUnit_maskInput_lo[3183:3168]},
     {otherUnit_maskInput_lo[3167:3152]},
     {otherUnit_maskInput_lo[3151:3136]},
     {otherUnit_maskInput_lo[3135:3120]},
     {otherUnit_maskInput_lo[3119:3104]},
     {otherUnit_maskInput_lo[3103:3088]},
     {otherUnit_maskInput_lo[3087:3072]},
     {otherUnit_maskInput_lo[3071:3056]},
     {otherUnit_maskInput_lo[3055:3040]},
     {otherUnit_maskInput_lo[3039:3024]},
     {otherUnit_maskInput_lo[3023:3008]},
     {otherUnit_maskInput_lo[3007:2992]},
     {otherUnit_maskInput_lo[2991:2976]},
     {otherUnit_maskInput_lo[2975:2960]},
     {otherUnit_maskInput_lo[2959:2944]},
     {otherUnit_maskInput_lo[2943:2928]},
     {otherUnit_maskInput_lo[2927:2912]},
     {otherUnit_maskInput_lo[2911:2896]},
     {otherUnit_maskInput_lo[2895:2880]},
     {otherUnit_maskInput_lo[2879:2864]},
     {otherUnit_maskInput_lo[2863:2848]},
     {otherUnit_maskInput_lo[2847:2832]},
     {otherUnit_maskInput_lo[2831:2816]},
     {otherUnit_maskInput_lo[2815:2800]},
     {otherUnit_maskInput_lo[2799:2784]},
     {otherUnit_maskInput_lo[2783:2768]},
     {otherUnit_maskInput_lo[2767:2752]},
     {otherUnit_maskInput_lo[2751:2736]},
     {otherUnit_maskInput_lo[2735:2720]},
     {otherUnit_maskInput_lo[2719:2704]},
     {otherUnit_maskInput_lo[2703:2688]},
     {otherUnit_maskInput_lo[2687:2672]},
     {otherUnit_maskInput_lo[2671:2656]},
     {otherUnit_maskInput_lo[2655:2640]},
     {otherUnit_maskInput_lo[2639:2624]},
     {otherUnit_maskInput_lo[2623:2608]},
     {otherUnit_maskInput_lo[2607:2592]},
     {otherUnit_maskInput_lo[2591:2576]},
     {otherUnit_maskInput_lo[2575:2560]},
     {otherUnit_maskInput_lo[2559:2544]},
     {otherUnit_maskInput_lo[2543:2528]},
     {otherUnit_maskInput_lo[2527:2512]},
     {otherUnit_maskInput_lo[2511:2496]},
     {otherUnit_maskInput_lo[2495:2480]},
     {otherUnit_maskInput_lo[2479:2464]},
     {otherUnit_maskInput_lo[2463:2448]},
     {otherUnit_maskInput_lo[2447:2432]},
     {otherUnit_maskInput_lo[2431:2416]},
     {otherUnit_maskInput_lo[2415:2400]},
     {otherUnit_maskInput_lo[2399:2384]},
     {otherUnit_maskInput_lo[2383:2368]},
     {otherUnit_maskInput_lo[2367:2352]},
     {otherUnit_maskInput_lo[2351:2336]},
     {otherUnit_maskInput_lo[2335:2320]},
     {otherUnit_maskInput_lo[2319:2304]},
     {otherUnit_maskInput_lo[2303:2288]},
     {otherUnit_maskInput_lo[2287:2272]},
     {otherUnit_maskInput_lo[2271:2256]},
     {otherUnit_maskInput_lo[2255:2240]},
     {otherUnit_maskInput_lo[2239:2224]},
     {otherUnit_maskInput_lo[2223:2208]},
     {otherUnit_maskInput_lo[2207:2192]},
     {otherUnit_maskInput_lo[2191:2176]},
     {otherUnit_maskInput_lo[2175:2160]},
     {otherUnit_maskInput_lo[2159:2144]},
     {otherUnit_maskInput_lo[2143:2128]},
     {otherUnit_maskInput_lo[2127:2112]},
     {otherUnit_maskInput_lo[2111:2096]},
     {otherUnit_maskInput_lo[2095:2080]},
     {otherUnit_maskInput_lo[2079:2064]},
     {otherUnit_maskInput_lo[2063:2048]},
     {otherUnit_maskInput_lo[2047:2032]},
     {otherUnit_maskInput_lo[2031:2016]},
     {otherUnit_maskInput_lo[2015:2000]},
     {otherUnit_maskInput_lo[1999:1984]},
     {otherUnit_maskInput_lo[1983:1968]},
     {otherUnit_maskInput_lo[1967:1952]},
     {otherUnit_maskInput_lo[1951:1936]},
     {otherUnit_maskInput_lo[1935:1920]},
     {otherUnit_maskInput_lo[1919:1904]},
     {otherUnit_maskInput_lo[1903:1888]},
     {otherUnit_maskInput_lo[1887:1872]},
     {otherUnit_maskInput_lo[1871:1856]},
     {otherUnit_maskInput_lo[1855:1840]},
     {otherUnit_maskInput_lo[1839:1824]},
     {otherUnit_maskInput_lo[1823:1808]},
     {otherUnit_maskInput_lo[1807:1792]},
     {otherUnit_maskInput_lo[1791:1776]},
     {otherUnit_maskInput_lo[1775:1760]},
     {otherUnit_maskInput_lo[1759:1744]},
     {otherUnit_maskInput_lo[1743:1728]},
     {otherUnit_maskInput_lo[1727:1712]},
     {otherUnit_maskInput_lo[1711:1696]},
     {otherUnit_maskInput_lo[1695:1680]},
     {otherUnit_maskInput_lo[1679:1664]},
     {otherUnit_maskInput_lo[1663:1648]},
     {otherUnit_maskInput_lo[1647:1632]},
     {otherUnit_maskInput_lo[1631:1616]},
     {otherUnit_maskInput_lo[1615:1600]},
     {otherUnit_maskInput_lo[1599:1584]},
     {otherUnit_maskInput_lo[1583:1568]},
     {otherUnit_maskInput_lo[1567:1552]},
     {otherUnit_maskInput_lo[1551:1536]},
     {otherUnit_maskInput_lo[1535:1520]},
     {otherUnit_maskInput_lo[1519:1504]},
     {otherUnit_maskInput_lo[1503:1488]},
     {otherUnit_maskInput_lo[1487:1472]},
     {otherUnit_maskInput_lo[1471:1456]},
     {otherUnit_maskInput_lo[1455:1440]},
     {otherUnit_maskInput_lo[1439:1424]},
     {otherUnit_maskInput_lo[1423:1408]},
     {otherUnit_maskInput_lo[1407:1392]},
     {otherUnit_maskInput_lo[1391:1376]},
     {otherUnit_maskInput_lo[1375:1360]},
     {otherUnit_maskInput_lo[1359:1344]},
     {otherUnit_maskInput_lo[1343:1328]},
     {otherUnit_maskInput_lo[1327:1312]},
     {otherUnit_maskInput_lo[1311:1296]},
     {otherUnit_maskInput_lo[1295:1280]},
     {otherUnit_maskInput_lo[1279:1264]},
     {otherUnit_maskInput_lo[1263:1248]},
     {otherUnit_maskInput_lo[1247:1232]},
     {otherUnit_maskInput_lo[1231:1216]},
     {otherUnit_maskInput_lo[1215:1200]},
     {otherUnit_maskInput_lo[1199:1184]},
     {otherUnit_maskInput_lo[1183:1168]},
     {otherUnit_maskInput_lo[1167:1152]},
     {otherUnit_maskInput_lo[1151:1136]},
     {otherUnit_maskInput_lo[1135:1120]},
     {otherUnit_maskInput_lo[1119:1104]},
     {otherUnit_maskInput_lo[1103:1088]},
     {otherUnit_maskInput_lo[1087:1072]},
     {otherUnit_maskInput_lo[1071:1056]},
     {otherUnit_maskInput_lo[1055:1040]},
     {otherUnit_maskInput_lo[1039:1024]},
     {otherUnit_maskInput_lo[1023:1008]},
     {otherUnit_maskInput_lo[1007:992]},
     {otherUnit_maskInput_lo[991:976]},
     {otherUnit_maskInput_lo[975:960]},
     {otherUnit_maskInput_lo[959:944]},
     {otherUnit_maskInput_lo[943:928]},
     {otherUnit_maskInput_lo[927:912]},
     {otherUnit_maskInput_lo[911:896]},
     {otherUnit_maskInput_lo[895:880]},
     {otherUnit_maskInput_lo[879:864]},
     {otherUnit_maskInput_lo[863:848]},
     {otherUnit_maskInput_lo[847:832]},
     {otherUnit_maskInput_lo[831:816]},
     {otherUnit_maskInput_lo[815:800]},
     {otherUnit_maskInput_lo[799:784]},
     {otherUnit_maskInput_lo[783:768]},
     {otherUnit_maskInput_lo[767:752]},
     {otherUnit_maskInput_lo[751:736]},
     {otherUnit_maskInput_lo[735:720]},
     {otherUnit_maskInput_lo[719:704]},
     {otherUnit_maskInput_lo[703:688]},
     {otherUnit_maskInput_lo[687:672]},
     {otherUnit_maskInput_lo[671:656]},
     {otherUnit_maskInput_lo[655:640]},
     {otherUnit_maskInput_lo[639:624]},
     {otherUnit_maskInput_lo[623:608]},
     {otherUnit_maskInput_lo[607:592]},
     {otherUnit_maskInput_lo[591:576]},
     {otherUnit_maskInput_lo[575:560]},
     {otherUnit_maskInput_lo[559:544]},
     {otherUnit_maskInput_lo[543:528]},
     {otherUnit_maskInput_lo[527:512]},
     {otherUnit_maskInput_lo[511:496]},
     {otherUnit_maskInput_lo[495:480]},
     {otherUnit_maskInput_lo[479:464]},
     {otherUnit_maskInput_lo[463:448]},
     {otherUnit_maskInput_lo[447:432]},
     {otherUnit_maskInput_lo[431:416]},
     {otherUnit_maskInput_lo[415:400]},
     {otherUnit_maskInput_lo[399:384]},
     {otherUnit_maskInput_lo[383:368]},
     {otherUnit_maskInput_lo[367:352]},
     {otherUnit_maskInput_lo[351:336]},
     {otherUnit_maskInput_lo[335:320]},
     {otherUnit_maskInput_lo[319:304]},
     {otherUnit_maskInput_lo[303:288]},
     {otherUnit_maskInput_lo[287:272]},
     {otherUnit_maskInput_lo[271:256]},
     {otherUnit_maskInput_lo[255:240]},
     {otherUnit_maskInput_lo[239:224]},
     {otherUnit_maskInput_lo[223:208]},
     {otherUnit_maskInput_lo[207:192]},
     {otherUnit_maskInput_lo[191:176]},
     {otherUnit_maskInput_lo[175:160]},
     {otherUnit_maskInput_lo[159:144]},
     {otherUnit_maskInput_lo[143:128]},
     {otherUnit_maskInput_lo[127:112]},
     {otherUnit_maskInput_lo[111:96]},
     {otherUnit_maskInput_lo[95:80]},
     {otherUnit_maskInput_lo[79:64]},
     {otherUnit_maskInput_lo[63:48]},
     {otherUnit_maskInput_lo[47:32]},
     {otherUnit_maskInput_lo[31:16]},
     {otherUnit_maskInput_lo[15:0]}};
  wire                vrfWritePort_0_valid_0 = writeQueueVec_0_deq_valid;
  wire [4:0]          vrfWritePort_0_bits_vd_0 = writeQueueVec_0_deq_bits_data_vd;
  wire [8:0]          vrfWritePort_0_bits_offset_0 = writeQueueVec_0_deq_bits_data_offset;
  wire [3:0]          vrfWritePort_0_bits_mask_0 = writeQueueVec_0_deq_bits_data_mask;
  wire [31:0]         vrfWritePort_0_bits_data_0 = writeQueueVec_0_deq_bits_data_data;
  wire                vrfWritePort_0_bits_last_0 = writeQueueVec_0_deq_bits_data_last;
  wire [2:0]          vrfWritePort_0_bits_instructionIndex_0 = writeQueueVec_0_deq_bits_data_instructionIndex;
  wire [2:0]          writeIndexQueue_enq_bits = writeQueueVec_0_deq_bits_data_instructionIndex;
  wire [31:0]         writeQueueVec_0_enq_bits_data_data;
  wire                writeQueueVec_0_enq_bits_data_last;
  wire [32:0]         writeQueueVec_dataIn_lo_hi = {writeQueueVec_0_enq_bits_data_data, writeQueueVec_0_enq_bits_data_last};
  wire [2:0]          writeQueueVec_0_enq_bits_data_instructionIndex;
  wire [35:0]         writeQueueVec_dataIn_lo = {writeQueueVec_dataIn_lo_hi, writeQueueVec_0_enq_bits_data_instructionIndex};
  wire [4:0]          writeQueueVec_0_enq_bits_data_vd;
  wire [8:0]          writeQueueVec_0_enq_bits_data_offset;
  wire [13:0]         writeQueueVec_dataIn_hi_hi = {writeQueueVec_0_enq_bits_data_vd, writeQueueVec_0_enq_bits_data_offset};
  wire [3:0]          writeQueueVec_0_enq_bits_data_mask;
  wire [17:0]         writeQueueVec_dataIn_hi = {writeQueueVec_dataIn_hi_hi, writeQueueVec_0_enq_bits_data_mask};
  wire [57:0]         writeQueueVec_dataIn = {writeQueueVec_dataIn_hi, writeQueueVec_dataIn_lo, 4'h1};
  wire [3:0]          writeQueueVec_dataOut_targetLane = _writeQueueVec_fifo_data_out[3:0];
  wire [2:0]          writeQueueVec_dataOut_data_instructionIndex = _writeQueueVec_fifo_data_out[6:4];
  wire                writeQueueVec_dataOut_data_last = _writeQueueVec_fifo_data_out[7];
  wire [31:0]         writeQueueVec_dataOut_data_data = _writeQueueVec_fifo_data_out[39:8];
  wire [3:0]          writeQueueVec_dataOut_data_mask = _writeQueueVec_fifo_data_out[43:40];
  wire [8:0]          writeQueueVec_dataOut_data_offset = _writeQueueVec_fifo_data_out[52:44];
  wire [4:0]          writeQueueVec_dataOut_data_vd = _writeQueueVec_fifo_data_out[57:53];
  wire                writeQueueVec_0_enq_ready = ~_writeQueueVec_fifo_full;
  wire                writeQueueVec_0_enq_valid;
  wire                _probeWire_slots_0_writeValid_T = writeQueueVec_0_enq_ready & writeQueueVec_0_enq_valid;
  assign writeQueueVec_0_deq_valid = ~_writeQueueVec_fifo_empty | writeQueueVec_0_enq_valid;
  assign writeQueueVec_0_deq_bits_data_vd = _writeQueueVec_fifo_empty ? writeQueueVec_0_enq_bits_data_vd : writeQueueVec_dataOut_data_vd;
  assign writeQueueVec_0_deq_bits_data_offset = _writeQueueVec_fifo_empty ? writeQueueVec_0_enq_bits_data_offset : writeQueueVec_dataOut_data_offset;
  assign writeQueueVec_0_deq_bits_data_mask = _writeQueueVec_fifo_empty ? writeQueueVec_0_enq_bits_data_mask : writeQueueVec_dataOut_data_mask;
  assign writeQueueVec_0_deq_bits_data_data = _writeQueueVec_fifo_empty ? writeQueueVec_0_enq_bits_data_data : writeQueueVec_dataOut_data_data;
  assign writeQueueVec_0_deq_bits_data_last = _writeQueueVec_fifo_empty ? writeQueueVec_0_enq_bits_data_last : writeQueueVec_dataOut_data_last;
  assign writeQueueVec_0_deq_bits_data_instructionIndex = _writeQueueVec_fifo_empty ? writeQueueVec_0_enq_bits_data_instructionIndex : writeQueueVec_dataOut_data_instructionIndex;
  wire [3:0]          writeQueueVec_0_deq_bits_targetLane = _writeQueueVec_fifo_empty ? 4'h1 : writeQueueVec_dataOut_targetLane;
  wire                vrfWritePort_1_valid_0 = writeQueueVec_1_deq_valid;
  wire [4:0]          vrfWritePort_1_bits_vd_0 = writeQueueVec_1_deq_bits_data_vd;
  wire [8:0]          vrfWritePort_1_bits_offset_0 = writeQueueVec_1_deq_bits_data_offset;
  wire [3:0]          vrfWritePort_1_bits_mask_0 = writeQueueVec_1_deq_bits_data_mask;
  wire [31:0]         vrfWritePort_1_bits_data_0 = writeQueueVec_1_deq_bits_data_data;
  wire                vrfWritePort_1_bits_last_0 = writeQueueVec_1_deq_bits_data_last;
  wire [2:0]          vrfWritePort_1_bits_instructionIndex_0 = writeQueueVec_1_deq_bits_data_instructionIndex;
  wire [2:0]          writeIndexQueue_1_enq_bits = writeQueueVec_1_deq_bits_data_instructionIndex;
  wire [31:0]         writeQueueVec_1_enq_bits_data_data;
  wire                writeQueueVec_1_enq_bits_data_last;
  wire [32:0]         writeQueueVec_dataIn_lo_hi_1 = {writeQueueVec_1_enq_bits_data_data, writeQueueVec_1_enq_bits_data_last};
  wire [2:0]          writeQueueVec_1_enq_bits_data_instructionIndex;
  wire [35:0]         writeQueueVec_dataIn_lo_1 = {writeQueueVec_dataIn_lo_hi_1, writeQueueVec_1_enq_bits_data_instructionIndex};
  wire [4:0]          writeQueueVec_1_enq_bits_data_vd;
  wire [8:0]          writeQueueVec_1_enq_bits_data_offset;
  wire [13:0]         writeQueueVec_dataIn_hi_hi_1 = {writeQueueVec_1_enq_bits_data_vd, writeQueueVec_1_enq_bits_data_offset};
  wire [3:0]          writeQueueVec_1_enq_bits_data_mask;
  wire [17:0]         writeQueueVec_dataIn_hi_1 = {writeQueueVec_dataIn_hi_hi_1, writeQueueVec_1_enq_bits_data_mask};
  wire [57:0]         writeQueueVec_dataIn_1 = {writeQueueVec_dataIn_hi_1, writeQueueVec_dataIn_lo_1, 4'h2};
  wire [3:0]          writeQueueVec_dataOut_1_targetLane = _writeQueueVec_fifo_1_data_out[3:0];
  wire [2:0]          writeQueueVec_dataOut_1_data_instructionIndex = _writeQueueVec_fifo_1_data_out[6:4];
  wire                writeQueueVec_dataOut_1_data_last = _writeQueueVec_fifo_1_data_out[7];
  wire [31:0]         writeQueueVec_dataOut_1_data_data = _writeQueueVec_fifo_1_data_out[39:8];
  wire [3:0]          writeQueueVec_dataOut_1_data_mask = _writeQueueVec_fifo_1_data_out[43:40];
  wire [8:0]          writeQueueVec_dataOut_1_data_offset = _writeQueueVec_fifo_1_data_out[52:44];
  wire [4:0]          writeQueueVec_dataOut_1_data_vd = _writeQueueVec_fifo_1_data_out[57:53];
  wire                writeQueueVec_1_enq_ready = ~_writeQueueVec_fifo_1_full;
  wire                writeQueueVec_1_enq_valid;
  wire                _probeWire_slots_1_writeValid_T = writeQueueVec_1_enq_ready & writeQueueVec_1_enq_valid;
  assign writeQueueVec_1_deq_valid = ~_writeQueueVec_fifo_1_empty | writeQueueVec_1_enq_valid;
  assign writeQueueVec_1_deq_bits_data_vd = _writeQueueVec_fifo_1_empty ? writeQueueVec_1_enq_bits_data_vd : writeQueueVec_dataOut_1_data_vd;
  assign writeQueueVec_1_deq_bits_data_offset = _writeQueueVec_fifo_1_empty ? writeQueueVec_1_enq_bits_data_offset : writeQueueVec_dataOut_1_data_offset;
  assign writeQueueVec_1_deq_bits_data_mask = _writeQueueVec_fifo_1_empty ? writeQueueVec_1_enq_bits_data_mask : writeQueueVec_dataOut_1_data_mask;
  assign writeQueueVec_1_deq_bits_data_data = _writeQueueVec_fifo_1_empty ? writeQueueVec_1_enq_bits_data_data : writeQueueVec_dataOut_1_data_data;
  assign writeQueueVec_1_deq_bits_data_last = _writeQueueVec_fifo_1_empty ? writeQueueVec_1_enq_bits_data_last : writeQueueVec_dataOut_1_data_last;
  assign writeQueueVec_1_deq_bits_data_instructionIndex = _writeQueueVec_fifo_1_empty ? writeQueueVec_1_enq_bits_data_instructionIndex : writeQueueVec_dataOut_1_data_instructionIndex;
  wire [3:0]          writeQueueVec_1_deq_bits_targetLane = _writeQueueVec_fifo_1_empty ? 4'h2 : writeQueueVec_dataOut_1_targetLane;
  wire                vrfWritePort_2_valid_0 = writeQueueVec_2_deq_valid;
  wire [4:0]          vrfWritePort_2_bits_vd_0 = writeQueueVec_2_deq_bits_data_vd;
  wire [8:0]          vrfWritePort_2_bits_offset_0 = writeQueueVec_2_deq_bits_data_offset;
  wire [3:0]          vrfWritePort_2_bits_mask_0 = writeQueueVec_2_deq_bits_data_mask;
  wire [31:0]         vrfWritePort_2_bits_data_0 = writeQueueVec_2_deq_bits_data_data;
  wire                vrfWritePort_2_bits_last_0 = writeQueueVec_2_deq_bits_data_last;
  wire [2:0]          vrfWritePort_2_bits_instructionIndex_0 = writeQueueVec_2_deq_bits_data_instructionIndex;
  wire [2:0]          writeIndexQueue_2_enq_bits = writeQueueVec_2_deq_bits_data_instructionIndex;
  wire [31:0]         writeQueueVec_2_enq_bits_data_data;
  wire                writeQueueVec_2_enq_bits_data_last;
  wire [32:0]         writeQueueVec_dataIn_lo_hi_2 = {writeQueueVec_2_enq_bits_data_data, writeQueueVec_2_enq_bits_data_last};
  wire [2:0]          writeQueueVec_2_enq_bits_data_instructionIndex;
  wire [35:0]         writeQueueVec_dataIn_lo_2 = {writeQueueVec_dataIn_lo_hi_2, writeQueueVec_2_enq_bits_data_instructionIndex};
  wire [4:0]          writeQueueVec_2_enq_bits_data_vd;
  wire [8:0]          writeQueueVec_2_enq_bits_data_offset;
  wire [13:0]         writeQueueVec_dataIn_hi_hi_2 = {writeQueueVec_2_enq_bits_data_vd, writeQueueVec_2_enq_bits_data_offset};
  wire [3:0]          writeQueueVec_2_enq_bits_data_mask;
  wire [17:0]         writeQueueVec_dataIn_hi_2 = {writeQueueVec_dataIn_hi_hi_2, writeQueueVec_2_enq_bits_data_mask};
  wire [57:0]         writeQueueVec_dataIn_2 = {writeQueueVec_dataIn_hi_2, writeQueueVec_dataIn_lo_2, 4'h4};
  wire [3:0]          writeQueueVec_dataOut_2_targetLane = _writeQueueVec_fifo_2_data_out[3:0];
  wire [2:0]          writeQueueVec_dataOut_2_data_instructionIndex = _writeQueueVec_fifo_2_data_out[6:4];
  wire                writeQueueVec_dataOut_2_data_last = _writeQueueVec_fifo_2_data_out[7];
  wire [31:0]         writeQueueVec_dataOut_2_data_data = _writeQueueVec_fifo_2_data_out[39:8];
  wire [3:0]          writeQueueVec_dataOut_2_data_mask = _writeQueueVec_fifo_2_data_out[43:40];
  wire [8:0]          writeQueueVec_dataOut_2_data_offset = _writeQueueVec_fifo_2_data_out[52:44];
  wire [4:0]          writeQueueVec_dataOut_2_data_vd = _writeQueueVec_fifo_2_data_out[57:53];
  wire                writeQueueVec_2_enq_ready = ~_writeQueueVec_fifo_2_full;
  wire                writeQueueVec_2_enq_valid;
  wire                _probeWire_slots_2_writeValid_T = writeQueueVec_2_enq_ready & writeQueueVec_2_enq_valid;
  assign writeQueueVec_2_deq_valid = ~_writeQueueVec_fifo_2_empty | writeQueueVec_2_enq_valid;
  assign writeQueueVec_2_deq_bits_data_vd = _writeQueueVec_fifo_2_empty ? writeQueueVec_2_enq_bits_data_vd : writeQueueVec_dataOut_2_data_vd;
  assign writeQueueVec_2_deq_bits_data_offset = _writeQueueVec_fifo_2_empty ? writeQueueVec_2_enq_bits_data_offset : writeQueueVec_dataOut_2_data_offset;
  assign writeQueueVec_2_deq_bits_data_mask = _writeQueueVec_fifo_2_empty ? writeQueueVec_2_enq_bits_data_mask : writeQueueVec_dataOut_2_data_mask;
  assign writeQueueVec_2_deq_bits_data_data = _writeQueueVec_fifo_2_empty ? writeQueueVec_2_enq_bits_data_data : writeQueueVec_dataOut_2_data_data;
  assign writeQueueVec_2_deq_bits_data_last = _writeQueueVec_fifo_2_empty ? writeQueueVec_2_enq_bits_data_last : writeQueueVec_dataOut_2_data_last;
  assign writeQueueVec_2_deq_bits_data_instructionIndex = _writeQueueVec_fifo_2_empty ? writeQueueVec_2_enq_bits_data_instructionIndex : writeQueueVec_dataOut_2_data_instructionIndex;
  wire [3:0]          writeQueueVec_2_deq_bits_targetLane = _writeQueueVec_fifo_2_empty ? 4'h4 : writeQueueVec_dataOut_2_targetLane;
  wire                vrfWritePort_3_valid_0 = writeQueueVec_3_deq_valid;
  wire [4:0]          vrfWritePort_3_bits_vd_0 = writeQueueVec_3_deq_bits_data_vd;
  wire [8:0]          vrfWritePort_3_bits_offset_0 = writeQueueVec_3_deq_bits_data_offset;
  wire [3:0]          vrfWritePort_3_bits_mask_0 = writeQueueVec_3_deq_bits_data_mask;
  wire [31:0]         vrfWritePort_3_bits_data_0 = writeQueueVec_3_deq_bits_data_data;
  wire                vrfWritePort_3_bits_last_0 = writeQueueVec_3_deq_bits_data_last;
  wire [2:0]          vrfWritePort_3_bits_instructionIndex_0 = writeQueueVec_3_deq_bits_data_instructionIndex;
  wire [2:0]          writeIndexQueue_3_enq_bits = writeQueueVec_3_deq_bits_data_instructionIndex;
  wire [31:0]         writeQueueVec_3_enq_bits_data_data;
  wire                writeQueueVec_3_enq_bits_data_last;
  wire [32:0]         writeQueueVec_dataIn_lo_hi_3 = {writeQueueVec_3_enq_bits_data_data, writeQueueVec_3_enq_bits_data_last};
  wire [2:0]          writeQueueVec_3_enq_bits_data_instructionIndex;
  wire [35:0]         writeQueueVec_dataIn_lo_3 = {writeQueueVec_dataIn_lo_hi_3, writeQueueVec_3_enq_bits_data_instructionIndex};
  wire [4:0]          writeQueueVec_3_enq_bits_data_vd;
  wire [8:0]          writeQueueVec_3_enq_bits_data_offset;
  wire [13:0]         writeQueueVec_dataIn_hi_hi_3 = {writeQueueVec_3_enq_bits_data_vd, writeQueueVec_3_enq_bits_data_offset};
  wire [3:0]          writeQueueVec_3_enq_bits_data_mask;
  wire [17:0]         writeQueueVec_dataIn_hi_3 = {writeQueueVec_dataIn_hi_hi_3, writeQueueVec_3_enq_bits_data_mask};
  wire [57:0]         writeQueueVec_dataIn_3 = {writeQueueVec_dataIn_hi_3, writeQueueVec_dataIn_lo_3, 4'h8};
  wire [3:0]          writeQueueVec_dataOut_3_targetLane = _writeQueueVec_fifo_3_data_out[3:0];
  wire [2:0]          writeQueueVec_dataOut_3_data_instructionIndex = _writeQueueVec_fifo_3_data_out[6:4];
  wire                writeQueueVec_dataOut_3_data_last = _writeQueueVec_fifo_3_data_out[7];
  wire [31:0]         writeQueueVec_dataOut_3_data_data = _writeQueueVec_fifo_3_data_out[39:8];
  wire [3:0]          writeQueueVec_dataOut_3_data_mask = _writeQueueVec_fifo_3_data_out[43:40];
  wire [8:0]          writeQueueVec_dataOut_3_data_offset = _writeQueueVec_fifo_3_data_out[52:44];
  wire [4:0]          writeQueueVec_dataOut_3_data_vd = _writeQueueVec_fifo_3_data_out[57:53];
  wire                writeQueueVec_3_enq_ready = ~_writeQueueVec_fifo_3_full;
  wire                writeQueueVec_3_enq_valid;
  wire                _probeWire_slots_3_writeValid_T = writeQueueVec_3_enq_ready & writeQueueVec_3_enq_valid;
  assign writeQueueVec_3_deq_valid = ~_writeQueueVec_fifo_3_empty | writeQueueVec_3_enq_valid;
  assign writeQueueVec_3_deq_bits_data_vd = _writeQueueVec_fifo_3_empty ? writeQueueVec_3_enq_bits_data_vd : writeQueueVec_dataOut_3_data_vd;
  assign writeQueueVec_3_deq_bits_data_offset = _writeQueueVec_fifo_3_empty ? writeQueueVec_3_enq_bits_data_offset : writeQueueVec_dataOut_3_data_offset;
  assign writeQueueVec_3_deq_bits_data_mask = _writeQueueVec_fifo_3_empty ? writeQueueVec_3_enq_bits_data_mask : writeQueueVec_dataOut_3_data_mask;
  assign writeQueueVec_3_deq_bits_data_data = _writeQueueVec_fifo_3_empty ? writeQueueVec_3_enq_bits_data_data : writeQueueVec_dataOut_3_data_data;
  assign writeQueueVec_3_deq_bits_data_last = _writeQueueVec_fifo_3_empty ? writeQueueVec_3_enq_bits_data_last : writeQueueVec_dataOut_3_data_last;
  assign writeQueueVec_3_deq_bits_data_instructionIndex = _writeQueueVec_fifo_3_empty ? writeQueueVec_3_enq_bits_data_instructionIndex : writeQueueVec_dataOut_3_data_instructionIndex;
  wire [3:0]          writeQueueVec_3_deq_bits_targetLane = _writeQueueVec_fifo_3_empty ? 4'h8 : writeQueueVec_dataOut_3_targetLane;
  wire                otherUnitTargetQueue_deq_valid;
  assign otherUnitTargetQueue_deq_valid = ~_otherUnitTargetQueue_fifo_empty;
  wire                otherUnitTargetQueue_deq_ready;
  wire                otherUnitTargetQueue_enq_ready = ~_otherUnitTargetQueue_fifo_full | otherUnitTargetQueue_deq_ready;
  wire                otherUnitTargetQueue_enq_valid;
  wire                otherUnitDataQueueVec_0_enq_ready = ~_otherUnitDataQueueVec_fifo_full;
  wire                otherUnitDataQueueVec_0_deq_ready;
  wire                otherUnitDataQueueVec_0_enq_valid;
  wire                otherUnitDataQueueVec_0_deq_valid = ~_otherUnitDataQueueVec_fifo_empty | otherUnitDataQueueVec_0_enq_valid;
  wire [31:0]         otherUnitDataQueueVec_0_deq_bits = _otherUnitDataQueueVec_fifo_empty ? otherUnitDataQueueVec_0_enq_bits : _otherUnitDataQueueVec_fifo_data_out;
  wire                otherUnitDataQueueVec_1_enq_ready = ~_otherUnitDataQueueVec_fifo_1_full;
  wire                otherUnitDataQueueVec_1_deq_ready;
  wire                otherUnitDataQueueVec_1_enq_valid;
  wire                otherUnitDataQueueVec_1_deq_valid = ~_otherUnitDataQueueVec_fifo_1_empty | otherUnitDataQueueVec_1_enq_valid;
  wire [31:0]         otherUnitDataQueueVec_1_deq_bits = _otherUnitDataQueueVec_fifo_1_empty ? otherUnitDataQueueVec_1_enq_bits : _otherUnitDataQueueVec_fifo_1_data_out;
  wire                otherUnitDataQueueVec_2_enq_ready = ~_otherUnitDataQueueVec_fifo_2_full;
  wire                otherUnitDataQueueVec_2_deq_ready;
  wire                otherUnitDataQueueVec_2_enq_valid;
  wire                otherUnitDataQueueVec_2_deq_valid = ~_otherUnitDataQueueVec_fifo_2_empty | otherUnitDataQueueVec_2_enq_valid;
  wire [31:0]         otherUnitDataQueueVec_2_deq_bits = _otherUnitDataQueueVec_fifo_2_empty ? otherUnitDataQueueVec_2_enq_bits : _otherUnitDataQueueVec_fifo_2_data_out;
  wire                otherUnitDataQueueVec_3_enq_ready = ~_otherUnitDataQueueVec_fifo_3_full;
  wire                otherUnitDataQueueVec_3_deq_ready;
  wire                otherUnitDataQueueVec_3_enq_valid;
  wire                otherUnitDataQueueVec_3_deq_valid = ~_otherUnitDataQueueVec_fifo_3_empty | otherUnitDataQueueVec_3_enq_valid;
  wire [31:0]         otherUnitDataQueueVec_3_deq_bits = _otherUnitDataQueueVec_fifo_3_empty ? otherUnitDataQueueVec_3_enq_bits : _otherUnitDataQueueVec_fifo_3_data_out;
  wire [3:0]          otherTryReadVrf = _otherUnit_vrfReadDataPorts_valid ? _otherUnit_status_targetLane : 4'h0;
  wire                vrfReadDataPorts_0_valid_0 = otherTryReadVrf[0] | _storeUnit_vrfReadDataPorts_0_valid;
  wire [4:0]          vrfReadDataPorts_0_bits_vs_0 = otherTryReadVrf[0] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_0_bits_vs;
  wire [8:0]          vrfReadDataPorts_0_bits_offset_0 = otherTryReadVrf[0] ? _otherUnit_vrfReadDataPorts_bits_offset : _storeUnit_vrfReadDataPorts_0_bits_offset;
  wire [2:0]          vrfReadDataPorts_0_bits_instructionIndex_0 = otherTryReadVrf[0] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_0_bits_instructionIndex;
  wire                otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_0_enq_valid = vrfReadResults_0_valid & ~otherUnitTargetQueue_empty;
  wire [3:0]          dataDeqFire;
  assign otherUnitDataQueueVec_0_deq_ready = dataDeqFire[0];
  wire                vrfReadDataPorts_1_valid_0 = otherTryReadVrf[1] | _storeUnit_vrfReadDataPorts_1_valid;
  wire [4:0]          vrfReadDataPorts_1_bits_vs_0 = otherTryReadVrf[1] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_1_bits_vs;
  wire [8:0]          vrfReadDataPorts_1_bits_offset_0 = otherTryReadVrf[1] ? _otherUnit_vrfReadDataPorts_bits_offset : _storeUnit_vrfReadDataPorts_1_bits_offset;
  wire [2:0]          vrfReadDataPorts_1_bits_instructionIndex_0 = otherTryReadVrf[1] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_1_bits_instructionIndex;
  assign otherUnitDataQueueVec_1_enq_valid = vrfReadResults_1_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_1_deq_ready = dataDeqFire[1];
  wire                vrfReadDataPorts_2_valid_0 = otherTryReadVrf[2] | _storeUnit_vrfReadDataPorts_2_valid;
  wire [4:0]          vrfReadDataPorts_2_bits_vs_0 = otherTryReadVrf[2] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_2_bits_vs;
  wire [8:0]          vrfReadDataPorts_2_bits_offset_0 = otherTryReadVrf[2] ? _otherUnit_vrfReadDataPorts_bits_offset : _storeUnit_vrfReadDataPorts_2_bits_offset;
  wire [2:0]          vrfReadDataPorts_2_bits_instructionIndex_0 = otherTryReadVrf[2] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_2_bits_instructionIndex;
  assign otherUnitDataQueueVec_2_enq_valid = vrfReadResults_2_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_2_deq_ready = dataDeqFire[2];
  wire                vrfReadDataPorts_3_valid_0 = otherTryReadVrf[3] | _storeUnit_vrfReadDataPorts_3_valid;
  wire [4:0]          vrfReadDataPorts_3_bits_vs_0 = otherTryReadVrf[3] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_3_bits_vs;
  wire [8:0]          vrfReadDataPorts_3_bits_offset_0 = otherTryReadVrf[3] ? _otherUnit_vrfReadDataPorts_bits_offset : _storeUnit_vrfReadDataPorts_3_bits_offset;
  wire [2:0]          vrfReadDataPorts_3_bits_instructionIndex_0 = otherTryReadVrf[3] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_3_bits_instructionIndex;
  assign otherUnitDataQueueVec_3_enq_valid = vrfReadResults_3_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_3_deq_ready = dataDeqFire[3];
  wire [1:0]          otherUnit_vrfReadDataPorts_ready_lo = {vrfReadDataPorts_1_ready_0, vrfReadDataPorts_0_ready_0};
  wire [1:0]          otherUnit_vrfReadDataPorts_ready_hi = {vrfReadDataPorts_3_ready_0, vrfReadDataPorts_2_ready_0};
  wire                otherUnit_vrfReadDataPorts_ready = (|(otherTryReadVrf & {otherUnit_vrfReadDataPorts_ready_hi, otherUnit_vrfReadDataPorts_ready_lo})) & otherUnitTargetQueue_enq_ready;
  assign otherUnitTargetQueue_enq_valid = otherUnit_vrfReadDataPorts_ready & _otherUnit_vrfReadDataPorts_valid;
  wire [3:0]          otherUnitTargetQueue_deq_bits;
  wire [1:0]          otherUnit_vrfReadResults_valid_lo = {otherUnitDataQueueVec_1_deq_valid, otherUnitDataQueueVec_0_deq_valid};
  wire [1:0]          otherUnit_vrfReadResults_valid_hi = {otherUnitDataQueueVec_3_deq_valid, otherUnitDataQueueVec_2_deq_valid};
  assign otherUnitTargetQueue_deq_ready = otherUnitTargetQueue_deq_valid & (|(otherUnitTargetQueue_deq_bits & {otherUnit_vrfReadResults_valid_hi, otherUnit_vrfReadResults_valid_lo}));
  assign dataDeqFire = otherUnitTargetQueue_deq_ready ? otherUnitTargetQueue_deq_bits : 4'h0;
  wire [3:0]          otherTryToWrite = _otherUnit_vrfWritePort_valid ? _otherUnit_status_targetLane : 4'h0;
  wire [1:0]          otherUnit_vrfWritePort_ready_lo = {writeQueueVec_1_enq_ready, writeQueueVec_0_enq_ready};
  wire [1:0]          otherUnit_vrfWritePort_ready_hi = {writeQueueVec_3_enq_ready, writeQueueVec_2_enq_ready};
  assign writeQueueVec_0_enq_valid = otherTryToWrite[0] | _loadUnit_vrfWritePort_0_valid;
  assign writeQueueVec_0_enq_bits_data_vd = otherTryToWrite[0] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_0_bits_vd;
  assign writeQueueVec_0_enq_bits_data_offset = otherTryToWrite[0] ? _otherUnit_vrfWritePort_bits_offset : _loadUnit_vrfWritePort_0_bits_offset;
  assign writeQueueVec_0_enq_bits_data_mask = otherTryToWrite[0] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_0_bits_mask;
  assign writeQueueVec_0_enq_bits_data_data = otherTryToWrite[0] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_0_bits_data;
  assign writeQueueVec_0_enq_bits_data_last = otherTryToWrite[0] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_0_enq_bits_data_instructionIndex = otherTryToWrite[0] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_0_bits_instructionIndex;
  assign writeQueueVec_1_enq_valid = otherTryToWrite[1] | _loadUnit_vrfWritePort_1_valid;
  assign writeQueueVec_1_enq_bits_data_vd = otherTryToWrite[1] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_1_bits_vd;
  assign writeQueueVec_1_enq_bits_data_offset = otherTryToWrite[1] ? _otherUnit_vrfWritePort_bits_offset : _loadUnit_vrfWritePort_1_bits_offset;
  assign writeQueueVec_1_enq_bits_data_mask = otherTryToWrite[1] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_1_bits_mask;
  assign writeQueueVec_1_enq_bits_data_data = otherTryToWrite[1] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_1_bits_data;
  assign writeQueueVec_1_enq_bits_data_last = otherTryToWrite[1] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_1_enq_bits_data_instructionIndex = otherTryToWrite[1] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_1_bits_instructionIndex;
  assign writeQueueVec_2_enq_valid = otherTryToWrite[2] | _loadUnit_vrfWritePort_2_valid;
  assign writeQueueVec_2_enq_bits_data_vd = otherTryToWrite[2] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_2_bits_vd;
  assign writeQueueVec_2_enq_bits_data_offset = otherTryToWrite[2] ? _otherUnit_vrfWritePort_bits_offset : _loadUnit_vrfWritePort_2_bits_offset;
  assign writeQueueVec_2_enq_bits_data_mask = otherTryToWrite[2] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_2_bits_mask;
  assign writeQueueVec_2_enq_bits_data_data = otherTryToWrite[2] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_2_bits_data;
  assign writeQueueVec_2_enq_bits_data_last = otherTryToWrite[2] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_2_enq_bits_data_instructionIndex = otherTryToWrite[2] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_2_bits_instructionIndex;
  assign writeQueueVec_3_enq_valid = otherTryToWrite[3] | _loadUnit_vrfWritePort_3_valid;
  assign writeQueueVec_3_enq_bits_data_vd = otherTryToWrite[3] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_3_bits_vd;
  assign writeQueueVec_3_enq_bits_data_offset = otherTryToWrite[3] ? _otherUnit_vrfWritePort_bits_offset : _loadUnit_vrfWritePort_3_bits_offset;
  assign writeQueueVec_3_enq_bits_data_mask = otherTryToWrite[3] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_3_bits_mask;
  assign writeQueueVec_3_enq_bits_data_data = otherTryToWrite[3] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_3_bits_data;
  assign writeQueueVec_3_enq_bits_data_last = otherTryToWrite[3] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_3_enq_bits_data_instructionIndex = otherTryToWrite[3] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_3_bits_instructionIndex;
  wire [7:0]          _GEN_1026 = {5'h0, _loadUnit_status_instructionIndex};
  wire [7:0]          _GEN_1027 = {5'h0, _otherUnit_status_instructionIndex};
  wire [7:0]          dataInMSHR = (_loadUnit_status_idle ? 8'h0 : 8'h1 << _GEN_1026) | (_otherUnit_status_idle | _otherUnit_status_isStore ? 8'h0 : 8'h1 << _GEN_1027);
  reg  [6:0]          queueCount_0;
  reg  [6:0]          queueCount_1;
  reg  [6:0]          queueCount_2;
  reg  [6:0]          queueCount_3;
  reg  [6:0]          queueCount_4;
  reg  [6:0]          queueCount_5;
  reg  [6:0]          queueCount_6;
  reg  [6:0]          queueCount_7;
  wire [7:0]          enqOH = 8'h1 << writeQueueVec_0_enq_bits_data_instructionIndex;
  wire [7:0]          queueEnq = _probeWire_slots_0_writeValid_T ? enqOH : 8'h0;
  wire                writeIndexQueue_deq_valid;
  assign writeIndexQueue_deq_valid = ~_writeIndexQueue_fifo_empty;
  wire                writeIndexQueue_enq_ready = ~_writeIndexQueue_fifo_full;
  wire                writeIndexQueue_enq_valid;
  assign writeIndexQueue_enq_valid = writeQueueVec_0_deq_ready & writeQueueVec_0_deq_valid;
  wire [2:0]          writeIndexQueue_deq_bits;
  wire [7:0]          queueDeq = writeIndexQueue_deq_ready & writeIndexQueue_deq_valid ? 8'h1 << writeIndexQueue_deq_bits : 8'h0;
  wire [6:0]          counterUpdate = queueEnq[0] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_1 = queueEnq[1] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_2 = queueEnq[2] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_3 = queueEnq[3] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_4 = queueEnq[4] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_5 = queueEnq[5] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_6 = queueEnq[6] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_7 = queueEnq[7] ? 7'h1 : 7'h7F;
  wire [1:0]          dataInWriteQueue_0_lo_lo = {|queueCount_1, |queueCount_0};
  wire [1:0]          dataInWriteQueue_0_lo_hi = {|queueCount_3, |queueCount_2};
  wire [3:0]          dataInWriteQueue_0_lo = {dataInWriteQueue_0_lo_hi, dataInWriteQueue_0_lo_lo};
  wire [1:0]          dataInWriteQueue_0_hi_lo = {|queueCount_5, |queueCount_4};
  wire [1:0]          dataInWriteQueue_0_hi_hi = {|queueCount_7, |queueCount_6};
  wire [3:0]          dataInWriteQueue_0_hi = {dataInWriteQueue_0_hi_hi, dataInWriteQueue_0_hi_lo};
  reg  [6:0]          queueCount_0_1;
  reg  [6:0]          queueCount_1_1;
  reg  [6:0]          queueCount_2_1;
  reg  [6:0]          queueCount_3_1;
  reg  [6:0]          queueCount_4_1;
  reg  [6:0]          queueCount_5_1;
  reg  [6:0]          queueCount_6_1;
  reg  [6:0]          queueCount_7_1;
  wire [7:0]          enqOH_1 = 8'h1 << writeQueueVec_1_enq_bits_data_instructionIndex;
  wire [7:0]          queueEnq_1 = _probeWire_slots_1_writeValid_T ? enqOH_1 : 8'h0;
  wire                writeIndexQueue_1_deq_valid;
  assign writeIndexQueue_1_deq_valid = ~_writeIndexQueue_fifo_1_empty;
  wire                writeIndexQueue_1_enq_ready = ~_writeIndexQueue_fifo_1_full;
  wire                writeIndexQueue_1_enq_valid;
  assign writeIndexQueue_1_enq_valid = writeQueueVec_1_deq_ready & writeQueueVec_1_deq_valid;
  wire [2:0]          writeIndexQueue_1_deq_bits;
  wire [7:0]          queueDeq_1 = writeIndexQueue_1_deq_ready & writeIndexQueue_1_deq_valid ? 8'h1 << writeIndexQueue_1_deq_bits : 8'h0;
  wire [6:0]          counterUpdate_8 = queueEnq_1[0] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_9 = queueEnq_1[1] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_10 = queueEnq_1[2] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_11 = queueEnq_1[3] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_12 = queueEnq_1[4] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_13 = queueEnq_1[5] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_14 = queueEnq_1[6] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_15 = queueEnq_1[7] ? 7'h1 : 7'h7F;
  wire [1:0]          dataInWriteQueue_1_lo_lo = {|queueCount_1_1, |queueCount_0_1};
  wire [1:0]          dataInWriteQueue_1_lo_hi = {|queueCount_3_1, |queueCount_2_1};
  wire [3:0]          dataInWriteQueue_1_lo = {dataInWriteQueue_1_lo_hi, dataInWriteQueue_1_lo_lo};
  wire [1:0]          dataInWriteQueue_1_hi_lo = {|queueCount_5_1, |queueCount_4_1};
  wire [1:0]          dataInWriteQueue_1_hi_hi = {|queueCount_7_1, |queueCount_6_1};
  wire [3:0]          dataInWriteQueue_1_hi = {dataInWriteQueue_1_hi_hi, dataInWriteQueue_1_hi_lo};
  reg  [6:0]          queueCount_0_2;
  reg  [6:0]          queueCount_1_2;
  reg  [6:0]          queueCount_2_2;
  reg  [6:0]          queueCount_3_2;
  reg  [6:0]          queueCount_4_2;
  reg  [6:0]          queueCount_5_2;
  reg  [6:0]          queueCount_6_2;
  reg  [6:0]          queueCount_7_2;
  wire [7:0]          enqOH_2 = 8'h1 << writeQueueVec_2_enq_bits_data_instructionIndex;
  wire [7:0]          queueEnq_2 = _probeWire_slots_2_writeValid_T ? enqOH_2 : 8'h0;
  wire                writeIndexQueue_2_deq_valid;
  assign writeIndexQueue_2_deq_valid = ~_writeIndexQueue_fifo_2_empty;
  wire                writeIndexQueue_2_enq_ready = ~_writeIndexQueue_fifo_2_full;
  wire                writeIndexQueue_2_enq_valid;
  assign writeIndexQueue_2_enq_valid = writeQueueVec_2_deq_ready & writeQueueVec_2_deq_valid;
  wire [2:0]          writeIndexQueue_2_deq_bits;
  wire [7:0]          queueDeq_2 = writeIndexQueue_2_deq_ready & writeIndexQueue_2_deq_valid ? 8'h1 << writeIndexQueue_2_deq_bits : 8'h0;
  wire [6:0]          counterUpdate_16 = queueEnq_2[0] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_17 = queueEnq_2[1] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_18 = queueEnq_2[2] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_19 = queueEnq_2[3] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_20 = queueEnq_2[4] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_21 = queueEnq_2[5] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_22 = queueEnq_2[6] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_23 = queueEnq_2[7] ? 7'h1 : 7'h7F;
  wire [1:0]          dataInWriteQueue_2_lo_lo = {|queueCount_1_2, |queueCount_0_2};
  wire [1:0]          dataInWriteQueue_2_lo_hi = {|queueCount_3_2, |queueCount_2_2};
  wire [3:0]          dataInWriteQueue_2_lo = {dataInWriteQueue_2_lo_hi, dataInWriteQueue_2_lo_lo};
  wire [1:0]          dataInWriteQueue_2_hi_lo = {|queueCount_5_2, |queueCount_4_2};
  wire [1:0]          dataInWriteQueue_2_hi_hi = {|queueCount_7_2, |queueCount_6_2};
  wire [3:0]          dataInWriteQueue_2_hi = {dataInWriteQueue_2_hi_hi, dataInWriteQueue_2_hi_lo};
  reg  [6:0]          queueCount_0_3;
  reg  [6:0]          queueCount_1_3;
  reg  [6:0]          queueCount_2_3;
  reg  [6:0]          queueCount_3_3;
  reg  [6:0]          queueCount_4_3;
  reg  [6:0]          queueCount_5_3;
  reg  [6:0]          queueCount_6_3;
  reg  [6:0]          queueCount_7_3;
  wire [7:0]          enqOH_3 = 8'h1 << writeQueueVec_3_enq_bits_data_instructionIndex;
  wire [7:0]          queueEnq_3 = _probeWire_slots_3_writeValid_T ? enqOH_3 : 8'h0;
  wire                writeIndexQueue_3_deq_valid;
  assign writeIndexQueue_3_deq_valid = ~_writeIndexQueue_fifo_3_empty;
  wire                writeIndexQueue_3_enq_ready = ~_writeIndexQueue_fifo_3_full;
  wire                writeIndexQueue_3_enq_valid;
  assign writeIndexQueue_3_enq_valid = writeQueueVec_3_deq_ready & writeQueueVec_3_deq_valid;
  wire [2:0]          writeIndexQueue_3_deq_bits;
  wire [7:0]          queueDeq_3 = writeIndexQueue_3_deq_ready & writeIndexQueue_3_deq_valid ? 8'h1 << writeIndexQueue_3_deq_bits : 8'h0;
  wire [6:0]          counterUpdate_24 = queueEnq_3[0] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_25 = queueEnq_3[1] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_26 = queueEnq_3[2] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_27 = queueEnq_3[3] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_28 = queueEnq_3[4] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_29 = queueEnq_3[5] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_30 = queueEnq_3[6] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_31 = queueEnq_3[7] ? 7'h1 : 7'h7F;
  wire [1:0]          dataInWriteQueue_3_lo_lo = {|queueCount_1_3, |queueCount_0_3};
  wire [1:0]          dataInWriteQueue_3_lo_hi = {|queueCount_3_3, |queueCount_2_3};
  wire [3:0]          dataInWriteQueue_3_lo = {dataInWriteQueue_3_lo_hi, dataInWriteQueue_3_lo_lo};
  wire [1:0]          dataInWriteQueue_3_hi_lo = {|queueCount_5_3, |queueCount_4_3};
  wire [1:0]          dataInWriteQueue_3_hi_hi = {|queueCount_7_3, |queueCount_6_3};
  wire [3:0]          dataInWriteQueue_3_hi = {dataInWriteQueue_3_hi_hi, dataInWriteQueue_3_hi_lo};
  wire                sourceQueue_deq_valid;
  assign sourceQueue_deq_valid = ~_sourceQueue_fifo_empty;
  wire                sourceQueue_enq_ready = ~_sourceQueue_fifo_full;
  wire                sourceQueue_enq_valid;
  wire                sourceQueue_deq_ready;
  wire                axi4Port_ar_valid_0 = _loadUnit_memRequest_valid & sourceQueue_enq_ready;
  wire                axi4Port_r_ready_0;
  assign sourceQueue_enq_valid = _loadUnit_memRequest_valid & axi4Port_ar_ready_0;
  assign sourceQueue_deq_ready = axi4Port_r_ready_0 & axi4Port_r_valid_0;
  assign dataQueue_deq_valid = ~_dataQueue_fifo_empty;
  wire                axi4Port_w_valid_0 = dataQueue_deq_valid;
  wire [127:0]        dataQueue_dataOut_data;
  wire [127:0]        axi4Port_w_bits_data_0 = dataQueue_deq_bits_data;
  wire [15:0]         dataQueue_dataOut_mask;
  wire [15:0]         axi4Port_w_bits_strb_0 = dataQueue_deq_bits_mask;
  wire [12:0]         dataQueue_dataOut_index;
  wire [31:0]         dataQueue_dataOut_address;
  wire [12:0]         dataQueue_enq_bits_index;
  wire [31:0]         dataQueue_enq_bits_address;
  wire [44:0]         dataQueue_dataIn_lo = {dataQueue_enq_bits_index, dataQueue_enq_bits_address};
  wire [127:0]        dataQueue_enq_bits_data;
  wire [15:0]         dataQueue_enq_bits_mask;
  wire [143:0]        dataQueue_dataIn_hi = {dataQueue_enq_bits_data, dataQueue_enq_bits_mask};
  wire [188:0]        dataQueue_dataIn = {dataQueue_dataIn_hi, dataQueue_dataIn_lo};
  assign dataQueue_dataOut_address = _dataQueue_fifo_data_out[31:0];
  assign dataQueue_dataOut_index = _dataQueue_fifo_data_out[44:32];
  assign dataQueue_dataOut_mask = _dataQueue_fifo_data_out[60:45];
  assign dataQueue_dataOut_data = _dataQueue_fifo_data_out[188:61];
  assign dataQueue_deq_bits_data = dataQueue_dataOut_data;
  assign dataQueue_deq_bits_mask = dataQueue_dataOut_mask;
  wire [12:0]         dataQueue_deq_bits_index = dataQueue_dataOut_index;
  wire [31:0]         dataQueue_deq_bits_address = dataQueue_dataOut_address;
  wire                dataQueue_enq_ready = ~_dataQueue_fifo_full;
  wire                dataQueue_enq_valid;
  wire                axi4Port_aw_valid_0 = _storeUnit_memRequest_valid & dataQueue_enq_ready;
  wire [1:0]          axi4Port_aw_bits_id_0 = _storeUnit_memRequest_bits_index[1:0];
  assign dataQueue_enq_valid = _storeUnit_memRequest_valid & axi4Port_aw_ready_0;
  wire                simpleSourceQueue_deq_valid;
  assign simpleSourceQueue_deq_valid = ~_simpleSourceQueue_fifo_empty;
  wire                simpleSourceQueue_enq_ready = ~_simpleSourceQueue_fifo_full;
  wire                simpleSourceQueue_enq_valid;
  wire                simpleSourceQueue_deq_ready;
  wire                simpleAccessPorts_ar_valid_0 = _otherUnit_memReadRequest_valid & simpleSourceQueue_enq_ready;
  wire                simpleAccessPorts_r_ready_0;
  assign simpleSourceQueue_enq_valid = _otherUnit_memReadRequest_valid & simpleAccessPorts_ar_ready_0;
  assign simpleSourceQueue_deq_ready = simpleAccessPorts_r_ready_0 & simpleAccessPorts_r_valid_0;
  assign simpleDataQueue_deq_valid = ~_simpleDataQueue_fifo_empty;
  wire                simpleAccessPorts_w_valid_0 = simpleDataQueue_deq_valid;
  wire [31:0]         simpleDataQueue_dataOut_data;
  wire [31:0]         simpleAccessPorts_w_bits_data_0 = simpleDataQueue_deq_bits_data;
  wire [3:0]          simpleDataQueue_dataOut_mask;
  wire [3:0]          simpleAccessPorts_w_bits_strb_0 = simpleDataQueue_deq_bits_mask;
  wire [7:0]          simpleDataQueue_dataOut_source;
  wire [31:0]         simpleDataQueue_dataOut_address;
  wire [1:0]          simpleDataQueue_dataOut_size;
  wire [31:0]         simpleDataQueue_enq_bits_address;
  wire [1:0]          simpleDataQueue_enq_bits_size;
  wire [33:0]         simpleDataQueue_dataIn_lo = {simpleDataQueue_enq_bits_address, simpleDataQueue_enq_bits_size};
  wire [31:0]         simpleDataQueue_enq_bits_data;
  wire [3:0]          simpleDataQueue_enq_bits_mask;
  wire [35:0]         simpleDataQueue_dataIn_hi_hi = {simpleDataQueue_enq_bits_data, simpleDataQueue_enq_bits_mask};
  wire [7:0]          simpleDataQueue_enq_bits_source;
  wire [43:0]         simpleDataQueue_dataIn_hi = {simpleDataQueue_dataIn_hi_hi, simpleDataQueue_enq_bits_source};
  wire [77:0]         simpleDataQueue_dataIn = {simpleDataQueue_dataIn_hi, simpleDataQueue_dataIn_lo};
  assign simpleDataQueue_dataOut_size = _simpleDataQueue_fifo_data_out[1:0];
  assign simpleDataQueue_dataOut_address = _simpleDataQueue_fifo_data_out[33:2];
  assign simpleDataQueue_dataOut_source = _simpleDataQueue_fifo_data_out[41:34];
  assign simpleDataQueue_dataOut_mask = _simpleDataQueue_fifo_data_out[45:42];
  assign simpleDataQueue_dataOut_data = _simpleDataQueue_fifo_data_out[77:46];
  assign simpleDataQueue_deq_bits_data = simpleDataQueue_dataOut_data;
  assign simpleDataQueue_deq_bits_mask = simpleDataQueue_dataOut_mask;
  wire [7:0]          simpleDataQueue_deq_bits_source = simpleDataQueue_dataOut_source;
  wire [31:0]         simpleDataQueue_deq_bits_address = simpleDataQueue_dataOut_address;
  wire [1:0]          simpleDataQueue_deq_bits_size = simpleDataQueue_dataOut_size;
  wire                simpleDataQueue_enq_ready = ~_simpleDataQueue_fifo_full;
  wire                simpleDataQueue_enq_valid;
  wire                simpleAccessPorts_aw_valid_0 = _otherUnit_memWriteRequest_valid & dataQueue_enq_ready;
  wire [2:0]          simpleAccessPorts_aw_bits_size_0 = {1'h0, _otherUnit_memWriteRequest_bits_size};
  wire [1:0]          simpleAccessPorts_aw_bits_id_0 = _otherUnit_memWriteRequest_bits_source[1:0];
  assign simpleDataQueue_enq_valid = _otherUnit_memWriteRequest_valid & simpleAccessPorts_aw_ready_0;
  wire [1:0]          tokenIO_offsetGroupRelease_lo = {_otherUnit_offsetRelease_1, _otherUnit_offsetRelease_0};
  wire [1:0]          tokenIO_offsetGroupRelease_hi = {_otherUnit_offsetRelease_3, _otherUnit_offsetRelease_2};
  wire                unitOrder =
    _loadUnit_status_instructionIndex == _storeUnit_status_instructionIndex | _loadUnit_status_instructionIndex[1:0] < _storeUnit_status_instructionIndex[1:0] ^ _loadUnit_status_instructionIndex[2] ^ _storeUnit_status_instructionIndex[2];
  wire                loadAddressConflict = _loadUnit_status_startAddress >= _storeUnit_status_startAddress & _loadUnit_status_startAddress <= _storeUnit_status_endAddress;
  wire                storeAddressConflict = _storeUnit_status_startAddress >= _loadUnit_status_startAddress & _storeUnit_status_startAddress <= _loadUnit_status_endAddress;
  wire                stallLoad = ~unitOrder & loadAddressConflict & ~_storeUnit_status_idle;
  wire                stallStore = unitOrder & storeAddressConflict & ~_loadUnit_status_idle;
  always @(posedge clock) begin
    if (reset) begin
      v0_0 <= 32'h0;
      v0_1 <= 32'h0;
      v0_2 <= 32'h0;
      v0_3 <= 32'h0;
      v0_4 <= 32'h0;
      v0_5 <= 32'h0;
      v0_6 <= 32'h0;
      v0_7 <= 32'h0;
      v0_8 <= 32'h0;
      v0_9 <= 32'h0;
      v0_10 <= 32'h0;
      v0_11 <= 32'h0;
      v0_12 <= 32'h0;
      v0_13 <= 32'h0;
      v0_14 <= 32'h0;
      v0_15 <= 32'h0;
      v0_16 <= 32'h0;
      v0_17 <= 32'h0;
      v0_18 <= 32'h0;
      v0_19 <= 32'h0;
      v0_20 <= 32'h0;
      v0_21 <= 32'h0;
      v0_22 <= 32'h0;
      v0_23 <= 32'h0;
      v0_24 <= 32'h0;
      v0_25 <= 32'h0;
      v0_26 <= 32'h0;
      v0_27 <= 32'h0;
      v0_28 <= 32'h0;
      v0_29 <= 32'h0;
      v0_30 <= 32'h0;
      v0_31 <= 32'h0;
      v0_32 <= 32'h0;
      v0_33 <= 32'h0;
      v0_34 <= 32'h0;
      v0_35 <= 32'h0;
      v0_36 <= 32'h0;
      v0_37 <= 32'h0;
      v0_38 <= 32'h0;
      v0_39 <= 32'h0;
      v0_40 <= 32'h0;
      v0_41 <= 32'h0;
      v0_42 <= 32'h0;
      v0_43 <= 32'h0;
      v0_44 <= 32'h0;
      v0_45 <= 32'h0;
      v0_46 <= 32'h0;
      v0_47 <= 32'h0;
      v0_48 <= 32'h0;
      v0_49 <= 32'h0;
      v0_50 <= 32'h0;
      v0_51 <= 32'h0;
      v0_52 <= 32'h0;
      v0_53 <= 32'h0;
      v0_54 <= 32'h0;
      v0_55 <= 32'h0;
      v0_56 <= 32'h0;
      v0_57 <= 32'h0;
      v0_58 <= 32'h0;
      v0_59 <= 32'h0;
      v0_60 <= 32'h0;
      v0_61 <= 32'h0;
      v0_62 <= 32'h0;
      v0_63 <= 32'h0;
      v0_64 <= 32'h0;
      v0_65 <= 32'h0;
      v0_66 <= 32'h0;
      v0_67 <= 32'h0;
      v0_68 <= 32'h0;
      v0_69 <= 32'h0;
      v0_70 <= 32'h0;
      v0_71 <= 32'h0;
      v0_72 <= 32'h0;
      v0_73 <= 32'h0;
      v0_74 <= 32'h0;
      v0_75 <= 32'h0;
      v0_76 <= 32'h0;
      v0_77 <= 32'h0;
      v0_78 <= 32'h0;
      v0_79 <= 32'h0;
      v0_80 <= 32'h0;
      v0_81 <= 32'h0;
      v0_82 <= 32'h0;
      v0_83 <= 32'h0;
      v0_84 <= 32'h0;
      v0_85 <= 32'h0;
      v0_86 <= 32'h0;
      v0_87 <= 32'h0;
      v0_88 <= 32'h0;
      v0_89 <= 32'h0;
      v0_90 <= 32'h0;
      v0_91 <= 32'h0;
      v0_92 <= 32'h0;
      v0_93 <= 32'h0;
      v0_94 <= 32'h0;
      v0_95 <= 32'h0;
      v0_96 <= 32'h0;
      v0_97 <= 32'h0;
      v0_98 <= 32'h0;
      v0_99 <= 32'h0;
      v0_100 <= 32'h0;
      v0_101 <= 32'h0;
      v0_102 <= 32'h0;
      v0_103 <= 32'h0;
      v0_104 <= 32'h0;
      v0_105 <= 32'h0;
      v0_106 <= 32'h0;
      v0_107 <= 32'h0;
      v0_108 <= 32'h0;
      v0_109 <= 32'h0;
      v0_110 <= 32'h0;
      v0_111 <= 32'h0;
      v0_112 <= 32'h0;
      v0_113 <= 32'h0;
      v0_114 <= 32'h0;
      v0_115 <= 32'h0;
      v0_116 <= 32'h0;
      v0_117 <= 32'h0;
      v0_118 <= 32'h0;
      v0_119 <= 32'h0;
      v0_120 <= 32'h0;
      v0_121 <= 32'h0;
      v0_122 <= 32'h0;
      v0_123 <= 32'h0;
      v0_124 <= 32'h0;
      v0_125 <= 32'h0;
      v0_126 <= 32'h0;
      v0_127 <= 32'h0;
      v0_128 <= 32'h0;
      v0_129 <= 32'h0;
      v0_130 <= 32'h0;
      v0_131 <= 32'h0;
      v0_132 <= 32'h0;
      v0_133 <= 32'h0;
      v0_134 <= 32'h0;
      v0_135 <= 32'h0;
      v0_136 <= 32'h0;
      v0_137 <= 32'h0;
      v0_138 <= 32'h0;
      v0_139 <= 32'h0;
      v0_140 <= 32'h0;
      v0_141 <= 32'h0;
      v0_142 <= 32'h0;
      v0_143 <= 32'h0;
      v0_144 <= 32'h0;
      v0_145 <= 32'h0;
      v0_146 <= 32'h0;
      v0_147 <= 32'h0;
      v0_148 <= 32'h0;
      v0_149 <= 32'h0;
      v0_150 <= 32'h0;
      v0_151 <= 32'h0;
      v0_152 <= 32'h0;
      v0_153 <= 32'h0;
      v0_154 <= 32'h0;
      v0_155 <= 32'h0;
      v0_156 <= 32'h0;
      v0_157 <= 32'h0;
      v0_158 <= 32'h0;
      v0_159 <= 32'h0;
      v0_160 <= 32'h0;
      v0_161 <= 32'h0;
      v0_162 <= 32'h0;
      v0_163 <= 32'h0;
      v0_164 <= 32'h0;
      v0_165 <= 32'h0;
      v0_166 <= 32'h0;
      v0_167 <= 32'h0;
      v0_168 <= 32'h0;
      v0_169 <= 32'h0;
      v0_170 <= 32'h0;
      v0_171 <= 32'h0;
      v0_172 <= 32'h0;
      v0_173 <= 32'h0;
      v0_174 <= 32'h0;
      v0_175 <= 32'h0;
      v0_176 <= 32'h0;
      v0_177 <= 32'h0;
      v0_178 <= 32'h0;
      v0_179 <= 32'h0;
      v0_180 <= 32'h0;
      v0_181 <= 32'h0;
      v0_182 <= 32'h0;
      v0_183 <= 32'h0;
      v0_184 <= 32'h0;
      v0_185 <= 32'h0;
      v0_186 <= 32'h0;
      v0_187 <= 32'h0;
      v0_188 <= 32'h0;
      v0_189 <= 32'h0;
      v0_190 <= 32'h0;
      v0_191 <= 32'h0;
      v0_192 <= 32'h0;
      v0_193 <= 32'h0;
      v0_194 <= 32'h0;
      v0_195 <= 32'h0;
      v0_196 <= 32'h0;
      v0_197 <= 32'h0;
      v0_198 <= 32'h0;
      v0_199 <= 32'h0;
      v0_200 <= 32'h0;
      v0_201 <= 32'h0;
      v0_202 <= 32'h0;
      v0_203 <= 32'h0;
      v0_204 <= 32'h0;
      v0_205 <= 32'h0;
      v0_206 <= 32'h0;
      v0_207 <= 32'h0;
      v0_208 <= 32'h0;
      v0_209 <= 32'h0;
      v0_210 <= 32'h0;
      v0_211 <= 32'h0;
      v0_212 <= 32'h0;
      v0_213 <= 32'h0;
      v0_214 <= 32'h0;
      v0_215 <= 32'h0;
      v0_216 <= 32'h0;
      v0_217 <= 32'h0;
      v0_218 <= 32'h0;
      v0_219 <= 32'h0;
      v0_220 <= 32'h0;
      v0_221 <= 32'h0;
      v0_222 <= 32'h0;
      v0_223 <= 32'h0;
      v0_224 <= 32'h0;
      v0_225 <= 32'h0;
      v0_226 <= 32'h0;
      v0_227 <= 32'h0;
      v0_228 <= 32'h0;
      v0_229 <= 32'h0;
      v0_230 <= 32'h0;
      v0_231 <= 32'h0;
      v0_232 <= 32'h0;
      v0_233 <= 32'h0;
      v0_234 <= 32'h0;
      v0_235 <= 32'h0;
      v0_236 <= 32'h0;
      v0_237 <= 32'h0;
      v0_238 <= 32'h0;
      v0_239 <= 32'h0;
      v0_240 <= 32'h0;
      v0_241 <= 32'h0;
      v0_242 <= 32'h0;
      v0_243 <= 32'h0;
      v0_244 <= 32'h0;
      v0_245 <= 32'h0;
      v0_246 <= 32'h0;
      v0_247 <= 32'h0;
      v0_248 <= 32'h0;
      v0_249 <= 32'h0;
      v0_250 <= 32'h0;
      v0_251 <= 32'h0;
      v0_252 <= 32'h0;
      v0_253 <= 32'h0;
      v0_254 <= 32'h0;
      v0_255 <= 32'h0;
      v0_256 <= 32'h0;
      v0_257 <= 32'h0;
      v0_258 <= 32'h0;
      v0_259 <= 32'h0;
      v0_260 <= 32'h0;
      v0_261 <= 32'h0;
      v0_262 <= 32'h0;
      v0_263 <= 32'h0;
      v0_264 <= 32'h0;
      v0_265 <= 32'h0;
      v0_266 <= 32'h0;
      v0_267 <= 32'h0;
      v0_268 <= 32'h0;
      v0_269 <= 32'h0;
      v0_270 <= 32'h0;
      v0_271 <= 32'h0;
      v0_272 <= 32'h0;
      v0_273 <= 32'h0;
      v0_274 <= 32'h0;
      v0_275 <= 32'h0;
      v0_276 <= 32'h0;
      v0_277 <= 32'h0;
      v0_278 <= 32'h0;
      v0_279 <= 32'h0;
      v0_280 <= 32'h0;
      v0_281 <= 32'h0;
      v0_282 <= 32'h0;
      v0_283 <= 32'h0;
      v0_284 <= 32'h0;
      v0_285 <= 32'h0;
      v0_286 <= 32'h0;
      v0_287 <= 32'h0;
      v0_288 <= 32'h0;
      v0_289 <= 32'h0;
      v0_290 <= 32'h0;
      v0_291 <= 32'h0;
      v0_292 <= 32'h0;
      v0_293 <= 32'h0;
      v0_294 <= 32'h0;
      v0_295 <= 32'h0;
      v0_296 <= 32'h0;
      v0_297 <= 32'h0;
      v0_298 <= 32'h0;
      v0_299 <= 32'h0;
      v0_300 <= 32'h0;
      v0_301 <= 32'h0;
      v0_302 <= 32'h0;
      v0_303 <= 32'h0;
      v0_304 <= 32'h0;
      v0_305 <= 32'h0;
      v0_306 <= 32'h0;
      v0_307 <= 32'h0;
      v0_308 <= 32'h0;
      v0_309 <= 32'h0;
      v0_310 <= 32'h0;
      v0_311 <= 32'h0;
      v0_312 <= 32'h0;
      v0_313 <= 32'h0;
      v0_314 <= 32'h0;
      v0_315 <= 32'h0;
      v0_316 <= 32'h0;
      v0_317 <= 32'h0;
      v0_318 <= 32'h0;
      v0_319 <= 32'h0;
      v0_320 <= 32'h0;
      v0_321 <= 32'h0;
      v0_322 <= 32'h0;
      v0_323 <= 32'h0;
      v0_324 <= 32'h0;
      v0_325 <= 32'h0;
      v0_326 <= 32'h0;
      v0_327 <= 32'h0;
      v0_328 <= 32'h0;
      v0_329 <= 32'h0;
      v0_330 <= 32'h0;
      v0_331 <= 32'h0;
      v0_332 <= 32'h0;
      v0_333 <= 32'h0;
      v0_334 <= 32'h0;
      v0_335 <= 32'h0;
      v0_336 <= 32'h0;
      v0_337 <= 32'h0;
      v0_338 <= 32'h0;
      v0_339 <= 32'h0;
      v0_340 <= 32'h0;
      v0_341 <= 32'h0;
      v0_342 <= 32'h0;
      v0_343 <= 32'h0;
      v0_344 <= 32'h0;
      v0_345 <= 32'h0;
      v0_346 <= 32'h0;
      v0_347 <= 32'h0;
      v0_348 <= 32'h0;
      v0_349 <= 32'h0;
      v0_350 <= 32'h0;
      v0_351 <= 32'h0;
      v0_352 <= 32'h0;
      v0_353 <= 32'h0;
      v0_354 <= 32'h0;
      v0_355 <= 32'h0;
      v0_356 <= 32'h0;
      v0_357 <= 32'h0;
      v0_358 <= 32'h0;
      v0_359 <= 32'h0;
      v0_360 <= 32'h0;
      v0_361 <= 32'h0;
      v0_362 <= 32'h0;
      v0_363 <= 32'h0;
      v0_364 <= 32'h0;
      v0_365 <= 32'h0;
      v0_366 <= 32'h0;
      v0_367 <= 32'h0;
      v0_368 <= 32'h0;
      v0_369 <= 32'h0;
      v0_370 <= 32'h0;
      v0_371 <= 32'h0;
      v0_372 <= 32'h0;
      v0_373 <= 32'h0;
      v0_374 <= 32'h0;
      v0_375 <= 32'h0;
      v0_376 <= 32'h0;
      v0_377 <= 32'h0;
      v0_378 <= 32'h0;
      v0_379 <= 32'h0;
      v0_380 <= 32'h0;
      v0_381 <= 32'h0;
      v0_382 <= 32'h0;
      v0_383 <= 32'h0;
      v0_384 <= 32'h0;
      v0_385 <= 32'h0;
      v0_386 <= 32'h0;
      v0_387 <= 32'h0;
      v0_388 <= 32'h0;
      v0_389 <= 32'h0;
      v0_390 <= 32'h0;
      v0_391 <= 32'h0;
      v0_392 <= 32'h0;
      v0_393 <= 32'h0;
      v0_394 <= 32'h0;
      v0_395 <= 32'h0;
      v0_396 <= 32'h0;
      v0_397 <= 32'h0;
      v0_398 <= 32'h0;
      v0_399 <= 32'h0;
      v0_400 <= 32'h0;
      v0_401 <= 32'h0;
      v0_402 <= 32'h0;
      v0_403 <= 32'h0;
      v0_404 <= 32'h0;
      v0_405 <= 32'h0;
      v0_406 <= 32'h0;
      v0_407 <= 32'h0;
      v0_408 <= 32'h0;
      v0_409 <= 32'h0;
      v0_410 <= 32'h0;
      v0_411 <= 32'h0;
      v0_412 <= 32'h0;
      v0_413 <= 32'h0;
      v0_414 <= 32'h0;
      v0_415 <= 32'h0;
      v0_416 <= 32'h0;
      v0_417 <= 32'h0;
      v0_418 <= 32'h0;
      v0_419 <= 32'h0;
      v0_420 <= 32'h0;
      v0_421 <= 32'h0;
      v0_422 <= 32'h0;
      v0_423 <= 32'h0;
      v0_424 <= 32'h0;
      v0_425 <= 32'h0;
      v0_426 <= 32'h0;
      v0_427 <= 32'h0;
      v0_428 <= 32'h0;
      v0_429 <= 32'h0;
      v0_430 <= 32'h0;
      v0_431 <= 32'h0;
      v0_432 <= 32'h0;
      v0_433 <= 32'h0;
      v0_434 <= 32'h0;
      v0_435 <= 32'h0;
      v0_436 <= 32'h0;
      v0_437 <= 32'h0;
      v0_438 <= 32'h0;
      v0_439 <= 32'h0;
      v0_440 <= 32'h0;
      v0_441 <= 32'h0;
      v0_442 <= 32'h0;
      v0_443 <= 32'h0;
      v0_444 <= 32'h0;
      v0_445 <= 32'h0;
      v0_446 <= 32'h0;
      v0_447 <= 32'h0;
      v0_448 <= 32'h0;
      v0_449 <= 32'h0;
      v0_450 <= 32'h0;
      v0_451 <= 32'h0;
      v0_452 <= 32'h0;
      v0_453 <= 32'h0;
      v0_454 <= 32'h0;
      v0_455 <= 32'h0;
      v0_456 <= 32'h0;
      v0_457 <= 32'h0;
      v0_458 <= 32'h0;
      v0_459 <= 32'h0;
      v0_460 <= 32'h0;
      v0_461 <= 32'h0;
      v0_462 <= 32'h0;
      v0_463 <= 32'h0;
      v0_464 <= 32'h0;
      v0_465 <= 32'h0;
      v0_466 <= 32'h0;
      v0_467 <= 32'h0;
      v0_468 <= 32'h0;
      v0_469 <= 32'h0;
      v0_470 <= 32'h0;
      v0_471 <= 32'h0;
      v0_472 <= 32'h0;
      v0_473 <= 32'h0;
      v0_474 <= 32'h0;
      v0_475 <= 32'h0;
      v0_476 <= 32'h0;
      v0_477 <= 32'h0;
      v0_478 <= 32'h0;
      v0_479 <= 32'h0;
      v0_480 <= 32'h0;
      v0_481 <= 32'h0;
      v0_482 <= 32'h0;
      v0_483 <= 32'h0;
      v0_484 <= 32'h0;
      v0_485 <= 32'h0;
      v0_486 <= 32'h0;
      v0_487 <= 32'h0;
      v0_488 <= 32'h0;
      v0_489 <= 32'h0;
      v0_490 <= 32'h0;
      v0_491 <= 32'h0;
      v0_492 <= 32'h0;
      v0_493 <= 32'h0;
      v0_494 <= 32'h0;
      v0_495 <= 32'h0;
      v0_496 <= 32'h0;
      v0_497 <= 32'h0;
      v0_498 <= 32'h0;
      v0_499 <= 32'h0;
      v0_500 <= 32'h0;
      v0_501 <= 32'h0;
      v0_502 <= 32'h0;
      v0_503 <= 32'h0;
      v0_504 <= 32'h0;
      v0_505 <= 32'h0;
      v0_506 <= 32'h0;
      v0_507 <= 32'h0;
      v0_508 <= 32'h0;
      v0_509 <= 32'h0;
      v0_510 <= 32'h0;
      v0_511 <= 32'h0;
      v0_512 <= 32'h0;
      v0_513 <= 32'h0;
      v0_514 <= 32'h0;
      v0_515 <= 32'h0;
      v0_516 <= 32'h0;
      v0_517 <= 32'h0;
      v0_518 <= 32'h0;
      v0_519 <= 32'h0;
      v0_520 <= 32'h0;
      v0_521 <= 32'h0;
      v0_522 <= 32'h0;
      v0_523 <= 32'h0;
      v0_524 <= 32'h0;
      v0_525 <= 32'h0;
      v0_526 <= 32'h0;
      v0_527 <= 32'h0;
      v0_528 <= 32'h0;
      v0_529 <= 32'h0;
      v0_530 <= 32'h0;
      v0_531 <= 32'h0;
      v0_532 <= 32'h0;
      v0_533 <= 32'h0;
      v0_534 <= 32'h0;
      v0_535 <= 32'h0;
      v0_536 <= 32'h0;
      v0_537 <= 32'h0;
      v0_538 <= 32'h0;
      v0_539 <= 32'h0;
      v0_540 <= 32'h0;
      v0_541 <= 32'h0;
      v0_542 <= 32'h0;
      v0_543 <= 32'h0;
      v0_544 <= 32'h0;
      v0_545 <= 32'h0;
      v0_546 <= 32'h0;
      v0_547 <= 32'h0;
      v0_548 <= 32'h0;
      v0_549 <= 32'h0;
      v0_550 <= 32'h0;
      v0_551 <= 32'h0;
      v0_552 <= 32'h0;
      v0_553 <= 32'h0;
      v0_554 <= 32'h0;
      v0_555 <= 32'h0;
      v0_556 <= 32'h0;
      v0_557 <= 32'h0;
      v0_558 <= 32'h0;
      v0_559 <= 32'h0;
      v0_560 <= 32'h0;
      v0_561 <= 32'h0;
      v0_562 <= 32'h0;
      v0_563 <= 32'h0;
      v0_564 <= 32'h0;
      v0_565 <= 32'h0;
      v0_566 <= 32'h0;
      v0_567 <= 32'h0;
      v0_568 <= 32'h0;
      v0_569 <= 32'h0;
      v0_570 <= 32'h0;
      v0_571 <= 32'h0;
      v0_572 <= 32'h0;
      v0_573 <= 32'h0;
      v0_574 <= 32'h0;
      v0_575 <= 32'h0;
      v0_576 <= 32'h0;
      v0_577 <= 32'h0;
      v0_578 <= 32'h0;
      v0_579 <= 32'h0;
      v0_580 <= 32'h0;
      v0_581 <= 32'h0;
      v0_582 <= 32'h0;
      v0_583 <= 32'h0;
      v0_584 <= 32'h0;
      v0_585 <= 32'h0;
      v0_586 <= 32'h0;
      v0_587 <= 32'h0;
      v0_588 <= 32'h0;
      v0_589 <= 32'h0;
      v0_590 <= 32'h0;
      v0_591 <= 32'h0;
      v0_592 <= 32'h0;
      v0_593 <= 32'h0;
      v0_594 <= 32'h0;
      v0_595 <= 32'h0;
      v0_596 <= 32'h0;
      v0_597 <= 32'h0;
      v0_598 <= 32'h0;
      v0_599 <= 32'h0;
      v0_600 <= 32'h0;
      v0_601 <= 32'h0;
      v0_602 <= 32'h0;
      v0_603 <= 32'h0;
      v0_604 <= 32'h0;
      v0_605 <= 32'h0;
      v0_606 <= 32'h0;
      v0_607 <= 32'h0;
      v0_608 <= 32'h0;
      v0_609 <= 32'h0;
      v0_610 <= 32'h0;
      v0_611 <= 32'h0;
      v0_612 <= 32'h0;
      v0_613 <= 32'h0;
      v0_614 <= 32'h0;
      v0_615 <= 32'h0;
      v0_616 <= 32'h0;
      v0_617 <= 32'h0;
      v0_618 <= 32'h0;
      v0_619 <= 32'h0;
      v0_620 <= 32'h0;
      v0_621 <= 32'h0;
      v0_622 <= 32'h0;
      v0_623 <= 32'h0;
      v0_624 <= 32'h0;
      v0_625 <= 32'h0;
      v0_626 <= 32'h0;
      v0_627 <= 32'h0;
      v0_628 <= 32'h0;
      v0_629 <= 32'h0;
      v0_630 <= 32'h0;
      v0_631 <= 32'h0;
      v0_632 <= 32'h0;
      v0_633 <= 32'h0;
      v0_634 <= 32'h0;
      v0_635 <= 32'h0;
      v0_636 <= 32'h0;
      v0_637 <= 32'h0;
      v0_638 <= 32'h0;
      v0_639 <= 32'h0;
      v0_640 <= 32'h0;
      v0_641 <= 32'h0;
      v0_642 <= 32'h0;
      v0_643 <= 32'h0;
      v0_644 <= 32'h0;
      v0_645 <= 32'h0;
      v0_646 <= 32'h0;
      v0_647 <= 32'h0;
      v0_648 <= 32'h0;
      v0_649 <= 32'h0;
      v0_650 <= 32'h0;
      v0_651 <= 32'h0;
      v0_652 <= 32'h0;
      v0_653 <= 32'h0;
      v0_654 <= 32'h0;
      v0_655 <= 32'h0;
      v0_656 <= 32'h0;
      v0_657 <= 32'h0;
      v0_658 <= 32'h0;
      v0_659 <= 32'h0;
      v0_660 <= 32'h0;
      v0_661 <= 32'h0;
      v0_662 <= 32'h0;
      v0_663 <= 32'h0;
      v0_664 <= 32'h0;
      v0_665 <= 32'h0;
      v0_666 <= 32'h0;
      v0_667 <= 32'h0;
      v0_668 <= 32'h0;
      v0_669 <= 32'h0;
      v0_670 <= 32'h0;
      v0_671 <= 32'h0;
      v0_672 <= 32'h0;
      v0_673 <= 32'h0;
      v0_674 <= 32'h0;
      v0_675 <= 32'h0;
      v0_676 <= 32'h0;
      v0_677 <= 32'h0;
      v0_678 <= 32'h0;
      v0_679 <= 32'h0;
      v0_680 <= 32'h0;
      v0_681 <= 32'h0;
      v0_682 <= 32'h0;
      v0_683 <= 32'h0;
      v0_684 <= 32'h0;
      v0_685 <= 32'h0;
      v0_686 <= 32'h0;
      v0_687 <= 32'h0;
      v0_688 <= 32'h0;
      v0_689 <= 32'h0;
      v0_690 <= 32'h0;
      v0_691 <= 32'h0;
      v0_692 <= 32'h0;
      v0_693 <= 32'h0;
      v0_694 <= 32'h0;
      v0_695 <= 32'h0;
      v0_696 <= 32'h0;
      v0_697 <= 32'h0;
      v0_698 <= 32'h0;
      v0_699 <= 32'h0;
      v0_700 <= 32'h0;
      v0_701 <= 32'h0;
      v0_702 <= 32'h0;
      v0_703 <= 32'h0;
      v0_704 <= 32'h0;
      v0_705 <= 32'h0;
      v0_706 <= 32'h0;
      v0_707 <= 32'h0;
      v0_708 <= 32'h0;
      v0_709 <= 32'h0;
      v0_710 <= 32'h0;
      v0_711 <= 32'h0;
      v0_712 <= 32'h0;
      v0_713 <= 32'h0;
      v0_714 <= 32'h0;
      v0_715 <= 32'h0;
      v0_716 <= 32'h0;
      v0_717 <= 32'h0;
      v0_718 <= 32'h0;
      v0_719 <= 32'h0;
      v0_720 <= 32'h0;
      v0_721 <= 32'h0;
      v0_722 <= 32'h0;
      v0_723 <= 32'h0;
      v0_724 <= 32'h0;
      v0_725 <= 32'h0;
      v0_726 <= 32'h0;
      v0_727 <= 32'h0;
      v0_728 <= 32'h0;
      v0_729 <= 32'h0;
      v0_730 <= 32'h0;
      v0_731 <= 32'h0;
      v0_732 <= 32'h0;
      v0_733 <= 32'h0;
      v0_734 <= 32'h0;
      v0_735 <= 32'h0;
      v0_736 <= 32'h0;
      v0_737 <= 32'h0;
      v0_738 <= 32'h0;
      v0_739 <= 32'h0;
      v0_740 <= 32'h0;
      v0_741 <= 32'h0;
      v0_742 <= 32'h0;
      v0_743 <= 32'h0;
      v0_744 <= 32'h0;
      v0_745 <= 32'h0;
      v0_746 <= 32'h0;
      v0_747 <= 32'h0;
      v0_748 <= 32'h0;
      v0_749 <= 32'h0;
      v0_750 <= 32'h0;
      v0_751 <= 32'h0;
      v0_752 <= 32'h0;
      v0_753 <= 32'h0;
      v0_754 <= 32'h0;
      v0_755 <= 32'h0;
      v0_756 <= 32'h0;
      v0_757 <= 32'h0;
      v0_758 <= 32'h0;
      v0_759 <= 32'h0;
      v0_760 <= 32'h0;
      v0_761 <= 32'h0;
      v0_762 <= 32'h0;
      v0_763 <= 32'h0;
      v0_764 <= 32'h0;
      v0_765 <= 32'h0;
      v0_766 <= 32'h0;
      v0_767 <= 32'h0;
      v0_768 <= 32'h0;
      v0_769 <= 32'h0;
      v0_770 <= 32'h0;
      v0_771 <= 32'h0;
      v0_772 <= 32'h0;
      v0_773 <= 32'h0;
      v0_774 <= 32'h0;
      v0_775 <= 32'h0;
      v0_776 <= 32'h0;
      v0_777 <= 32'h0;
      v0_778 <= 32'h0;
      v0_779 <= 32'h0;
      v0_780 <= 32'h0;
      v0_781 <= 32'h0;
      v0_782 <= 32'h0;
      v0_783 <= 32'h0;
      v0_784 <= 32'h0;
      v0_785 <= 32'h0;
      v0_786 <= 32'h0;
      v0_787 <= 32'h0;
      v0_788 <= 32'h0;
      v0_789 <= 32'h0;
      v0_790 <= 32'h0;
      v0_791 <= 32'h0;
      v0_792 <= 32'h0;
      v0_793 <= 32'h0;
      v0_794 <= 32'h0;
      v0_795 <= 32'h0;
      v0_796 <= 32'h0;
      v0_797 <= 32'h0;
      v0_798 <= 32'h0;
      v0_799 <= 32'h0;
      v0_800 <= 32'h0;
      v0_801 <= 32'h0;
      v0_802 <= 32'h0;
      v0_803 <= 32'h0;
      v0_804 <= 32'h0;
      v0_805 <= 32'h0;
      v0_806 <= 32'h0;
      v0_807 <= 32'h0;
      v0_808 <= 32'h0;
      v0_809 <= 32'h0;
      v0_810 <= 32'h0;
      v0_811 <= 32'h0;
      v0_812 <= 32'h0;
      v0_813 <= 32'h0;
      v0_814 <= 32'h0;
      v0_815 <= 32'h0;
      v0_816 <= 32'h0;
      v0_817 <= 32'h0;
      v0_818 <= 32'h0;
      v0_819 <= 32'h0;
      v0_820 <= 32'h0;
      v0_821 <= 32'h0;
      v0_822 <= 32'h0;
      v0_823 <= 32'h0;
      v0_824 <= 32'h0;
      v0_825 <= 32'h0;
      v0_826 <= 32'h0;
      v0_827 <= 32'h0;
      v0_828 <= 32'h0;
      v0_829 <= 32'h0;
      v0_830 <= 32'h0;
      v0_831 <= 32'h0;
      v0_832 <= 32'h0;
      v0_833 <= 32'h0;
      v0_834 <= 32'h0;
      v0_835 <= 32'h0;
      v0_836 <= 32'h0;
      v0_837 <= 32'h0;
      v0_838 <= 32'h0;
      v0_839 <= 32'h0;
      v0_840 <= 32'h0;
      v0_841 <= 32'h0;
      v0_842 <= 32'h0;
      v0_843 <= 32'h0;
      v0_844 <= 32'h0;
      v0_845 <= 32'h0;
      v0_846 <= 32'h0;
      v0_847 <= 32'h0;
      v0_848 <= 32'h0;
      v0_849 <= 32'h0;
      v0_850 <= 32'h0;
      v0_851 <= 32'h0;
      v0_852 <= 32'h0;
      v0_853 <= 32'h0;
      v0_854 <= 32'h0;
      v0_855 <= 32'h0;
      v0_856 <= 32'h0;
      v0_857 <= 32'h0;
      v0_858 <= 32'h0;
      v0_859 <= 32'h0;
      v0_860 <= 32'h0;
      v0_861 <= 32'h0;
      v0_862 <= 32'h0;
      v0_863 <= 32'h0;
      v0_864 <= 32'h0;
      v0_865 <= 32'h0;
      v0_866 <= 32'h0;
      v0_867 <= 32'h0;
      v0_868 <= 32'h0;
      v0_869 <= 32'h0;
      v0_870 <= 32'h0;
      v0_871 <= 32'h0;
      v0_872 <= 32'h0;
      v0_873 <= 32'h0;
      v0_874 <= 32'h0;
      v0_875 <= 32'h0;
      v0_876 <= 32'h0;
      v0_877 <= 32'h0;
      v0_878 <= 32'h0;
      v0_879 <= 32'h0;
      v0_880 <= 32'h0;
      v0_881 <= 32'h0;
      v0_882 <= 32'h0;
      v0_883 <= 32'h0;
      v0_884 <= 32'h0;
      v0_885 <= 32'h0;
      v0_886 <= 32'h0;
      v0_887 <= 32'h0;
      v0_888 <= 32'h0;
      v0_889 <= 32'h0;
      v0_890 <= 32'h0;
      v0_891 <= 32'h0;
      v0_892 <= 32'h0;
      v0_893 <= 32'h0;
      v0_894 <= 32'h0;
      v0_895 <= 32'h0;
      v0_896 <= 32'h0;
      v0_897 <= 32'h0;
      v0_898 <= 32'h0;
      v0_899 <= 32'h0;
      v0_900 <= 32'h0;
      v0_901 <= 32'h0;
      v0_902 <= 32'h0;
      v0_903 <= 32'h0;
      v0_904 <= 32'h0;
      v0_905 <= 32'h0;
      v0_906 <= 32'h0;
      v0_907 <= 32'h0;
      v0_908 <= 32'h0;
      v0_909 <= 32'h0;
      v0_910 <= 32'h0;
      v0_911 <= 32'h0;
      v0_912 <= 32'h0;
      v0_913 <= 32'h0;
      v0_914 <= 32'h0;
      v0_915 <= 32'h0;
      v0_916 <= 32'h0;
      v0_917 <= 32'h0;
      v0_918 <= 32'h0;
      v0_919 <= 32'h0;
      v0_920 <= 32'h0;
      v0_921 <= 32'h0;
      v0_922 <= 32'h0;
      v0_923 <= 32'h0;
      v0_924 <= 32'h0;
      v0_925 <= 32'h0;
      v0_926 <= 32'h0;
      v0_927 <= 32'h0;
      v0_928 <= 32'h0;
      v0_929 <= 32'h0;
      v0_930 <= 32'h0;
      v0_931 <= 32'h0;
      v0_932 <= 32'h0;
      v0_933 <= 32'h0;
      v0_934 <= 32'h0;
      v0_935 <= 32'h0;
      v0_936 <= 32'h0;
      v0_937 <= 32'h0;
      v0_938 <= 32'h0;
      v0_939 <= 32'h0;
      v0_940 <= 32'h0;
      v0_941 <= 32'h0;
      v0_942 <= 32'h0;
      v0_943 <= 32'h0;
      v0_944 <= 32'h0;
      v0_945 <= 32'h0;
      v0_946 <= 32'h0;
      v0_947 <= 32'h0;
      v0_948 <= 32'h0;
      v0_949 <= 32'h0;
      v0_950 <= 32'h0;
      v0_951 <= 32'h0;
      v0_952 <= 32'h0;
      v0_953 <= 32'h0;
      v0_954 <= 32'h0;
      v0_955 <= 32'h0;
      v0_956 <= 32'h0;
      v0_957 <= 32'h0;
      v0_958 <= 32'h0;
      v0_959 <= 32'h0;
      v0_960 <= 32'h0;
      v0_961 <= 32'h0;
      v0_962 <= 32'h0;
      v0_963 <= 32'h0;
      v0_964 <= 32'h0;
      v0_965 <= 32'h0;
      v0_966 <= 32'h0;
      v0_967 <= 32'h0;
      v0_968 <= 32'h0;
      v0_969 <= 32'h0;
      v0_970 <= 32'h0;
      v0_971 <= 32'h0;
      v0_972 <= 32'h0;
      v0_973 <= 32'h0;
      v0_974 <= 32'h0;
      v0_975 <= 32'h0;
      v0_976 <= 32'h0;
      v0_977 <= 32'h0;
      v0_978 <= 32'h0;
      v0_979 <= 32'h0;
      v0_980 <= 32'h0;
      v0_981 <= 32'h0;
      v0_982 <= 32'h0;
      v0_983 <= 32'h0;
      v0_984 <= 32'h0;
      v0_985 <= 32'h0;
      v0_986 <= 32'h0;
      v0_987 <= 32'h0;
      v0_988 <= 32'h0;
      v0_989 <= 32'h0;
      v0_990 <= 32'h0;
      v0_991 <= 32'h0;
      v0_992 <= 32'h0;
      v0_993 <= 32'h0;
      v0_994 <= 32'h0;
      v0_995 <= 32'h0;
      v0_996 <= 32'h0;
      v0_997 <= 32'h0;
      v0_998 <= 32'h0;
      v0_999 <= 32'h0;
      v0_1000 <= 32'h0;
      v0_1001 <= 32'h0;
      v0_1002 <= 32'h0;
      v0_1003 <= 32'h0;
      v0_1004 <= 32'h0;
      v0_1005 <= 32'h0;
      v0_1006 <= 32'h0;
      v0_1007 <= 32'h0;
      v0_1008 <= 32'h0;
      v0_1009 <= 32'h0;
      v0_1010 <= 32'h0;
      v0_1011 <= 32'h0;
      v0_1012 <= 32'h0;
      v0_1013 <= 32'h0;
      v0_1014 <= 32'h0;
      v0_1015 <= 32'h0;
      v0_1016 <= 32'h0;
      v0_1017 <= 32'h0;
      v0_1018 <= 32'h0;
      v0_1019 <= 32'h0;
      v0_1020 <= 32'h0;
      v0_1021 <= 32'h0;
      v0_1022 <= 32'h0;
      v0_1023 <= 32'h0;
      v0_1024 <= 32'h0;
      v0_1025 <= 32'h0;
      v0_1026 <= 32'h0;
      v0_1027 <= 32'h0;
      v0_1028 <= 32'h0;
      v0_1029 <= 32'h0;
      v0_1030 <= 32'h0;
      v0_1031 <= 32'h0;
      v0_1032 <= 32'h0;
      v0_1033 <= 32'h0;
      v0_1034 <= 32'h0;
      v0_1035 <= 32'h0;
      v0_1036 <= 32'h0;
      v0_1037 <= 32'h0;
      v0_1038 <= 32'h0;
      v0_1039 <= 32'h0;
      v0_1040 <= 32'h0;
      v0_1041 <= 32'h0;
      v0_1042 <= 32'h0;
      v0_1043 <= 32'h0;
      v0_1044 <= 32'h0;
      v0_1045 <= 32'h0;
      v0_1046 <= 32'h0;
      v0_1047 <= 32'h0;
      v0_1048 <= 32'h0;
      v0_1049 <= 32'h0;
      v0_1050 <= 32'h0;
      v0_1051 <= 32'h0;
      v0_1052 <= 32'h0;
      v0_1053 <= 32'h0;
      v0_1054 <= 32'h0;
      v0_1055 <= 32'h0;
      v0_1056 <= 32'h0;
      v0_1057 <= 32'h0;
      v0_1058 <= 32'h0;
      v0_1059 <= 32'h0;
      v0_1060 <= 32'h0;
      v0_1061 <= 32'h0;
      v0_1062 <= 32'h0;
      v0_1063 <= 32'h0;
      v0_1064 <= 32'h0;
      v0_1065 <= 32'h0;
      v0_1066 <= 32'h0;
      v0_1067 <= 32'h0;
      v0_1068 <= 32'h0;
      v0_1069 <= 32'h0;
      v0_1070 <= 32'h0;
      v0_1071 <= 32'h0;
      v0_1072 <= 32'h0;
      v0_1073 <= 32'h0;
      v0_1074 <= 32'h0;
      v0_1075 <= 32'h0;
      v0_1076 <= 32'h0;
      v0_1077 <= 32'h0;
      v0_1078 <= 32'h0;
      v0_1079 <= 32'h0;
      v0_1080 <= 32'h0;
      v0_1081 <= 32'h0;
      v0_1082 <= 32'h0;
      v0_1083 <= 32'h0;
      v0_1084 <= 32'h0;
      v0_1085 <= 32'h0;
      v0_1086 <= 32'h0;
      v0_1087 <= 32'h0;
      v0_1088 <= 32'h0;
      v0_1089 <= 32'h0;
      v0_1090 <= 32'h0;
      v0_1091 <= 32'h0;
      v0_1092 <= 32'h0;
      v0_1093 <= 32'h0;
      v0_1094 <= 32'h0;
      v0_1095 <= 32'h0;
      v0_1096 <= 32'h0;
      v0_1097 <= 32'h0;
      v0_1098 <= 32'h0;
      v0_1099 <= 32'h0;
      v0_1100 <= 32'h0;
      v0_1101 <= 32'h0;
      v0_1102 <= 32'h0;
      v0_1103 <= 32'h0;
      v0_1104 <= 32'h0;
      v0_1105 <= 32'h0;
      v0_1106 <= 32'h0;
      v0_1107 <= 32'h0;
      v0_1108 <= 32'h0;
      v0_1109 <= 32'h0;
      v0_1110 <= 32'h0;
      v0_1111 <= 32'h0;
      v0_1112 <= 32'h0;
      v0_1113 <= 32'h0;
      v0_1114 <= 32'h0;
      v0_1115 <= 32'h0;
      v0_1116 <= 32'h0;
      v0_1117 <= 32'h0;
      v0_1118 <= 32'h0;
      v0_1119 <= 32'h0;
      v0_1120 <= 32'h0;
      v0_1121 <= 32'h0;
      v0_1122 <= 32'h0;
      v0_1123 <= 32'h0;
      v0_1124 <= 32'h0;
      v0_1125 <= 32'h0;
      v0_1126 <= 32'h0;
      v0_1127 <= 32'h0;
      v0_1128 <= 32'h0;
      v0_1129 <= 32'h0;
      v0_1130 <= 32'h0;
      v0_1131 <= 32'h0;
      v0_1132 <= 32'h0;
      v0_1133 <= 32'h0;
      v0_1134 <= 32'h0;
      v0_1135 <= 32'h0;
      v0_1136 <= 32'h0;
      v0_1137 <= 32'h0;
      v0_1138 <= 32'h0;
      v0_1139 <= 32'h0;
      v0_1140 <= 32'h0;
      v0_1141 <= 32'h0;
      v0_1142 <= 32'h0;
      v0_1143 <= 32'h0;
      v0_1144 <= 32'h0;
      v0_1145 <= 32'h0;
      v0_1146 <= 32'h0;
      v0_1147 <= 32'h0;
      v0_1148 <= 32'h0;
      v0_1149 <= 32'h0;
      v0_1150 <= 32'h0;
      v0_1151 <= 32'h0;
      v0_1152 <= 32'h0;
      v0_1153 <= 32'h0;
      v0_1154 <= 32'h0;
      v0_1155 <= 32'h0;
      v0_1156 <= 32'h0;
      v0_1157 <= 32'h0;
      v0_1158 <= 32'h0;
      v0_1159 <= 32'h0;
      v0_1160 <= 32'h0;
      v0_1161 <= 32'h0;
      v0_1162 <= 32'h0;
      v0_1163 <= 32'h0;
      v0_1164 <= 32'h0;
      v0_1165 <= 32'h0;
      v0_1166 <= 32'h0;
      v0_1167 <= 32'h0;
      v0_1168 <= 32'h0;
      v0_1169 <= 32'h0;
      v0_1170 <= 32'h0;
      v0_1171 <= 32'h0;
      v0_1172 <= 32'h0;
      v0_1173 <= 32'h0;
      v0_1174 <= 32'h0;
      v0_1175 <= 32'h0;
      v0_1176 <= 32'h0;
      v0_1177 <= 32'h0;
      v0_1178 <= 32'h0;
      v0_1179 <= 32'h0;
      v0_1180 <= 32'h0;
      v0_1181 <= 32'h0;
      v0_1182 <= 32'h0;
      v0_1183 <= 32'h0;
      v0_1184 <= 32'h0;
      v0_1185 <= 32'h0;
      v0_1186 <= 32'h0;
      v0_1187 <= 32'h0;
      v0_1188 <= 32'h0;
      v0_1189 <= 32'h0;
      v0_1190 <= 32'h0;
      v0_1191 <= 32'h0;
      v0_1192 <= 32'h0;
      v0_1193 <= 32'h0;
      v0_1194 <= 32'h0;
      v0_1195 <= 32'h0;
      v0_1196 <= 32'h0;
      v0_1197 <= 32'h0;
      v0_1198 <= 32'h0;
      v0_1199 <= 32'h0;
      v0_1200 <= 32'h0;
      v0_1201 <= 32'h0;
      v0_1202 <= 32'h0;
      v0_1203 <= 32'h0;
      v0_1204 <= 32'h0;
      v0_1205 <= 32'h0;
      v0_1206 <= 32'h0;
      v0_1207 <= 32'h0;
      v0_1208 <= 32'h0;
      v0_1209 <= 32'h0;
      v0_1210 <= 32'h0;
      v0_1211 <= 32'h0;
      v0_1212 <= 32'h0;
      v0_1213 <= 32'h0;
      v0_1214 <= 32'h0;
      v0_1215 <= 32'h0;
      v0_1216 <= 32'h0;
      v0_1217 <= 32'h0;
      v0_1218 <= 32'h0;
      v0_1219 <= 32'h0;
      v0_1220 <= 32'h0;
      v0_1221 <= 32'h0;
      v0_1222 <= 32'h0;
      v0_1223 <= 32'h0;
      v0_1224 <= 32'h0;
      v0_1225 <= 32'h0;
      v0_1226 <= 32'h0;
      v0_1227 <= 32'h0;
      v0_1228 <= 32'h0;
      v0_1229 <= 32'h0;
      v0_1230 <= 32'h0;
      v0_1231 <= 32'h0;
      v0_1232 <= 32'h0;
      v0_1233 <= 32'h0;
      v0_1234 <= 32'h0;
      v0_1235 <= 32'h0;
      v0_1236 <= 32'h0;
      v0_1237 <= 32'h0;
      v0_1238 <= 32'h0;
      v0_1239 <= 32'h0;
      v0_1240 <= 32'h0;
      v0_1241 <= 32'h0;
      v0_1242 <= 32'h0;
      v0_1243 <= 32'h0;
      v0_1244 <= 32'h0;
      v0_1245 <= 32'h0;
      v0_1246 <= 32'h0;
      v0_1247 <= 32'h0;
      v0_1248 <= 32'h0;
      v0_1249 <= 32'h0;
      v0_1250 <= 32'h0;
      v0_1251 <= 32'h0;
      v0_1252 <= 32'h0;
      v0_1253 <= 32'h0;
      v0_1254 <= 32'h0;
      v0_1255 <= 32'h0;
      v0_1256 <= 32'h0;
      v0_1257 <= 32'h0;
      v0_1258 <= 32'h0;
      v0_1259 <= 32'h0;
      v0_1260 <= 32'h0;
      v0_1261 <= 32'h0;
      v0_1262 <= 32'h0;
      v0_1263 <= 32'h0;
      v0_1264 <= 32'h0;
      v0_1265 <= 32'h0;
      v0_1266 <= 32'h0;
      v0_1267 <= 32'h0;
      v0_1268 <= 32'h0;
      v0_1269 <= 32'h0;
      v0_1270 <= 32'h0;
      v0_1271 <= 32'h0;
      v0_1272 <= 32'h0;
      v0_1273 <= 32'h0;
      v0_1274 <= 32'h0;
      v0_1275 <= 32'h0;
      v0_1276 <= 32'h0;
      v0_1277 <= 32'h0;
      v0_1278 <= 32'h0;
      v0_1279 <= 32'h0;
      v0_1280 <= 32'h0;
      v0_1281 <= 32'h0;
      v0_1282 <= 32'h0;
      v0_1283 <= 32'h0;
      v0_1284 <= 32'h0;
      v0_1285 <= 32'h0;
      v0_1286 <= 32'h0;
      v0_1287 <= 32'h0;
      v0_1288 <= 32'h0;
      v0_1289 <= 32'h0;
      v0_1290 <= 32'h0;
      v0_1291 <= 32'h0;
      v0_1292 <= 32'h0;
      v0_1293 <= 32'h0;
      v0_1294 <= 32'h0;
      v0_1295 <= 32'h0;
      v0_1296 <= 32'h0;
      v0_1297 <= 32'h0;
      v0_1298 <= 32'h0;
      v0_1299 <= 32'h0;
      v0_1300 <= 32'h0;
      v0_1301 <= 32'h0;
      v0_1302 <= 32'h0;
      v0_1303 <= 32'h0;
      v0_1304 <= 32'h0;
      v0_1305 <= 32'h0;
      v0_1306 <= 32'h0;
      v0_1307 <= 32'h0;
      v0_1308 <= 32'h0;
      v0_1309 <= 32'h0;
      v0_1310 <= 32'h0;
      v0_1311 <= 32'h0;
      v0_1312 <= 32'h0;
      v0_1313 <= 32'h0;
      v0_1314 <= 32'h0;
      v0_1315 <= 32'h0;
      v0_1316 <= 32'h0;
      v0_1317 <= 32'h0;
      v0_1318 <= 32'h0;
      v0_1319 <= 32'h0;
      v0_1320 <= 32'h0;
      v0_1321 <= 32'h0;
      v0_1322 <= 32'h0;
      v0_1323 <= 32'h0;
      v0_1324 <= 32'h0;
      v0_1325 <= 32'h0;
      v0_1326 <= 32'h0;
      v0_1327 <= 32'h0;
      v0_1328 <= 32'h0;
      v0_1329 <= 32'h0;
      v0_1330 <= 32'h0;
      v0_1331 <= 32'h0;
      v0_1332 <= 32'h0;
      v0_1333 <= 32'h0;
      v0_1334 <= 32'h0;
      v0_1335 <= 32'h0;
      v0_1336 <= 32'h0;
      v0_1337 <= 32'h0;
      v0_1338 <= 32'h0;
      v0_1339 <= 32'h0;
      v0_1340 <= 32'h0;
      v0_1341 <= 32'h0;
      v0_1342 <= 32'h0;
      v0_1343 <= 32'h0;
      v0_1344 <= 32'h0;
      v0_1345 <= 32'h0;
      v0_1346 <= 32'h0;
      v0_1347 <= 32'h0;
      v0_1348 <= 32'h0;
      v0_1349 <= 32'h0;
      v0_1350 <= 32'h0;
      v0_1351 <= 32'h0;
      v0_1352 <= 32'h0;
      v0_1353 <= 32'h0;
      v0_1354 <= 32'h0;
      v0_1355 <= 32'h0;
      v0_1356 <= 32'h0;
      v0_1357 <= 32'h0;
      v0_1358 <= 32'h0;
      v0_1359 <= 32'h0;
      v0_1360 <= 32'h0;
      v0_1361 <= 32'h0;
      v0_1362 <= 32'h0;
      v0_1363 <= 32'h0;
      v0_1364 <= 32'h0;
      v0_1365 <= 32'h0;
      v0_1366 <= 32'h0;
      v0_1367 <= 32'h0;
      v0_1368 <= 32'h0;
      v0_1369 <= 32'h0;
      v0_1370 <= 32'h0;
      v0_1371 <= 32'h0;
      v0_1372 <= 32'h0;
      v0_1373 <= 32'h0;
      v0_1374 <= 32'h0;
      v0_1375 <= 32'h0;
      v0_1376 <= 32'h0;
      v0_1377 <= 32'h0;
      v0_1378 <= 32'h0;
      v0_1379 <= 32'h0;
      v0_1380 <= 32'h0;
      v0_1381 <= 32'h0;
      v0_1382 <= 32'h0;
      v0_1383 <= 32'h0;
      v0_1384 <= 32'h0;
      v0_1385 <= 32'h0;
      v0_1386 <= 32'h0;
      v0_1387 <= 32'h0;
      v0_1388 <= 32'h0;
      v0_1389 <= 32'h0;
      v0_1390 <= 32'h0;
      v0_1391 <= 32'h0;
      v0_1392 <= 32'h0;
      v0_1393 <= 32'h0;
      v0_1394 <= 32'h0;
      v0_1395 <= 32'h0;
      v0_1396 <= 32'h0;
      v0_1397 <= 32'h0;
      v0_1398 <= 32'h0;
      v0_1399 <= 32'h0;
      v0_1400 <= 32'h0;
      v0_1401 <= 32'h0;
      v0_1402 <= 32'h0;
      v0_1403 <= 32'h0;
      v0_1404 <= 32'h0;
      v0_1405 <= 32'h0;
      v0_1406 <= 32'h0;
      v0_1407 <= 32'h0;
      v0_1408 <= 32'h0;
      v0_1409 <= 32'h0;
      v0_1410 <= 32'h0;
      v0_1411 <= 32'h0;
      v0_1412 <= 32'h0;
      v0_1413 <= 32'h0;
      v0_1414 <= 32'h0;
      v0_1415 <= 32'h0;
      v0_1416 <= 32'h0;
      v0_1417 <= 32'h0;
      v0_1418 <= 32'h0;
      v0_1419 <= 32'h0;
      v0_1420 <= 32'h0;
      v0_1421 <= 32'h0;
      v0_1422 <= 32'h0;
      v0_1423 <= 32'h0;
      v0_1424 <= 32'h0;
      v0_1425 <= 32'h0;
      v0_1426 <= 32'h0;
      v0_1427 <= 32'h0;
      v0_1428 <= 32'h0;
      v0_1429 <= 32'h0;
      v0_1430 <= 32'h0;
      v0_1431 <= 32'h0;
      v0_1432 <= 32'h0;
      v0_1433 <= 32'h0;
      v0_1434 <= 32'h0;
      v0_1435 <= 32'h0;
      v0_1436 <= 32'h0;
      v0_1437 <= 32'h0;
      v0_1438 <= 32'h0;
      v0_1439 <= 32'h0;
      v0_1440 <= 32'h0;
      v0_1441 <= 32'h0;
      v0_1442 <= 32'h0;
      v0_1443 <= 32'h0;
      v0_1444 <= 32'h0;
      v0_1445 <= 32'h0;
      v0_1446 <= 32'h0;
      v0_1447 <= 32'h0;
      v0_1448 <= 32'h0;
      v0_1449 <= 32'h0;
      v0_1450 <= 32'h0;
      v0_1451 <= 32'h0;
      v0_1452 <= 32'h0;
      v0_1453 <= 32'h0;
      v0_1454 <= 32'h0;
      v0_1455 <= 32'h0;
      v0_1456 <= 32'h0;
      v0_1457 <= 32'h0;
      v0_1458 <= 32'h0;
      v0_1459 <= 32'h0;
      v0_1460 <= 32'h0;
      v0_1461 <= 32'h0;
      v0_1462 <= 32'h0;
      v0_1463 <= 32'h0;
      v0_1464 <= 32'h0;
      v0_1465 <= 32'h0;
      v0_1466 <= 32'h0;
      v0_1467 <= 32'h0;
      v0_1468 <= 32'h0;
      v0_1469 <= 32'h0;
      v0_1470 <= 32'h0;
      v0_1471 <= 32'h0;
      v0_1472 <= 32'h0;
      v0_1473 <= 32'h0;
      v0_1474 <= 32'h0;
      v0_1475 <= 32'h0;
      v0_1476 <= 32'h0;
      v0_1477 <= 32'h0;
      v0_1478 <= 32'h0;
      v0_1479 <= 32'h0;
      v0_1480 <= 32'h0;
      v0_1481 <= 32'h0;
      v0_1482 <= 32'h0;
      v0_1483 <= 32'h0;
      v0_1484 <= 32'h0;
      v0_1485 <= 32'h0;
      v0_1486 <= 32'h0;
      v0_1487 <= 32'h0;
      v0_1488 <= 32'h0;
      v0_1489 <= 32'h0;
      v0_1490 <= 32'h0;
      v0_1491 <= 32'h0;
      v0_1492 <= 32'h0;
      v0_1493 <= 32'h0;
      v0_1494 <= 32'h0;
      v0_1495 <= 32'h0;
      v0_1496 <= 32'h0;
      v0_1497 <= 32'h0;
      v0_1498 <= 32'h0;
      v0_1499 <= 32'h0;
      v0_1500 <= 32'h0;
      v0_1501 <= 32'h0;
      v0_1502 <= 32'h0;
      v0_1503 <= 32'h0;
      v0_1504 <= 32'h0;
      v0_1505 <= 32'h0;
      v0_1506 <= 32'h0;
      v0_1507 <= 32'h0;
      v0_1508 <= 32'h0;
      v0_1509 <= 32'h0;
      v0_1510 <= 32'h0;
      v0_1511 <= 32'h0;
      v0_1512 <= 32'h0;
      v0_1513 <= 32'h0;
      v0_1514 <= 32'h0;
      v0_1515 <= 32'h0;
      v0_1516 <= 32'h0;
      v0_1517 <= 32'h0;
      v0_1518 <= 32'h0;
      v0_1519 <= 32'h0;
      v0_1520 <= 32'h0;
      v0_1521 <= 32'h0;
      v0_1522 <= 32'h0;
      v0_1523 <= 32'h0;
      v0_1524 <= 32'h0;
      v0_1525 <= 32'h0;
      v0_1526 <= 32'h0;
      v0_1527 <= 32'h0;
      v0_1528 <= 32'h0;
      v0_1529 <= 32'h0;
      v0_1530 <= 32'h0;
      v0_1531 <= 32'h0;
      v0_1532 <= 32'h0;
      v0_1533 <= 32'h0;
      v0_1534 <= 32'h0;
      v0_1535 <= 32'h0;
      v0_1536 <= 32'h0;
      v0_1537 <= 32'h0;
      v0_1538 <= 32'h0;
      v0_1539 <= 32'h0;
      v0_1540 <= 32'h0;
      v0_1541 <= 32'h0;
      v0_1542 <= 32'h0;
      v0_1543 <= 32'h0;
      v0_1544 <= 32'h0;
      v0_1545 <= 32'h0;
      v0_1546 <= 32'h0;
      v0_1547 <= 32'h0;
      v0_1548 <= 32'h0;
      v0_1549 <= 32'h0;
      v0_1550 <= 32'h0;
      v0_1551 <= 32'h0;
      v0_1552 <= 32'h0;
      v0_1553 <= 32'h0;
      v0_1554 <= 32'h0;
      v0_1555 <= 32'h0;
      v0_1556 <= 32'h0;
      v0_1557 <= 32'h0;
      v0_1558 <= 32'h0;
      v0_1559 <= 32'h0;
      v0_1560 <= 32'h0;
      v0_1561 <= 32'h0;
      v0_1562 <= 32'h0;
      v0_1563 <= 32'h0;
      v0_1564 <= 32'h0;
      v0_1565 <= 32'h0;
      v0_1566 <= 32'h0;
      v0_1567 <= 32'h0;
      v0_1568 <= 32'h0;
      v0_1569 <= 32'h0;
      v0_1570 <= 32'h0;
      v0_1571 <= 32'h0;
      v0_1572 <= 32'h0;
      v0_1573 <= 32'h0;
      v0_1574 <= 32'h0;
      v0_1575 <= 32'h0;
      v0_1576 <= 32'h0;
      v0_1577 <= 32'h0;
      v0_1578 <= 32'h0;
      v0_1579 <= 32'h0;
      v0_1580 <= 32'h0;
      v0_1581 <= 32'h0;
      v0_1582 <= 32'h0;
      v0_1583 <= 32'h0;
      v0_1584 <= 32'h0;
      v0_1585 <= 32'h0;
      v0_1586 <= 32'h0;
      v0_1587 <= 32'h0;
      v0_1588 <= 32'h0;
      v0_1589 <= 32'h0;
      v0_1590 <= 32'h0;
      v0_1591 <= 32'h0;
      v0_1592 <= 32'h0;
      v0_1593 <= 32'h0;
      v0_1594 <= 32'h0;
      v0_1595 <= 32'h0;
      v0_1596 <= 32'h0;
      v0_1597 <= 32'h0;
      v0_1598 <= 32'h0;
      v0_1599 <= 32'h0;
      v0_1600 <= 32'h0;
      v0_1601 <= 32'h0;
      v0_1602 <= 32'h0;
      v0_1603 <= 32'h0;
      v0_1604 <= 32'h0;
      v0_1605 <= 32'h0;
      v0_1606 <= 32'h0;
      v0_1607 <= 32'h0;
      v0_1608 <= 32'h0;
      v0_1609 <= 32'h0;
      v0_1610 <= 32'h0;
      v0_1611 <= 32'h0;
      v0_1612 <= 32'h0;
      v0_1613 <= 32'h0;
      v0_1614 <= 32'h0;
      v0_1615 <= 32'h0;
      v0_1616 <= 32'h0;
      v0_1617 <= 32'h0;
      v0_1618 <= 32'h0;
      v0_1619 <= 32'h0;
      v0_1620 <= 32'h0;
      v0_1621 <= 32'h0;
      v0_1622 <= 32'h0;
      v0_1623 <= 32'h0;
      v0_1624 <= 32'h0;
      v0_1625 <= 32'h0;
      v0_1626 <= 32'h0;
      v0_1627 <= 32'h0;
      v0_1628 <= 32'h0;
      v0_1629 <= 32'h0;
      v0_1630 <= 32'h0;
      v0_1631 <= 32'h0;
      v0_1632 <= 32'h0;
      v0_1633 <= 32'h0;
      v0_1634 <= 32'h0;
      v0_1635 <= 32'h0;
      v0_1636 <= 32'h0;
      v0_1637 <= 32'h0;
      v0_1638 <= 32'h0;
      v0_1639 <= 32'h0;
      v0_1640 <= 32'h0;
      v0_1641 <= 32'h0;
      v0_1642 <= 32'h0;
      v0_1643 <= 32'h0;
      v0_1644 <= 32'h0;
      v0_1645 <= 32'h0;
      v0_1646 <= 32'h0;
      v0_1647 <= 32'h0;
      v0_1648 <= 32'h0;
      v0_1649 <= 32'h0;
      v0_1650 <= 32'h0;
      v0_1651 <= 32'h0;
      v0_1652 <= 32'h0;
      v0_1653 <= 32'h0;
      v0_1654 <= 32'h0;
      v0_1655 <= 32'h0;
      v0_1656 <= 32'h0;
      v0_1657 <= 32'h0;
      v0_1658 <= 32'h0;
      v0_1659 <= 32'h0;
      v0_1660 <= 32'h0;
      v0_1661 <= 32'h0;
      v0_1662 <= 32'h0;
      v0_1663 <= 32'h0;
      v0_1664 <= 32'h0;
      v0_1665 <= 32'h0;
      v0_1666 <= 32'h0;
      v0_1667 <= 32'h0;
      v0_1668 <= 32'h0;
      v0_1669 <= 32'h0;
      v0_1670 <= 32'h0;
      v0_1671 <= 32'h0;
      v0_1672 <= 32'h0;
      v0_1673 <= 32'h0;
      v0_1674 <= 32'h0;
      v0_1675 <= 32'h0;
      v0_1676 <= 32'h0;
      v0_1677 <= 32'h0;
      v0_1678 <= 32'h0;
      v0_1679 <= 32'h0;
      v0_1680 <= 32'h0;
      v0_1681 <= 32'h0;
      v0_1682 <= 32'h0;
      v0_1683 <= 32'h0;
      v0_1684 <= 32'h0;
      v0_1685 <= 32'h0;
      v0_1686 <= 32'h0;
      v0_1687 <= 32'h0;
      v0_1688 <= 32'h0;
      v0_1689 <= 32'h0;
      v0_1690 <= 32'h0;
      v0_1691 <= 32'h0;
      v0_1692 <= 32'h0;
      v0_1693 <= 32'h0;
      v0_1694 <= 32'h0;
      v0_1695 <= 32'h0;
      v0_1696 <= 32'h0;
      v0_1697 <= 32'h0;
      v0_1698 <= 32'h0;
      v0_1699 <= 32'h0;
      v0_1700 <= 32'h0;
      v0_1701 <= 32'h0;
      v0_1702 <= 32'h0;
      v0_1703 <= 32'h0;
      v0_1704 <= 32'h0;
      v0_1705 <= 32'h0;
      v0_1706 <= 32'h0;
      v0_1707 <= 32'h0;
      v0_1708 <= 32'h0;
      v0_1709 <= 32'h0;
      v0_1710 <= 32'h0;
      v0_1711 <= 32'h0;
      v0_1712 <= 32'h0;
      v0_1713 <= 32'h0;
      v0_1714 <= 32'h0;
      v0_1715 <= 32'h0;
      v0_1716 <= 32'h0;
      v0_1717 <= 32'h0;
      v0_1718 <= 32'h0;
      v0_1719 <= 32'h0;
      v0_1720 <= 32'h0;
      v0_1721 <= 32'h0;
      v0_1722 <= 32'h0;
      v0_1723 <= 32'h0;
      v0_1724 <= 32'h0;
      v0_1725 <= 32'h0;
      v0_1726 <= 32'h0;
      v0_1727 <= 32'h0;
      v0_1728 <= 32'h0;
      v0_1729 <= 32'h0;
      v0_1730 <= 32'h0;
      v0_1731 <= 32'h0;
      v0_1732 <= 32'h0;
      v0_1733 <= 32'h0;
      v0_1734 <= 32'h0;
      v0_1735 <= 32'h0;
      v0_1736 <= 32'h0;
      v0_1737 <= 32'h0;
      v0_1738 <= 32'h0;
      v0_1739 <= 32'h0;
      v0_1740 <= 32'h0;
      v0_1741 <= 32'h0;
      v0_1742 <= 32'h0;
      v0_1743 <= 32'h0;
      v0_1744 <= 32'h0;
      v0_1745 <= 32'h0;
      v0_1746 <= 32'h0;
      v0_1747 <= 32'h0;
      v0_1748 <= 32'h0;
      v0_1749 <= 32'h0;
      v0_1750 <= 32'h0;
      v0_1751 <= 32'h0;
      v0_1752 <= 32'h0;
      v0_1753 <= 32'h0;
      v0_1754 <= 32'h0;
      v0_1755 <= 32'h0;
      v0_1756 <= 32'h0;
      v0_1757 <= 32'h0;
      v0_1758 <= 32'h0;
      v0_1759 <= 32'h0;
      v0_1760 <= 32'h0;
      v0_1761 <= 32'h0;
      v0_1762 <= 32'h0;
      v0_1763 <= 32'h0;
      v0_1764 <= 32'h0;
      v0_1765 <= 32'h0;
      v0_1766 <= 32'h0;
      v0_1767 <= 32'h0;
      v0_1768 <= 32'h0;
      v0_1769 <= 32'h0;
      v0_1770 <= 32'h0;
      v0_1771 <= 32'h0;
      v0_1772 <= 32'h0;
      v0_1773 <= 32'h0;
      v0_1774 <= 32'h0;
      v0_1775 <= 32'h0;
      v0_1776 <= 32'h0;
      v0_1777 <= 32'h0;
      v0_1778 <= 32'h0;
      v0_1779 <= 32'h0;
      v0_1780 <= 32'h0;
      v0_1781 <= 32'h0;
      v0_1782 <= 32'h0;
      v0_1783 <= 32'h0;
      v0_1784 <= 32'h0;
      v0_1785 <= 32'h0;
      v0_1786 <= 32'h0;
      v0_1787 <= 32'h0;
      v0_1788 <= 32'h0;
      v0_1789 <= 32'h0;
      v0_1790 <= 32'h0;
      v0_1791 <= 32'h0;
      v0_1792 <= 32'h0;
      v0_1793 <= 32'h0;
      v0_1794 <= 32'h0;
      v0_1795 <= 32'h0;
      v0_1796 <= 32'h0;
      v0_1797 <= 32'h0;
      v0_1798 <= 32'h0;
      v0_1799 <= 32'h0;
      v0_1800 <= 32'h0;
      v0_1801 <= 32'h0;
      v0_1802 <= 32'h0;
      v0_1803 <= 32'h0;
      v0_1804 <= 32'h0;
      v0_1805 <= 32'h0;
      v0_1806 <= 32'h0;
      v0_1807 <= 32'h0;
      v0_1808 <= 32'h0;
      v0_1809 <= 32'h0;
      v0_1810 <= 32'h0;
      v0_1811 <= 32'h0;
      v0_1812 <= 32'h0;
      v0_1813 <= 32'h0;
      v0_1814 <= 32'h0;
      v0_1815 <= 32'h0;
      v0_1816 <= 32'h0;
      v0_1817 <= 32'h0;
      v0_1818 <= 32'h0;
      v0_1819 <= 32'h0;
      v0_1820 <= 32'h0;
      v0_1821 <= 32'h0;
      v0_1822 <= 32'h0;
      v0_1823 <= 32'h0;
      v0_1824 <= 32'h0;
      v0_1825 <= 32'h0;
      v0_1826 <= 32'h0;
      v0_1827 <= 32'h0;
      v0_1828 <= 32'h0;
      v0_1829 <= 32'h0;
      v0_1830 <= 32'h0;
      v0_1831 <= 32'h0;
      v0_1832 <= 32'h0;
      v0_1833 <= 32'h0;
      v0_1834 <= 32'h0;
      v0_1835 <= 32'h0;
      v0_1836 <= 32'h0;
      v0_1837 <= 32'h0;
      v0_1838 <= 32'h0;
      v0_1839 <= 32'h0;
      v0_1840 <= 32'h0;
      v0_1841 <= 32'h0;
      v0_1842 <= 32'h0;
      v0_1843 <= 32'h0;
      v0_1844 <= 32'h0;
      v0_1845 <= 32'h0;
      v0_1846 <= 32'h0;
      v0_1847 <= 32'h0;
      v0_1848 <= 32'h0;
      v0_1849 <= 32'h0;
      v0_1850 <= 32'h0;
      v0_1851 <= 32'h0;
      v0_1852 <= 32'h0;
      v0_1853 <= 32'h0;
      v0_1854 <= 32'h0;
      v0_1855 <= 32'h0;
      v0_1856 <= 32'h0;
      v0_1857 <= 32'h0;
      v0_1858 <= 32'h0;
      v0_1859 <= 32'h0;
      v0_1860 <= 32'h0;
      v0_1861 <= 32'h0;
      v0_1862 <= 32'h0;
      v0_1863 <= 32'h0;
      v0_1864 <= 32'h0;
      v0_1865 <= 32'h0;
      v0_1866 <= 32'h0;
      v0_1867 <= 32'h0;
      v0_1868 <= 32'h0;
      v0_1869 <= 32'h0;
      v0_1870 <= 32'h0;
      v0_1871 <= 32'h0;
      v0_1872 <= 32'h0;
      v0_1873 <= 32'h0;
      v0_1874 <= 32'h0;
      v0_1875 <= 32'h0;
      v0_1876 <= 32'h0;
      v0_1877 <= 32'h0;
      v0_1878 <= 32'h0;
      v0_1879 <= 32'h0;
      v0_1880 <= 32'h0;
      v0_1881 <= 32'h0;
      v0_1882 <= 32'h0;
      v0_1883 <= 32'h0;
      v0_1884 <= 32'h0;
      v0_1885 <= 32'h0;
      v0_1886 <= 32'h0;
      v0_1887 <= 32'h0;
      v0_1888 <= 32'h0;
      v0_1889 <= 32'h0;
      v0_1890 <= 32'h0;
      v0_1891 <= 32'h0;
      v0_1892 <= 32'h0;
      v0_1893 <= 32'h0;
      v0_1894 <= 32'h0;
      v0_1895 <= 32'h0;
      v0_1896 <= 32'h0;
      v0_1897 <= 32'h0;
      v0_1898 <= 32'h0;
      v0_1899 <= 32'h0;
      v0_1900 <= 32'h0;
      v0_1901 <= 32'h0;
      v0_1902 <= 32'h0;
      v0_1903 <= 32'h0;
      v0_1904 <= 32'h0;
      v0_1905 <= 32'h0;
      v0_1906 <= 32'h0;
      v0_1907 <= 32'h0;
      v0_1908 <= 32'h0;
      v0_1909 <= 32'h0;
      v0_1910 <= 32'h0;
      v0_1911 <= 32'h0;
      v0_1912 <= 32'h0;
      v0_1913 <= 32'h0;
      v0_1914 <= 32'h0;
      v0_1915 <= 32'h0;
      v0_1916 <= 32'h0;
      v0_1917 <= 32'h0;
      v0_1918 <= 32'h0;
      v0_1919 <= 32'h0;
      v0_1920 <= 32'h0;
      v0_1921 <= 32'h0;
      v0_1922 <= 32'h0;
      v0_1923 <= 32'h0;
      v0_1924 <= 32'h0;
      v0_1925 <= 32'h0;
      v0_1926 <= 32'h0;
      v0_1927 <= 32'h0;
      v0_1928 <= 32'h0;
      v0_1929 <= 32'h0;
      v0_1930 <= 32'h0;
      v0_1931 <= 32'h0;
      v0_1932 <= 32'h0;
      v0_1933 <= 32'h0;
      v0_1934 <= 32'h0;
      v0_1935 <= 32'h0;
      v0_1936 <= 32'h0;
      v0_1937 <= 32'h0;
      v0_1938 <= 32'h0;
      v0_1939 <= 32'h0;
      v0_1940 <= 32'h0;
      v0_1941 <= 32'h0;
      v0_1942 <= 32'h0;
      v0_1943 <= 32'h0;
      v0_1944 <= 32'h0;
      v0_1945 <= 32'h0;
      v0_1946 <= 32'h0;
      v0_1947 <= 32'h0;
      v0_1948 <= 32'h0;
      v0_1949 <= 32'h0;
      v0_1950 <= 32'h0;
      v0_1951 <= 32'h0;
      v0_1952 <= 32'h0;
      v0_1953 <= 32'h0;
      v0_1954 <= 32'h0;
      v0_1955 <= 32'h0;
      v0_1956 <= 32'h0;
      v0_1957 <= 32'h0;
      v0_1958 <= 32'h0;
      v0_1959 <= 32'h0;
      v0_1960 <= 32'h0;
      v0_1961 <= 32'h0;
      v0_1962 <= 32'h0;
      v0_1963 <= 32'h0;
      v0_1964 <= 32'h0;
      v0_1965 <= 32'h0;
      v0_1966 <= 32'h0;
      v0_1967 <= 32'h0;
      v0_1968 <= 32'h0;
      v0_1969 <= 32'h0;
      v0_1970 <= 32'h0;
      v0_1971 <= 32'h0;
      v0_1972 <= 32'h0;
      v0_1973 <= 32'h0;
      v0_1974 <= 32'h0;
      v0_1975 <= 32'h0;
      v0_1976 <= 32'h0;
      v0_1977 <= 32'h0;
      v0_1978 <= 32'h0;
      v0_1979 <= 32'h0;
      v0_1980 <= 32'h0;
      v0_1981 <= 32'h0;
      v0_1982 <= 32'h0;
      v0_1983 <= 32'h0;
      v0_1984 <= 32'h0;
      v0_1985 <= 32'h0;
      v0_1986 <= 32'h0;
      v0_1987 <= 32'h0;
      v0_1988 <= 32'h0;
      v0_1989 <= 32'h0;
      v0_1990 <= 32'h0;
      v0_1991 <= 32'h0;
      v0_1992 <= 32'h0;
      v0_1993 <= 32'h0;
      v0_1994 <= 32'h0;
      v0_1995 <= 32'h0;
      v0_1996 <= 32'h0;
      v0_1997 <= 32'h0;
      v0_1998 <= 32'h0;
      v0_1999 <= 32'h0;
      v0_2000 <= 32'h0;
      v0_2001 <= 32'h0;
      v0_2002 <= 32'h0;
      v0_2003 <= 32'h0;
      v0_2004 <= 32'h0;
      v0_2005 <= 32'h0;
      v0_2006 <= 32'h0;
      v0_2007 <= 32'h0;
      v0_2008 <= 32'h0;
      v0_2009 <= 32'h0;
      v0_2010 <= 32'h0;
      v0_2011 <= 32'h0;
      v0_2012 <= 32'h0;
      v0_2013 <= 32'h0;
      v0_2014 <= 32'h0;
      v0_2015 <= 32'h0;
      v0_2016 <= 32'h0;
      v0_2017 <= 32'h0;
      v0_2018 <= 32'h0;
      v0_2019 <= 32'h0;
      v0_2020 <= 32'h0;
      v0_2021 <= 32'h0;
      v0_2022 <= 32'h0;
      v0_2023 <= 32'h0;
      v0_2024 <= 32'h0;
      v0_2025 <= 32'h0;
      v0_2026 <= 32'h0;
      v0_2027 <= 32'h0;
      v0_2028 <= 32'h0;
      v0_2029 <= 32'h0;
      v0_2030 <= 32'h0;
      v0_2031 <= 32'h0;
      v0_2032 <= 32'h0;
      v0_2033 <= 32'h0;
      v0_2034 <= 32'h0;
      v0_2035 <= 32'h0;
      v0_2036 <= 32'h0;
      v0_2037 <= 32'h0;
      v0_2038 <= 32'h0;
      v0_2039 <= 32'h0;
      v0_2040 <= 32'h0;
      v0_2041 <= 32'h0;
      v0_2042 <= 32'h0;
      v0_2043 <= 32'h0;
      v0_2044 <= 32'h0;
      v0_2045 <= 32'h0;
      v0_2046 <= 32'h0;
      v0_2047 <= 32'h0;
      queueCount_0 <= 7'h0;
      queueCount_1 <= 7'h0;
      queueCount_2 <= 7'h0;
      queueCount_3 <= 7'h0;
      queueCount_4 <= 7'h0;
      queueCount_5 <= 7'h0;
      queueCount_6 <= 7'h0;
      queueCount_7 <= 7'h0;
      queueCount_0_1 <= 7'h0;
      queueCount_1_1 <= 7'h0;
      queueCount_2_1 <= 7'h0;
      queueCount_3_1 <= 7'h0;
      queueCount_4_1 <= 7'h0;
      queueCount_5_1 <= 7'h0;
      queueCount_6_1 <= 7'h0;
      queueCount_7_1 <= 7'h0;
      queueCount_0_2 <= 7'h0;
      queueCount_1_2 <= 7'h0;
      queueCount_2_2 <= 7'h0;
      queueCount_3_2 <= 7'h0;
      queueCount_4_2 <= 7'h0;
      queueCount_5_2 <= 7'h0;
      queueCount_6_2 <= 7'h0;
      queueCount_7_2 <= 7'h0;
      queueCount_0_3 <= 7'h0;
      queueCount_1_3 <= 7'h0;
      queueCount_2_3 <= 7'h0;
      queueCount_3_3 <= 7'h0;
      queueCount_4_3 <= 7'h0;
      queueCount_5_3 <= 7'h0;
      queueCount_6_3 <= 7'h0;
      queueCount_7_3 <= 7'h0;
    end
    else begin
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h0)
        v0_0 <= v0_0 & ~maskExt | maskExt & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h0)
        v0_1 <= v0_1 & ~maskExt_1 | maskExt_1 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h0)
        v0_2 <= v0_2 & ~maskExt_2 | maskExt_2 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h0)
        v0_3 <= v0_3 & ~maskExt_3 | maskExt_3 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1)
        v0_4 <= v0_4 & ~maskExt_4 | maskExt_4 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1)
        v0_5 <= v0_5 & ~maskExt_5 | maskExt_5 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1)
        v0_6 <= v0_6 & ~maskExt_6 | maskExt_6 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1)
        v0_7 <= v0_7 & ~maskExt_7 | maskExt_7 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h2)
        v0_8 <= v0_8 & ~maskExt_8 | maskExt_8 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h2)
        v0_9 <= v0_9 & ~maskExt_9 | maskExt_9 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h2)
        v0_10 <= v0_10 & ~maskExt_10 | maskExt_10 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h2)
        v0_11 <= v0_11 & ~maskExt_11 | maskExt_11 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h3)
        v0_12 <= v0_12 & ~maskExt_12 | maskExt_12 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h3)
        v0_13 <= v0_13 & ~maskExt_13 | maskExt_13 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h3)
        v0_14 <= v0_14 & ~maskExt_14 | maskExt_14 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h3)
        v0_15 <= v0_15 & ~maskExt_15 | maskExt_15 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h4)
        v0_16 <= v0_16 & ~maskExt_16 | maskExt_16 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h4)
        v0_17 <= v0_17 & ~maskExt_17 | maskExt_17 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h4)
        v0_18 <= v0_18 & ~maskExt_18 | maskExt_18 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h4)
        v0_19 <= v0_19 & ~maskExt_19 | maskExt_19 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h5)
        v0_20 <= v0_20 & ~maskExt_20 | maskExt_20 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h5)
        v0_21 <= v0_21 & ~maskExt_21 | maskExt_21 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h5)
        v0_22 <= v0_22 & ~maskExt_22 | maskExt_22 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h5)
        v0_23 <= v0_23 & ~maskExt_23 | maskExt_23 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h6)
        v0_24 <= v0_24 & ~maskExt_24 | maskExt_24 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h6)
        v0_25 <= v0_25 & ~maskExt_25 | maskExt_25 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h6)
        v0_26 <= v0_26 & ~maskExt_26 | maskExt_26 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h6)
        v0_27 <= v0_27 & ~maskExt_27 | maskExt_27 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h7)
        v0_28 <= v0_28 & ~maskExt_28 | maskExt_28 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h7)
        v0_29 <= v0_29 & ~maskExt_29 | maskExt_29 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h7)
        v0_30 <= v0_30 & ~maskExt_30 | maskExt_30 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h7)
        v0_31 <= v0_31 & ~maskExt_31 | maskExt_31 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h8)
        v0_32 <= v0_32 & ~maskExt_32 | maskExt_32 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h8)
        v0_33 <= v0_33 & ~maskExt_33 | maskExt_33 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h8)
        v0_34 <= v0_34 & ~maskExt_34 | maskExt_34 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h8)
        v0_35 <= v0_35 & ~maskExt_35 | maskExt_35 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h9)
        v0_36 <= v0_36 & ~maskExt_36 | maskExt_36 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h9)
        v0_37 <= v0_37 & ~maskExt_37 | maskExt_37 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h9)
        v0_38 <= v0_38 & ~maskExt_38 | maskExt_38 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h9)
        v0_39 <= v0_39 & ~maskExt_39 | maskExt_39 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hA)
        v0_40 <= v0_40 & ~maskExt_40 | maskExt_40 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hA)
        v0_41 <= v0_41 & ~maskExt_41 | maskExt_41 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hA)
        v0_42 <= v0_42 & ~maskExt_42 | maskExt_42 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hA)
        v0_43 <= v0_43 & ~maskExt_43 | maskExt_43 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hB)
        v0_44 <= v0_44 & ~maskExt_44 | maskExt_44 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hB)
        v0_45 <= v0_45 & ~maskExt_45 | maskExt_45 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hB)
        v0_46 <= v0_46 & ~maskExt_46 | maskExt_46 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hB)
        v0_47 <= v0_47 & ~maskExt_47 | maskExt_47 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hC)
        v0_48 <= v0_48 & ~maskExt_48 | maskExt_48 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hC)
        v0_49 <= v0_49 & ~maskExt_49 | maskExt_49 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hC)
        v0_50 <= v0_50 & ~maskExt_50 | maskExt_50 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hC)
        v0_51 <= v0_51 & ~maskExt_51 | maskExt_51 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hD)
        v0_52 <= v0_52 & ~maskExt_52 | maskExt_52 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hD)
        v0_53 <= v0_53 & ~maskExt_53 | maskExt_53 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hD)
        v0_54 <= v0_54 & ~maskExt_54 | maskExt_54 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hD)
        v0_55 <= v0_55 & ~maskExt_55 | maskExt_55 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hE)
        v0_56 <= v0_56 & ~maskExt_56 | maskExt_56 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hE)
        v0_57 <= v0_57 & ~maskExt_57 | maskExt_57 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hE)
        v0_58 <= v0_58 & ~maskExt_58 | maskExt_58 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hE)
        v0_59 <= v0_59 & ~maskExt_59 | maskExt_59 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hF)
        v0_60 <= v0_60 & ~maskExt_60 | maskExt_60 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hF)
        v0_61 <= v0_61 & ~maskExt_61 | maskExt_61 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hF)
        v0_62 <= v0_62 & ~maskExt_62 | maskExt_62 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hF)
        v0_63 <= v0_63 & ~maskExt_63 | maskExt_63 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h10)
        v0_64 <= v0_64 & ~maskExt_64 | maskExt_64 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h10)
        v0_65 <= v0_65 & ~maskExt_65 | maskExt_65 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h10)
        v0_66 <= v0_66 & ~maskExt_66 | maskExt_66 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h10)
        v0_67 <= v0_67 & ~maskExt_67 | maskExt_67 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h11)
        v0_68 <= v0_68 & ~maskExt_68 | maskExt_68 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h11)
        v0_69 <= v0_69 & ~maskExt_69 | maskExt_69 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h11)
        v0_70 <= v0_70 & ~maskExt_70 | maskExt_70 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h11)
        v0_71 <= v0_71 & ~maskExt_71 | maskExt_71 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h12)
        v0_72 <= v0_72 & ~maskExt_72 | maskExt_72 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h12)
        v0_73 <= v0_73 & ~maskExt_73 | maskExt_73 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h12)
        v0_74 <= v0_74 & ~maskExt_74 | maskExt_74 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h12)
        v0_75 <= v0_75 & ~maskExt_75 | maskExt_75 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h13)
        v0_76 <= v0_76 & ~maskExt_76 | maskExt_76 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h13)
        v0_77 <= v0_77 & ~maskExt_77 | maskExt_77 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h13)
        v0_78 <= v0_78 & ~maskExt_78 | maskExt_78 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h13)
        v0_79 <= v0_79 & ~maskExt_79 | maskExt_79 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h14)
        v0_80 <= v0_80 & ~maskExt_80 | maskExt_80 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h14)
        v0_81 <= v0_81 & ~maskExt_81 | maskExt_81 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h14)
        v0_82 <= v0_82 & ~maskExt_82 | maskExt_82 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h14)
        v0_83 <= v0_83 & ~maskExt_83 | maskExt_83 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h15)
        v0_84 <= v0_84 & ~maskExt_84 | maskExt_84 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h15)
        v0_85 <= v0_85 & ~maskExt_85 | maskExt_85 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h15)
        v0_86 <= v0_86 & ~maskExt_86 | maskExt_86 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h15)
        v0_87 <= v0_87 & ~maskExt_87 | maskExt_87 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h16)
        v0_88 <= v0_88 & ~maskExt_88 | maskExt_88 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h16)
        v0_89 <= v0_89 & ~maskExt_89 | maskExt_89 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h16)
        v0_90 <= v0_90 & ~maskExt_90 | maskExt_90 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h16)
        v0_91 <= v0_91 & ~maskExt_91 | maskExt_91 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h17)
        v0_92 <= v0_92 & ~maskExt_92 | maskExt_92 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h17)
        v0_93 <= v0_93 & ~maskExt_93 | maskExt_93 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h17)
        v0_94 <= v0_94 & ~maskExt_94 | maskExt_94 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h17)
        v0_95 <= v0_95 & ~maskExt_95 | maskExt_95 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h18)
        v0_96 <= v0_96 & ~maskExt_96 | maskExt_96 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h18)
        v0_97 <= v0_97 & ~maskExt_97 | maskExt_97 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h18)
        v0_98 <= v0_98 & ~maskExt_98 | maskExt_98 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h18)
        v0_99 <= v0_99 & ~maskExt_99 | maskExt_99 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h19)
        v0_100 <= v0_100 & ~maskExt_100 | maskExt_100 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h19)
        v0_101 <= v0_101 & ~maskExt_101 | maskExt_101 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h19)
        v0_102 <= v0_102 & ~maskExt_102 | maskExt_102 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h19)
        v0_103 <= v0_103 & ~maskExt_103 | maskExt_103 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1A)
        v0_104 <= v0_104 & ~maskExt_104 | maskExt_104 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1A)
        v0_105 <= v0_105 & ~maskExt_105 | maskExt_105 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1A)
        v0_106 <= v0_106 & ~maskExt_106 | maskExt_106 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1A)
        v0_107 <= v0_107 & ~maskExt_107 | maskExt_107 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1B)
        v0_108 <= v0_108 & ~maskExt_108 | maskExt_108 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1B)
        v0_109 <= v0_109 & ~maskExt_109 | maskExt_109 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1B)
        v0_110 <= v0_110 & ~maskExt_110 | maskExt_110 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1B)
        v0_111 <= v0_111 & ~maskExt_111 | maskExt_111 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1C)
        v0_112 <= v0_112 & ~maskExt_112 | maskExt_112 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1C)
        v0_113 <= v0_113 & ~maskExt_113 | maskExt_113 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1C)
        v0_114 <= v0_114 & ~maskExt_114 | maskExt_114 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1C)
        v0_115 <= v0_115 & ~maskExt_115 | maskExt_115 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1D)
        v0_116 <= v0_116 & ~maskExt_116 | maskExt_116 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1D)
        v0_117 <= v0_117 & ~maskExt_117 | maskExt_117 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1D)
        v0_118 <= v0_118 & ~maskExt_118 | maskExt_118 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1D)
        v0_119 <= v0_119 & ~maskExt_119 | maskExt_119 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1E)
        v0_120 <= v0_120 & ~maskExt_120 | maskExt_120 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1E)
        v0_121 <= v0_121 & ~maskExt_121 | maskExt_121 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1E)
        v0_122 <= v0_122 & ~maskExt_122 | maskExt_122 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1E)
        v0_123 <= v0_123 & ~maskExt_123 | maskExt_123 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1F)
        v0_124 <= v0_124 & ~maskExt_124 | maskExt_124 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1F)
        v0_125 <= v0_125 & ~maskExt_125 | maskExt_125 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1F)
        v0_126 <= v0_126 & ~maskExt_126 | maskExt_126 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1F)
        v0_127 <= v0_127 & ~maskExt_127 | maskExt_127 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h20)
        v0_128 <= v0_128 & ~maskExt_128 | maskExt_128 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h20)
        v0_129 <= v0_129 & ~maskExt_129 | maskExt_129 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h20)
        v0_130 <= v0_130 & ~maskExt_130 | maskExt_130 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h20)
        v0_131 <= v0_131 & ~maskExt_131 | maskExt_131 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h21)
        v0_132 <= v0_132 & ~maskExt_132 | maskExt_132 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h21)
        v0_133 <= v0_133 & ~maskExt_133 | maskExt_133 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h21)
        v0_134 <= v0_134 & ~maskExt_134 | maskExt_134 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h21)
        v0_135 <= v0_135 & ~maskExt_135 | maskExt_135 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h22)
        v0_136 <= v0_136 & ~maskExt_136 | maskExt_136 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h22)
        v0_137 <= v0_137 & ~maskExt_137 | maskExt_137 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h22)
        v0_138 <= v0_138 & ~maskExt_138 | maskExt_138 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h22)
        v0_139 <= v0_139 & ~maskExt_139 | maskExt_139 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h23)
        v0_140 <= v0_140 & ~maskExt_140 | maskExt_140 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h23)
        v0_141 <= v0_141 & ~maskExt_141 | maskExt_141 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h23)
        v0_142 <= v0_142 & ~maskExt_142 | maskExt_142 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h23)
        v0_143 <= v0_143 & ~maskExt_143 | maskExt_143 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h24)
        v0_144 <= v0_144 & ~maskExt_144 | maskExt_144 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h24)
        v0_145 <= v0_145 & ~maskExt_145 | maskExt_145 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h24)
        v0_146 <= v0_146 & ~maskExt_146 | maskExt_146 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h24)
        v0_147 <= v0_147 & ~maskExt_147 | maskExt_147 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h25)
        v0_148 <= v0_148 & ~maskExt_148 | maskExt_148 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h25)
        v0_149 <= v0_149 & ~maskExt_149 | maskExt_149 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h25)
        v0_150 <= v0_150 & ~maskExt_150 | maskExt_150 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h25)
        v0_151 <= v0_151 & ~maskExt_151 | maskExt_151 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h26)
        v0_152 <= v0_152 & ~maskExt_152 | maskExt_152 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h26)
        v0_153 <= v0_153 & ~maskExt_153 | maskExt_153 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h26)
        v0_154 <= v0_154 & ~maskExt_154 | maskExt_154 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h26)
        v0_155 <= v0_155 & ~maskExt_155 | maskExt_155 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h27)
        v0_156 <= v0_156 & ~maskExt_156 | maskExt_156 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h27)
        v0_157 <= v0_157 & ~maskExt_157 | maskExt_157 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h27)
        v0_158 <= v0_158 & ~maskExt_158 | maskExt_158 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h27)
        v0_159 <= v0_159 & ~maskExt_159 | maskExt_159 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h28)
        v0_160 <= v0_160 & ~maskExt_160 | maskExt_160 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h28)
        v0_161 <= v0_161 & ~maskExt_161 | maskExt_161 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h28)
        v0_162 <= v0_162 & ~maskExt_162 | maskExt_162 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h28)
        v0_163 <= v0_163 & ~maskExt_163 | maskExt_163 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h29)
        v0_164 <= v0_164 & ~maskExt_164 | maskExt_164 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h29)
        v0_165 <= v0_165 & ~maskExt_165 | maskExt_165 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h29)
        v0_166 <= v0_166 & ~maskExt_166 | maskExt_166 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h29)
        v0_167 <= v0_167 & ~maskExt_167 | maskExt_167 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h2A)
        v0_168 <= v0_168 & ~maskExt_168 | maskExt_168 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h2A)
        v0_169 <= v0_169 & ~maskExt_169 | maskExt_169 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h2A)
        v0_170 <= v0_170 & ~maskExt_170 | maskExt_170 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h2A)
        v0_171 <= v0_171 & ~maskExt_171 | maskExt_171 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h2B)
        v0_172 <= v0_172 & ~maskExt_172 | maskExt_172 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h2B)
        v0_173 <= v0_173 & ~maskExt_173 | maskExt_173 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h2B)
        v0_174 <= v0_174 & ~maskExt_174 | maskExt_174 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h2B)
        v0_175 <= v0_175 & ~maskExt_175 | maskExt_175 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h2C)
        v0_176 <= v0_176 & ~maskExt_176 | maskExt_176 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h2C)
        v0_177 <= v0_177 & ~maskExt_177 | maskExt_177 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h2C)
        v0_178 <= v0_178 & ~maskExt_178 | maskExt_178 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h2C)
        v0_179 <= v0_179 & ~maskExt_179 | maskExt_179 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h2D)
        v0_180 <= v0_180 & ~maskExt_180 | maskExt_180 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h2D)
        v0_181 <= v0_181 & ~maskExt_181 | maskExt_181 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h2D)
        v0_182 <= v0_182 & ~maskExt_182 | maskExt_182 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h2D)
        v0_183 <= v0_183 & ~maskExt_183 | maskExt_183 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h2E)
        v0_184 <= v0_184 & ~maskExt_184 | maskExt_184 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h2E)
        v0_185 <= v0_185 & ~maskExt_185 | maskExt_185 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h2E)
        v0_186 <= v0_186 & ~maskExt_186 | maskExt_186 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h2E)
        v0_187 <= v0_187 & ~maskExt_187 | maskExt_187 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h2F)
        v0_188 <= v0_188 & ~maskExt_188 | maskExt_188 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h2F)
        v0_189 <= v0_189 & ~maskExt_189 | maskExt_189 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h2F)
        v0_190 <= v0_190 & ~maskExt_190 | maskExt_190 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h2F)
        v0_191 <= v0_191 & ~maskExt_191 | maskExt_191 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h30)
        v0_192 <= v0_192 & ~maskExt_192 | maskExt_192 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h30)
        v0_193 <= v0_193 & ~maskExt_193 | maskExt_193 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h30)
        v0_194 <= v0_194 & ~maskExt_194 | maskExt_194 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h30)
        v0_195 <= v0_195 & ~maskExt_195 | maskExt_195 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h31)
        v0_196 <= v0_196 & ~maskExt_196 | maskExt_196 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h31)
        v0_197 <= v0_197 & ~maskExt_197 | maskExt_197 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h31)
        v0_198 <= v0_198 & ~maskExt_198 | maskExt_198 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h31)
        v0_199 <= v0_199 & ~maskExt_199 | maskExt_199 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h32)
        v0_200 <= v0_200 & ~maskExt_200 | maskExt_200 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h32)
        v0_201 <= v0_201 & ~maskExt_201 | maskExt_201 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h32)
        v0_202 <= v0_202 & ~maskExt_202 | maskExt_202 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h32)
        v0_203 <= v0_203 & ~maskExt_203 | maskExt_203 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h33)
        v0_204 <= v0_204 & ~maskExt_204 | maskExt_204 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h33)
        v0_205 <= v0_205 & ~maskExt_205 | maskExt_205 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h33)
        v0_206 <= v0_206 & ~maskExt_206 | maskExt_206 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h33)
        v0_207 <= v0_207 & ~maskExt_207 | maskExt_207 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h34)
        v0_208 <= v0_208 & ~maskExt_208 | maskExt_208 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h34)
        v0_209 <= v0_209 & ~maskExt_209 | maskExt_209 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h34)
        v0_210 <= v0_210 & ~maskExt_210 | maskExt_210 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h34)
        v0_211 <= v0_211 & ~maskExt_211 | maskExt_211 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h35)
        v0_212 <= v0_212 & ~maskExt_212 | maskExt_212 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h35)
        v0_213 <= v0_213 & ~maskExt_213 | maskExt_213 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h35)
        v0_214 <= v0_214 & ~maskExt_214 | maskExt_214 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h35)
        v0_215 <= v0_215 & ~maskExt_215 | maskExt_215 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h36)
        v0_216 <= v0_216 & ~maskExt_216 | maskExt_216 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h36)
        v0_217 <= v0_217 & ~maskExt_217 | maskExt_217 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h36)
        v0_218 <= v0_218 & ~maskExt_218 | maskExt_218 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h36)
        v0_219 <= v0_219 & ~maskExt_219 | maskExt_219 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h37)
        v0_220 <= v0_220 & ~maskExt_220 | maskExt_220 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h37)
        v0_221 <= v0_221 & ~maskExt_221 | maskExt_221 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h37)
        v0_222 <= v0_222 & ~maskExt_222 | maskExt_222 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h37)
        v0_223 <= v0_223 & ~maskExt_223 | maskExt_223 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h38)
        v0_224 <= v0_224 & ~maskExt_224 | maskExt_224 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h38)
        v0_225 <= v0_225 & ~maskExt_225 | maskExt_225 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h38)
        v0_226 <= v0_226 & ~maskExt_226 | maskExt_226 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h38)
        v0_227 <= v0_227 & ~maskExt_227 | maskExt_227 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h39)
        v0_228 <= v0_228 & ~maskExt_228 | maskExt_228 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h39)
        v0_229 <= v0_229 & ~maskExt_229 | maskExt_229 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h39)
        v0_230 <= v0_230 & ~maskExt_230 | maskExt_230 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h39)
        v0_231 <= v0_231 & ~maskExt_231 | maskExt_231 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h3A)
        v0_232 <= v0_232 & ~maskExt_232 | maskExt_232 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h3A)
        v0_233 <= v0_233 & ~maskExt_233 | maskExt_233 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h3A)
        v0_234 <= v0_234 & ~maskExt_234 | maskExt_234 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h3A)
        v0_235 <= v0_235 & ~maskExt_235 | maskExt_235 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h3B)
        v0_236 <= v0_236 & ~maskExt_236 | maskExt_236 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h3B)
        v0_237 <= v0_237 & ~maskExt_237 | maskExt_237 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h3B)
        v0_238 <= v0_238 & ~maskExt_238 | maskExt_238 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h3B)
        v0_239 <= v0_239 & ~maskExt_239 | maskExt_239 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h3C)
        v0_240 <= v0_240 & ~maskExt_240 | maskExt_240 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h3C)
        v0_241 <= v0_241 & ~maskExt_241 | maskExt_241 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h3C)
        v0_242 <= v0_242 & ~maskExt_242 | maskExt_242 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h3C)
        v0_243 <= v0_243 & ~maskExt_243 | maskExt_243 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h3D)
        v0_244 <= v0_244 & ~maskExt_244 | maskExt_244 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h3D)
        v0_245 <= v0_245 & ~maskExt_245 | maskExt_245 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h3D)
        v0_246 <= v0_246 & ~maskExt_246 | maskExt_246 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h3D)
        v0_247 <= v0_247 & ~maskExt_247 | maskExt_247 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h3E)
        v0_248 <= v0_248 & ~maskExt_248 | maskExt_248 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h3E)
        v0_249 <= v0_249 & ~maskExt_249 | maskExt_249 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h3E)
        v0_250 <= v0_250 & ~maskExt_250 | maskExt_250 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h3E)
        v0_251 <= v0_251 & ~maskExt_251 | maskExt_251 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h3F)
        v0_252 <= v0_252 & ~maskExt_252 | maskExt_252 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h3F)
        v0_253 <= v0_253 & ~maskExt_253 | maskExt_253 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h3F)
        v0_254 <= v0_254 & ~maskExt_254 | maskExt_254 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h3F)
        v0_255 <= v0_255 & ~maskExt_255 | maskExt_255 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h40)
        v0_256 <= v0_256 & ~maskExt_256 | maskExt_256 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h40)
        v0_257 <= v0_257 & ~maskExt_257 | maskExt_257 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h40)
        v0_258 <= v0_258 & ~maskExt_258 | maskExt_258 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h40)
        v0_259 <= v0_259 & ~maskExt_259 | maskExt_259 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h41)
        v0_260 <= v0_260 & ~maskExt_260 | maskExt_260 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h41)
        v0_261 <= v0_261 & ~maskExt_261 | maskExt_261 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h41)
        v0_262 <= v0_262 & ~maskExt_262 | maskExt_262 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h41)
        v0_263 <= v0_263 & ~maskExt_263 | maskExt_263 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h42)
        v0_264 <= v0_264 & ~maskExt_264 | maskExt_264 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h42)
        v0_265 <= v0_265 & ~maskExt_265 | maskExt_265 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h42)
        v0_266 <= v0_266 & ~maskExt_266 | maskExt_266 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h42)
        v0_267 <= v0_267 & ~maskExt_267 | maskExt_267 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h43)
        v0_268 <= v0_268 & ~maskExt_268 | maskExt_268 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h43)
        v0_269 <= v0_269 & ~maskExt_269 | maskExt_269 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h43)
        v0_270 <= v0_270 & ~maskExt_270 | maskExt_270 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h43)
        v0_271 <= v0_271 & ~maskExt_271 | maskExt_271 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h44)
        v0_272 <= v0_272 & ~maskExt_272 | maskExt_272 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h44)
        v0_273 <= v0_273 & ~maskExt_273 | maskExt_273 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h44)
        v0_274 <= v0_274 & ~maskExt_274 | maskExt_274 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h44)
        v0_275 <= v0_275 & ~maskExt_275 | maskExt_275 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h45)
        v0_276 <= v0_276 & ~maskExt_276 | maskExt_276 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h45)
        v0_277 <= v0_277 & ~maskExt_277 | maskExt_277 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h45)
        v0_278 <= v0_278 & ~maskExt_278 | maskExt_278 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h45)
        v0_279 <= v0_279 & ~maskExt_279 | maskExt_279 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h46)
        v0_280 <= v0_280 & ~maskExt_280 | maskExt_280 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h46)
        v0_281 <= v0_281 & ~maskExt_281 | maskExt_281 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h46)
        v0_282 <= v0_282 & ~maskExt_282 | maskExt_282 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h46)
        v0_283 <= v0_283 & ~maskExt_283 | maskExt_283 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h47)
        v0_284 <= v0_284 & ~maskExt_284 | maskExt_284 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h47)
        v0_285 <= v0_285 & ~maskExt_285 | maskExt_285 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h47)
        v0_286 <= v0_286 & ~maskExt_286 | maskExt_286 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h47)
        v0_287 <= v0_287 & ~maskExt_287 | maskExt_287 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h48)
        v0_288 <= v0_288 & ~maskExt_288 | maskExt_288 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h48)
        v0_289 <= v0_289 & ~maskExt_289 | maskExt_289 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h48)
        v0_290 <= v0_290 & ~maskExt_290 | maskExt_290 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h48)
        v0_291 <= v0_291 & ~maskExt_291 | maskExt_291 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h49)
        v0_292 <= v0_292 & ~maskExt_292 | maskExt_292 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h49)
        v0_293 <= v0_293 & ~maskExt_293 | maskExt_293 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h49)
        v0_294 <= v0_294 & ~maskExt_294 | maskExt_294 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h49)
        v0_295 <= v0_295 & ~maskExt_295 | maskExt_295 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h4A)
        v0_296 <= v0_296 & ~maskExt_296 | maskExt_296 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h4A)
        v0_297 <= v0_297 & ~maskExt_297 | maskExt_297 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h4A)
        v0_298 <= v0_298 & ~maskExt_298 | maskExt_298 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h4A)
        v0_299 <= v0_299 & ~maskExt_299 | maskExt_299 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h4B)
        v0_300 <= v0_300 & ~maskExt_300 | maskExt_300 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h4B)
        v0_301 <= v0_301 & ~maskExt_301 | maskExt_301 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h4B)
        v0_302 <= v0_302 & ~maskExt_302 | maskExt_302 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h4B)
        v0_303 <= v0_303 & ~maskExt_303 | maskExt_303 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h4C)
        v0_304 <= v0_304 & ~maskExt_304 | maskExt_304 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h4C)
        v0_305 <= v0_305 & ~maskExt_305 | maskExt_305 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h4C)
        v0_306 <= v0_306 & ~maskExt_306 | maskExt_306 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h4C)
        v0_307 <= v0_307 & ~maskExt_307 | maskExt_307 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h4D)
        v0_308 <= v0_308 & ~maskExt_308 | maskExt_308 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h4D)
        v0_309 <= v0_309 & ~maskExt_309 | maskExt_309 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h4D)
        v0_310 <= v0_310 & ~maskExt_310 | maskExt_310 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h4D)
        v0_311 <= v0_311 & ~maskExt_311 | maskExt_311 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h4E)
        v0_312 <= v0_312 & ~maskExt_312 | maskExt_312 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h4E)
        v0_313 <= v0_313 & ~maskExt_313 | maskExt_313 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h4E)
        v0_314 <= v0_314 & ~maskExt_314 | maskExt_314 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h4E)
        v0_315 <= v0_315 & ~maskExt_315 | maskExt_315 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h4F)
        v0_316 <= v0_316 & ~maskExt_316 | maskExt_316 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h4F)
        v0_317 <= v0_317 & ~maskExt_317 | maskExt_317 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h4F)
        v0_318 <= v0_318 & ~maskExt_318 | maskExt_318 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h4F)
        v0_319 <= v0_319 & ~maskExt_319 | maskExt_319 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h50)
        v0_320 <= v0_320 & ~maskExt_320 | maskExt_320 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h50)
        v0_321 <= v0_321 & ~maskExt_321 | maskExt_321 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h50)
        v0_322 <= v0_322 & ~maskExt_322 | maskExt_322 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h50)
        v0_323 <= v0_323 & ~maskExt_323 | maskExt_323 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h51)
        v0_324 <= v0_324 & ~maskExt_324 | maskExt_324 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h51)
        v0_325 <= v0_325 & ~maskExt_325 | maskExt_325 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h51)
        v0_326 <= v0_326 & ~maskExt_326 | maskExt_326 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h51)
        v0_327 <= v0_327 & ~maskExt_327 | maskExt_327 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h52)
        v0_328 <= v0_328 & ~maskExt_328 | maskExt_328 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h52)
        v0_329 <= v0_329 & ~maskExt_329 | maskExt_329 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h52)
        v0_330 <= v0_330 & ~maskExt_330 | maskExt_330 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h52)
        v0_331 <= v0_331 & ~maskExt_331 | maskExt_331 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h53)
        v0_332 <= v0_332 & ~maskExt_332 | maskExt_332 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h53)
        v0_333 <= v0_333 & ~maskExt_333 | maskExt_333 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h53)
        v0_334 <= v0_334 & ~maskExt_334 | maskExt_334 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h53)
        v0_335 <= v0_335 & ~maskExt_335 | maskExt_335 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h54)
        v0_336 <= v0_336 & ~maskExt_336 | maskExt_336 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h54)
        v0_337 <= v0_337 & ~maskExt_337 | maskExt_337 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h54)
        v0_338 <= v0_338 & ~maskExt_338 | maskExt_338 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h54)
        v0_339 <= v0_339 & ~maskExt_339 | maskExt_339 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h55)
        v0_340 <= v0_340 & ~maskExt_340 | maskExt_340 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h55)
        v0_341 <= v0_341 & ~maskExt_341 | maskExt_341 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h55)
        v0_342 <= v0_342 & ~maskExt_342 | maskExt_342 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h55)
        v0_343 <= v0_343 & ~maskExt_343 | maskExt_343 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h56)
        v0_344 <= v0_344 & ~maskExt_344 | maskExt_344 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h56)
        v0_345 <= v0_345 & ~maskExt_345 | maskExt_345 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h56)
        v0_346 <= v0_346 & ~maskExt_346 | maskExt_346 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h56)
        v0_347 <= v0_347 & ~maskExt_347 | maskExt_347 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h57)
        v0_348 <= v0_348 & ~maskExt_348 | maskExt_348 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h57)
        v0_349 <= v0_349 & ~maskExt_349 | maskExt_349 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h57)
        v0_350 <= v0_350 & ~maskExt_350 | maskExt_350 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h57)
        v0_351 <= v0_351 & ~maskExt_351 | maskExt_351 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h58)
        v0_352 <= v0_352 & ~maskExt_352 | maskExt_352 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h58)
        v0_353 <= v0_353 & ~maskExt_353 | maskExt_353 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h58)
        v0_354 <= v0_354 & ~maskExt_354 | maskExt_354 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h58)
        v0_355 <= v0_355 & ~maskExt_355 | maskExt_355 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h59)
        v0_356 <= v0_356 & ~maskExt_356 | maskExt_356 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h59)
        v0_357 <= v0_357 & ~maskExt_357 | maskExt_357 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h59)
        v0_358 <= v0_358 & ~maskExt_358 | maskExt_358 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h59)
        v0_359 <= v0_359 & ~maskExt_359 | maskExt_359 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h5A)
        v0_360 <= v0_360 & ~maskExt_360 | maskExt_360 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h5A)
        v0_361 <= v0_361 & ~maskExt_361 | maskExt_361 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h5A)
        v0_362 <= v0_362 & ~maskExt_362 | maskExt_362 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h5A)
        v0_363 <= v0_363 & ~maskExt_363 | maskExt_363 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h5B)
        v0_364 <= v0_364 & ~maskExt_364 | maskExt_364 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h5B)
        v0_365 <= v0_365 & ~maskExt_365 | maskExt_365 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h5B)
        v0_366 <= v0_366 & ~maskExt_366 | maskExt_366 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h5B)
        v0_367 <= v0_367 & ~maskExt_367 | maskExt_367 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h5C)
        v0_368 <= v0_368 & ~maskExt_368 | maskExt_368 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h5C)
        v0_369 <= v0_369 & ~maskExt_369 | maskExt_369 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h5C)
        v0_370 <= v0_370 & ~maskExt_370 | maskExt_370 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h5C)
        v0_371 <= v0_371 & ~maskExt_371 | maskExt_371 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h5D)
        v0_372 <= v0_372 & ~maskExt_372 | maskExt_372 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h5D)
        v0_373 <= v0_373 & ~maskExt_373 | maskExt_373 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h5D)
        v0_374 <= v0_374 & ~maskExt_374 | maskExt_374 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h5D)
        v0_375 <= v0_375 & ~maskExt_375 | maskExt_375 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h5E)
        v0_376 <= v0_376 & ~maskExt_376 | maskExt_376 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h5E)
        v0_377 <= v0_377 & ~maskExt_377 | maskExt_377 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h5E)
        v0_378 <= v0_378 & ~maskExt_378 | maskExt_378 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h5E)
        v0_379 <= v0_379 & ~maskExt_379 | maskExt_379 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h5F)
        v0_380 <= v0_380 & ~maskExt_380 | maskExt_380 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h5F)
        v0_381 <= v0_381 & ~maskExt_381 | maskExt_381 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h5F)
        v0_382 <= v0_382 & ~maskExt_382 | maskExt_382 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h5F)
        v0_383 <= v0_383 & ~maskExt_383 | maskExt_383 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h60)
        v0_384 <= v0_384 & ~maskExt_384 | maskExt_384 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h60)
        v0_385 <= v0_385 & ~maskExt_385 | maskExt_385 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h60)
        v0_386 <= v0_386 & ~maskExt_386 | maskExt_386 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h60)
        v0_387 <= v0_387 & ~maskExt_387 | maskExt_387 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h61)
        v0_388 <= v0_388 & ~maskExt_388 | maskExt_388 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h61)
        v0_389 <= v0_389 & ~maskExt_389 | maskExt_389 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h61)
        v0_390 <= v0_390 & ~maskExt_390 | maskExt_390 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h61)
        v0_391 <= v0_391 & ~maskExt_391 | maskExt_391 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h62)
        v0_392 <= v0_392 & ~maskExt_392 | maskExt_392 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h62)
        v0_393 <= v0_393 & ~maskExt_393 | maskExt_393 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h62)
        v0_394 <= v0_394 & ~maskExt_394 | maskExt_394 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h62)
        v0_395 <= v0_395 & ~maskExt_395 | maskExt_395 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h63)
        v0_396 <= v0_396 & ~maskExt_396 | maskExt_396 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h63)
        v0_397 <= v0_397 & ~maskExt_397 | maskExt_397 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h63)
        v0_398 <= v0_398 & ~maskExt_398 | maskExt_398 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h63)
        v0_399 <= v0_399 & ~maskExt_399 | maskExt_399 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h64)
        v0_400 <= v0_400 & ~maskExt_400 | maskExt_400 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h64)
        v0_401 <= v0_401 & ~maskExt_401 | maskExt_401 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h64)
        v0_402 <= v0_402 & ~maskExt_402 | maskExt_402 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h64)
        v0_403 <= v0_403 & ~maskExt_403 | maskExt_403 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h65)
        v0_404 <= v0_404 & ~maskExt_404 | maskExt_404 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h65)
        v0_405 <= v0_405 & ~maskExt_405 | maskExt_405 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h65)
        v0_406 <= v0_406 & ~maskExt_406 | maskExt_406 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h65)
        v0_407 <= v0_407 & ~maskExt_407 | maskExt_407 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h66)
        v0_408 <= v0_408 & ~maskExt_408 | maskExt_408 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h66)
        v0_409 <= v0_409 & ~maskExt_409 | maskExt_409 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h66)
        v0_410 <= v0_410 & ~maskExt_410 | maskExt_410 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h66)
        v0_411 <= v0_411 & ~maskExt_411 | maskExt_411 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h67)
        v0_412 <= v0_412 & ~maskExt_412 | maskExt_412 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h67)
        v0_413 <= v0_413 & ~maskExt_413 | maskExt_413 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h67)
        v0_414 <= v0_414 & ~maskExt_414 | maskExt_414 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h67)
        v0_415 <= v0_415 & ~maskExt_415 | maskExt_415 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h68)
        v0_416 <= v0_416 & ~maskExt_416 | maskExt_416 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h68)
        v0_417 <= v0_417 & ~maskExt_417 | maskExt_417 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h68)
        v0_418 <= v0_418 & ~maskExt_418 | maskExt_418 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h68)
        v0_419 <= v0_419 & ~maskExt_419 | maskExt_419 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h69)
        v0_420 <= v0_420 & ~maskExt_420 | maskExt_420 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h69)
        v0_421 <= v0_421 & ~maskExt_421 | maskExt_421 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h69)
        v0_422 <= v0_422 & ~maskExt_422 | maskExt_422 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h69)
        v0_423 <= v0_423 & ~maskExt_423 | maskExt_423 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h6A)
        v0_424 <= v0_424 & ~maskExt_424 | maskExt_424 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h6A)
        v0_425 <= v0_425 & ~maskExt_425 | maskExt_425 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h6A)
        v0_426 <= v0_426 & ~maskExt_426 | maskExt_426 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h6A)
        v0_427 <= v0_427 & ~maskExt_427 | maskExt_427 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h6B)
        v0_428 <= v0_428 & ~maskExt_428 | maskExt_428 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h6B)
        v0_429 <= v0_429 & ~maskExt_429 | maskExt_429 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h6B)
        v0_430 <= v0_430 & ~maskExt_430 | maskExt_430 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h6B)
        v0_431 <= v0_431 & ~maskExt_431 | maskExt_431 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h6C)
        v0_432 <= v0_432 & ~maskExt_432 | maskExt_432 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h6C)
        v0_433 <= v0_433 & ~maskExt_433 | maskExt_433 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h6C)
        v0_434 <= v0_434 & ~maskExt_434 | maskExt_434 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h6C)
        v0_435 <= v0_435 & ~maskExt_435 | maskExt_435 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h6D)
        v0_436 <= v0_436 & ~maskExt_436 | maskExt_436 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h6D)
        v0_437 <= v0_437 & ~maskExt_437 | maskExt_437 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h6D)
        v0_438 <= v0_438 & ~maskExt_438 | maskExt_438 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h6D)
        v0_439 <= v0_439 & ~maskExt_439 | maskExt_439 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h6E)
        v0_440 <= v0_440 & ~maskExt_440 | maskExt_440 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h6E)
        v0_441 <= v0_441 & ~maskExt_441 | maskExt_441 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h6E)
        v0_442 <= v0_442 & ~maskExt_442 | maskExt_442 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h6E)
        v0_443 <= v0_443 & ~maskExt_443 | maskExt_443 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h6F)
        v0_444 <= v0_444 & ~maskExt_444 | maskExt_444 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h6F)
        v0_445 <= v0_445 & ~maskExt_445 | maskExt_445 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h6F)
        v0_446 <= v0_446 & ~maskExt_446 | maskExt_446 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h6F)
        v0_447 <= v0_447 & ~maskExt_447 | maskExt_447 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h70)
        v0_448 <= v0_448 & ~maskExt_448 | maskExt_448 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h70)
        v0_449 <= v0_449 & ~maskExt_449 | maskExt_449 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h70)
        v0_450 <= v0_450 & ~maskExt_450 | maskExt_450 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h70)
        v0_451 <= v0_451 & ~maskExt_451 | maskExt_451 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h71)
        v0_452 <= v0_452 & ~maskExt_452 | maskExt_452 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h71)
        v0_453 <= v0_453 & ~maskExt_453 | maskExt_453 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h71)
        v0_454 <= v0_454 & ~maskExt_454 | maskExt_454 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h71)
        v0_455 <= v0_455 & ~maskExt_455 | maskExt_455 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h72)
        v0_456 <= v0_456 & ~maskExt_456 | maskExt_456 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h72)
        v0_457 <= v0_457 & ~maskExt_457 | maskExt_457 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h72)
        v0_458 <= v0_458 & ~maskExt_458 | maskExt_458 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h72)
        v0_459 <= v0_459 & ~maskExt_459 | maskExt_459 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h73)
        v0_460 <= v0_460 & ~maskExt_460 | maskExt_460 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h73)
        v0_461 <= v0_461 & ~maskExt_461 | maskExt_461 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h73)
        v0_462 <= v0_462 & ~maskExt_462 | maskExt_462 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h73)
        v0_463 <= v0_463 & ~maskExt_463 | maskExt_463 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h74)
        v0_464 <= v0_464 & ~maskExt_464 | maskExt_464 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h74)
        v0_465 <= v0_465 & ~maskExt_465 | maskExt_465 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h74)
        v0_466 <= v0_466 & ~maskExt_466 | maskExt_466 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h74)
        v0_467 <= v0_467 & ~maskExt_467 | maskExt_467 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h75)
        v0_468 <= v0_468 & ~maskExt_468 | maskExt_468 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h75)
        v0_469 <= v0_469 & ~maskExt_469 | maskExt_469 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h75)
        v0_470 <= v0_470 & ~maskExt_470 | maskExt_470 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h75)
        v0_471 <= v0_471 & ~maskExt_471 | maskExt_471 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h76)
        v0_472 <= v0_472 & ~maskExt_472 | maskExt_472 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h76)
        v0_473 <= v0_473 & ~maskExt_473 | maskExt_473 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h76)
        v0_474 <= v0_474 & ~maskExt_474 | maskExt_474 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h76)
        v0_475 <= v0_475 & ~maskExt_475 | maskExt_475 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h77)
        v0_476 <= v0_476 & ~maskExt_476 | maskExt_476 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h77)
        v0_477 <= v0_477 & ~maskExt_477 | maskExt_477 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h77)
        v0_478 <= v0_478 & ~maskExt_478 | maskExt_478 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h77)
        v0_479 <= v0_479 & ~maskExt_479 | maskExt_479 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h78)
        v0_480 <= v0_480 & ~maskExt_480 | maskExt_480 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h78)
        v0_481 <= v0_481 & ~maskExt_481 | maskExt_481 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h78)
        v0_482 <= v0_482 & ~maskExt_482 | maskExt_482 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h78)
        v0_483 <= v0_483 & ~maskExt_483 | maskExt_483 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h79)
        v0_484 <= v0_484 & ~maskExt_484 | maskExt_484 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h79)
        v0_485 <= v0_485 & ~maskExt_485 | maskExt_485 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h79)
        v0_486 <= v0_486 & ~maskExt_486 | maskExt_486 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h79)
        v0_487 <= v0_487 & ~maskExt_487 | maskExt_487 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h7A)
        v0_488 <= v0_488 & ~maskExt_488 | maskExt_488 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h7A)
        v0_489 <= v0_489 & ~maskExt_489 | maskExt_489 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h7A)
        v0_490 <= v0_490 & ~maskExt_490 | maskExt_490 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h7A)
        v0_491 <= v0_491 & ~maskExt_491 | maskExt_491 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h7B)
        v0_492 <= v0_492 & ~maskExt_492 | maskExt_492 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h7B)
        v0_493 <= v0_493 & ~maskExt_493 | maskExt_493 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h7B)
        v0_494 <= v0_494 & ~maskExt_494 | maskExt_494 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h7B)
        v0_495 <= v0_495 & ~maskExt_495 | maskExt_495 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h7C)
        v0_496 <= v0_496 & ~maskExt_496 | maskExt_496 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h7C)
        v0_497 <= v0_497 & ~maskExt_497 | maskExt_497 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h7C)
        v0_498 <= v0_498 & ~maskExt_498 | maskExt_498 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h7C)
        v0_499 <= v0_499 & ~maskExt_499 | maskExt_499 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h7D)
        v0_500 <= v0_500 & ~maskExt_500 | maskExt_500 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h7D)
        v0_501 <= v0_501 & ~maskExt_501 | maskExt_501 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h7D)
        v0_502 <= v0_502 & ~maskExt_502 | maskExt_502 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h7D)
        v0_503 <= v0_503 & ~maskExt_503 | maskExt_503 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h7E)
        v0_504 <= v0_504 & ~maskExt_504 | maskExt_504 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h7E)
        v0_505 <= v0_505 & ~maskExt_505 | maskExt_505 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h7E)
        v0_506 <= v0_506 & ~maskExt_506 | maskExt_506 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h7E)
        v0_507 <= v0_507 & ~maskExt_507 | maskExt_507 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h7F)
        v0_508 <= v0_508 & ~maskExt_508 | maskExt_508 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h7F)
        v0_509 <= v0_509 & ~maskExt_509 | maskExt_509 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h7F)
        v0_510 <= v0_510 & ~maskExt_510 | maskExt_510 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h7F)
        v0_511 <= v0_511 & ~maskExt_511 | maskExt_511 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h80)
        v0_512 <= v0_512 & ~maskExt_512 | maskExt_512 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h80)
        v0_513 <= v0_513 & ~maskExt_513 | maskExt_513 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h80)
        v0_514 <= v0_514 & ~maskExt_514 | maskExt_514 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h80)
        v0_515 <= v0_515 & ~maskExt_515 | maskExt_515 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h81)
        v0_516 <= v0_516 & ~maskExt_516 | maskExt_516 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h81)
        v0_517 <= v0_517 & ~maskExt_517 | maskExt_517 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h81)
        v0_518 <= v0_518 & ~maskExt_518 | maskExt_518 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h81)
        v0_519 <= v0_519 & ~maskExt_519 | maskExt_519 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h82)
        v0_520 <= v0_520 & ~maskExt_520 | maskExt_520 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h82)
        v0_521 <= v0_521 & ~maskExt_521 | maskExt_521 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h82)
        v0_522 <= v0_522 & ~maskExt_522 | maskExt_522 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h82)
        v0_523 <= v0_523 & ~maskExt_523 | maskExt_523 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h83)
        v0_524 <= v0_524 & ~maskExt_524 | maskExt_524 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h83)
        v0_525 <= v0_525 & ~maskExt_525 | maskExt_525 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h83)
        v0_526 <= v0_526 & ~maskExt_526 | maskExt_526 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h83)
        v0_527 <= v0_527 & ~maskExt_527 | maskExt_527 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h84)
        v0_528 <= v0_528 & ~maskExt_528 | maskExt_528 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h84)
        v0_529 <= v0_529 & ~maskExt_529 | maskExt_529 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h84)
        v0_530 <= v0_530 & ~maskExt_530 | maskExt_530 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h84)
        v0_531 <= v0_531 & ~maskExt_531 | maskExt_531 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h85)
        v0_532 <= v0_532 & ~maskExt_532 | maskExt_532 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h85)
        v0_533 <= v0_533 & ~maskExt_533 | maskExt_533 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h85)
        v0_534 <= v0_534 & ~maskExt_534 | maskExt_534 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h85)
        v0_535 <= v0_535 & ~maskExt_535 | maskExt_535 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h86)
        v0_536 <= v0_536 & ~maskExt_536 | maskExt_536 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h86)
        v0_537 <= v0_537 & ~maskExt_537 | maskExt_537 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h86)
        v0_538 <= v0_538 & ~maskExt_538 | maskExt_538 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h86)
        v0_539 <= v0_539 & ~maskExt_539 | maskExt_539 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h87)
        v0_540 <= v0_540 & ~maskExt_540 | maskExt_540 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h87)
        v0_541 <= v0_541 & ~maskExt_541 | maskExt_541 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h87)
        v0_542 <= v0_542 & ~maskExt_542 | maskExt_542 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h87)
        v0_543 <= v0_543 & ~maskExt_543 | maskExt_543 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h88)
        v0_544 <= v0_544 & ~maskExt_544 | maskExt_544 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h88)
        v0_545 <= v0_545 & ~maskExt_545 | maskExt_545 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h88)
        v0_546 <= v0_546 & ~maskExt_546 | maskExt_546 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h88)
        v0_547 <= v0_547 & ~maskExt_547 | maskExt_547 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h89)
        v0_548 <= v0_548 & ~maskExt_548 | maskExt_548 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h89)
        v0_549 <= v0_549 & ~maskExt_549 | maskExt_549 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h89)
        v0_550 <= v0_550 & ~maskExt_550 | maskExt_550 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h89)
        v0_551 <= v0_551 & ~maskExt_551 | maskExt_551 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h8A)
        v0_552 <= v0_552 & ~maskExt_552 | maskExt_552 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h8A)
        v0_553 <= v0_553 & ~maskExt_553 | maskExt_553 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h8A)
        v0_554 <= v0_554 & ~maskExt_554 | maskExt_554 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h8A)
        v0_555 <= v0_555 & ~maskExt_555 | maskExt_555 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h8B)
        v0_556 <= v0_556 & ~maskExt_556 | maskExt_556 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h8B)
        v0_557 <= v0_557 & ~maskExt_557 | maskExt_557 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h8B)
        v0_558 <= v0_558 & ~maskExt_558 | maskExt_558 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h8B)
        v0_559 <= v0_559 & ~maskExt_559 | maskExt_559 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h8C)
        v0_560 <= v0_560 & ~maskExt_560 | maskExt_560 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h8C)
        v0_561 <= v0_561 & ~maskExt_561 | maskExt_561 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h8C)
        v0_562 <= v0_562 & ~maskExt_562 | maskExt_562 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h8C)
        v0_563 <= v0_563 & ~maskExt_563 | maskExt_563 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h8D)
        v0_564 <= v0_564 & ~maskExt_564 | maskExt_564 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h8D)
        v0_565 <= v0_565 & ~maskExt_565 | maskExt_565 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h8D)
        v0_566 <= v0_566 & ~maskExt_566 | maskExt_566 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h8D)
        v0_567 <= v0_567 & ~maskExt_567 | maskExt_567 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h8E)
        v0_568 <= v0_568 & ~maskExt_568 | maskExt_568 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h8E)
        v0_569 <= v0_569 & ~maskExt_569 | maskExt_569 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h8E)
        v0_570 <= v0_570 & ~maskExt_570 | maskExt_570 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h8E)
        v0_571 <= v0_571 & ~maskExt_571 | maskExt_571 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h8F)
        v0_572 <= v0_572 & ~maskExt_572 | maskExt_572 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h8F)
        v0_573 <= v0_573 & ~maskExt_573 | maskExt_573 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h8F)
        v0_574 <= v0_574 & ~maskExt_574 | maskExt_574 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h8F)
        v0_575 <= v0_575 & ~maskExt_575 | maskExt_575 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h90)
        v0_576 <= v0_576 & ~maskExt_576 | maskExt_576 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h90)
        v0_577 <= v0_577 & ~maskExt_577 | maskExt_577 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h90)
        v0_578 <= v0_578 & ~maskExt_578 | maskExt_578 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h90)
        v0_579 <= v0_579 & ~maskExt_579 | maskExt_579 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h91)
        v0_580 <= v0_580 & ~maskExt_580 | maskExt_580 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h91)
        v0_581 <= v0_581 & ~maskExt_581 | maskExt_581 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h91)
        v0_582 <= v0_582 & ~maskExt_582 | maskExt_582 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h91)
        v0_583 <= v0_583 & ~maskExt_583 | maskExt_583 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h92)
        v0_584 <= v0_584 & ~maskExt_584 | maskExt_584 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h92)
        v0_585 <= v0_585 & ~maskExt_585 | maskExt_585 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h92)
        v0_586 <= v0_586 & ~maskExt_586 | maskExt_586 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h92)
        v0_587 <= v0_587 & ~maskExt_587 | maskExt_587 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h93)
        v0_588 <= v0_588 & ~maskExt_588 | maskExt_588 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h93)
        v0_589 <= v0_589 & ~maskExt_589 | maskExt_589 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h93)
        v0_590 <= v0_590 & ~maskExt_590 | maskExt_590 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h93)
        v0_591 <= v0_591 & ~maskExt_591 | maskExt_591 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h94)
        v0_592 <= v0_592 & ~maskExt_592 | maskExt_592 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h94)
        v0_593 <= v0_593 & ~maskExt_593 | maskExt_593 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h94)
        v0_594 <= v0_594 & ~maskExt_594 | maskExt_594 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h94)
        v0_595 <= v0_595 & ~maskExt_595 | maskExt_595 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h95)
        v0_596 <= v0_596 & ~maskExt_596 | maskExt_596 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h95)
        v0_597 <= v0_597 & ~maskExt_597 | maskExt_597 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h95)
        v0_598 <= v0_598 & ~maskExt_598 | maskExt_598 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h95)
        v0_599 <= v0_599 & ~maskExt_599 | maskExt_599 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h96)
        v0_600 <= v0_600 & ~maskExt_600 | maskExt_600 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h96)
        v0_601 <= v0_601 & ~maskExt_601 | maskExt_601 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h96)
        v0_602 <= v0_602 & ~maskExt_602 | maskExt_602 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h96)
        v0_603 <= v0_603 & ~maskExt_603 | maskExt_603 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h97)
        v0_604 <= v0_604 & ~maskExt_604 | maskExt_604 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h97)
        v0_605 <= v0_605 & ~maskExt_605 | maskExt_605 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h97)
        v0_606 <= v0_606 & ~maskExt_606 | maskExt_606 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h97)
        v0_607 <= v0_607 & ~maskExt_607 | maskExt_607 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h98)
        v0_608 <= v0_608 & ~maskExt_608 | maskExt_608 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h98)
        v0_609 <= v0_609 & ~maskExt_609 | maskExt_609 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h98)
        v0_610 <= v0_610 & ~maskExt_610 | maskExt_610 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h98)
        v0_611 <= v0_611 & ~maskExt_611 | maskExt_611 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h99)
        v0_612 <= v0_612 & ~maskExt_612 | maskExt_612 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h99)
        v0_613 <= v0_613 & ~maskExt_613 | maskExt_613 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h99)
        v0_614 <= v0_614 & ~maskExt_614 | maskExt_614 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h99)
        v0_615 <= v0_615 & ~maskExt_615 | maskExt_615 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h9A)
        v0_616 <= v0_616 & ~maskExt_616 | maskExt_616 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h9A)
        v0_617 <= v0_617 & ~maskExt_617 | maskExt_617 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h9A)
        v0_618 <= v0_618 & ~maskExt_618 | maskExt_618 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h9A)
        v0_619 <= v0_619 & ~maskExt_619 | maskExt_619 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h9B)
        v0_620 <= v0_620 & ~maskExt_620 | maskExt_620 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h9B)
        v0_621 <= v0_621 & ~maskExt_621 | maskExt_621 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h9B)
        v0_622 <= v0_622 & ~maskExt_622 | maskExt_622 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h9B)
        v0_623 <= v0_623 & ~maskExt_623 | maskExt_623 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h9C)
        v0_624 <= v0_624 & ~maskExt_624 | maskExt_624 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h9C)
        v0_625 <= v0_625 & ~maskExt_625 | maskExt_625 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h9C)
        v0_626 <= v0_626 & ~maskExt_626 | maskExt_626 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h9C)
        v0_627 <= v0_627 & ~maskExt_627 | maskExt_627 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h9D)
        v0_628 <= v0_628 & ~maskExt_628 | maskExt_628 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h9D)
        v0_629 <= v0_629 & ~maskExt_629 | maskExt_629 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h9D)
        v0_630 <= v0_630 & ~maskExt_630 | maskExt_630 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h9D)
        v0_631 <= v0_631 & ~maskExt_631 | maskExt_631 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h9E)
        v0_632 <= v0_632 & ~maskExt_632 | maskExt_632 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h9E)
        v0_633 <= v0_633 & ~maskExt_633 | maskExt_633 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h9E)
        v0_634 <= v0_634 & ~maskExt_634 | maskExt_634 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h9E)
        v0_635 <= v0_635 & ~maskExt_635 | maskExt_635 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h9F)
        v0_636 <= v0_636 & ~maskExt_636 | maskExt_636 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h9F)
        v0_637 <= v0_637 & ~maskExt_637 | maskExt_637 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h9F)
        v0_638 <= v0_638 & ~maskExt_638 | maskExt_638 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h9F)
        v0_639 <= v0_639 & ~maskExt_639 | maskExt_639 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hA0)
        v0_640 <= v0_640 & ~maskExt_640 | maskExt_640 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hA0)
        v0_641 <= v0_641 & ~maskExt_641 | maskExt_641 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hA0)
        v0_642 <= v0_642 & ~maskExt_642 | maskExt_642 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hA0)
        v0_643 <= v0_643 & ~maskExt_643 | maskExt_643 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hA1)
        v0_644 <= v0_644 & ~maskExt_644 | maskExt_644 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hA1)
        v0_645 <= v0_645 & ~maskExt_645 | maskExt_645 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hA1)
        v0_646 <= v0_646 & ~maskExt_646 | maskExt_646 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hA1)
        v0_647 <= v0_647 & ~maskExt_647 | maskExt_647 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hA2)
        v0_648 <= v0_648 & ~maskExt_648 | maskExt_648 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hA2)
        v0_649 <= v0_649 & ~maskExt_649 | maskExt_649 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hA2)
        v0_650 <= v0_650 & ~maskExt_650 | maskExt_650 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hA2)
        v0_651 <= v0_651 & ~maskExt_651 | maskExt_651 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hA3)
        v0_652 <= v0_652 & ~maskExt_652 | maskExt_652 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hA3)
        v0_653 <= v0_653 & ~maskExt_653 | maskExt_653 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hA3)
        v0_654 <= v0_654 & ~maskExt_654 | maskExt_654 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hA3)
        v0_655 <= v0_655 & ~maskExt_655 | maskExt_655 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hA4)
        v0_656 <= v0_656 & ~maskExt_656 | maskExt_656 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hA4)
        v0_657 <= v0_657 & ~maskExt_657 | maskExt_657 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hA4)
        v0_658 <= v0_658 & ~maskExt_658 | maskExt_658 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hA4)
        v0_659 <= v0_659 & ~maskExt_659 | maskExt_659 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hA5)
        v0_660 <= v0_660 & ~maskExt_660 | maskExt_660 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hA5)
        v0_661 <= v0_661 & ~maskExt_661 | maskExt_661 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hA5)
        v0_662 <= v0_662 & ~maskExt_662 | maskExt_662 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hA5)
        v0_663 <= v0_663 & ~maskExt_663 | maskExt_663 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hA6)
        v0_664 <= v0_664 & ~maskExt_664 | maskExt_664 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hA6)
        v0_665 <= v0_665 & ~maskExt_665 | maskExt_665 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hA6)
        v0_666 <= v0_666 & ~maskExt_666 | maskExt_666 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hA6)
        v0_667 <= v0_667 & ~maskExt_667 | maskExt_667 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hA7)
        v0_668 <= v0_668 & ~maskExt_668 | maskExt_668 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hA7)
        v0_669 <= v0_669 & ~maskExt_669 | maskExt_669 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hA7)
        v0_670 <= v0_670 & ~maskExt_670 | maskExt_670 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hA7)
        v0_671 <= v0_671 & ~maskExt_671 | maskExt_671 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hA8)
        v0_672 <= v0_672 & ~maskExt_672 | maskExt_672 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hA8)
        v0_673 <= v0_673 & ~maskExt_673 | maskExt_673 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hA8)
        v0_674 <= v0_674 & ~maskExt_674 | maskExt_674 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hA8)
        v0_675 <= v0_675 & ~maskExt_675 | maskExt_675 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hA9)
        v0_676 <= v0_676 & ~maskExt_676 | maskExt_676 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hA9)
        v0_677 <= v0_677 & ~maskExt_677 | maskExt_677 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hA9)
        v0_678 <= v0_678 & ~maskExt_678 | maskExt_678 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hA9)
        v0_679 <= v0_679 & ~maskExt_679 | maskExt_679 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hAA)
        v0_680 <= v0_680 & ~maskExt_680 | maskExt_680 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hAA)
        v0_681 <= v0_681 & ~maskExt_681 | maskExt_681 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hAA)
        v0_682 <= v0_682 & ~maskExt_682 | maskExt_682 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hAA)
        v0_683 <= v0_683 & ~maskExt_683 | maskExt_683 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hAB)
        v0_684 <= v0_684 & ~maskExt_684 | maskExt_684 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hAB)
        v0_685 <= v0_685 & ~maskExt_685 | maskExt_685 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hAB)
        v0_686 <= v0_686 & ~maskExt_686 | maskExt_686 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hAB)
        v0_687 <= v0_687 & ~maskExt_687 | maskExt_687 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hAC)
        v0_688 <= v0_688 & ~maskExt_688 | maskExt_688 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hAC)
        v0_689 <= v0_689 & ~maskExt_689 | maskExt_689 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hAC)
        v0_690 <= v0_690 & ~maskExt_690 | maskExt_690 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hAC)
        v0_691 <= v0_691 & ~maskExt_691 | maskExt_691 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hAD)
        v0_692 <= v0_692 & ~maskExt_692 | maskExt_692 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hAD)
        v0_693 <= v0_693 & ~maskExt_693 | maskExt_693 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hAD)
        v0_694 <= v0_694 & ~maskExt_694 | maskExt_694 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hAD)
        v0_695 <= v0_695 & ~maskExt_695 | maskExt_695 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hAE)
        v0_696 <= v0_696 & ~maskExt_696 | maskExt_696 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hAE)
        v0_697 <= v0_697 & ~maskExt_697 | maskExt_697 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hAE)
        v0_698 <= v0_698 & ~maskExt_698 | maskExt_698 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hAE)
        v0_699 <= v0_699 & ~maskExt_699 | maskExt_699 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hAF)
        v0_700 <= v0_700 & ~maskExt_700 | maskExt_700 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hAF)
        v0_701 <= v0_701 & ~maskExt_701 | maskExt_701 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hAF)
        v0_702 <= v0_702 & ~maskExt_702 | maskExt_702 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hAF)
        v0_703 <= v0_703 & ~maskExt_703 | maskExt_703 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hB0)
        v0_704 <= v0_704 & ~maskExt_704 | maskExt_704 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hB0)
        v0_705 <= v0_705 & ~maskExt_705 | maskExt_705 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hB0)
        v0_706 <= v0_706 & ~maskExt_706 | maskExt_706 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hB0)
        v0_707 <= v0_707 & ~maskExt_707 | maskExt_707 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hB1)
        v0_708 <= v0_708 & ~maskExt_708 | maskExt_708 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hB1)
        v0_709 <= v0_709 & ~maskExt_709 | maskExt_709 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hB1)
        v0_710 <= v0_710 & ~maskExt_710 | maskExt_710 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hB1)
        v0_711 <= v0_711 & ~maskExt_711 | maskExt_711 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hB2)
        v0_712 <= v0_712 & ~maskExt_712 | maskExt_712 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hB2)
        v0_713 <= v0_713 & ~maskExt_713 | maskExt_713 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hB2)
        v0_714 <= v0_714 & ~maskExt_714 | maskExt_714 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hB2)
        v0_715 <= v0_715 & ~maskExt_715 | maskExt_715 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hB3)
        v0_716 <= v0_716 & ~maskExt_716 | maskExt_716 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hB3)
        v0_717 <= v0_717 & ~maskExt_717 | maskExt_717 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hB3)
        v0_718 <= v0_718 & ~maskExt_718 | maskExt_718 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hB3)
        v0_719 <= v0_719 & ~maskExt_719 | maskExt_719 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hB4)
        v0_720 <= v0_720 & ~maskExt_720 | maskExt_720 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hB4)
        v0_721 <= v0_721 & ~maskExt_721 | maskExt_721 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hB4)
        v0_722 <= v0_722 & ~maskExt_722 | maskExt_722 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hB4)
        v0_723 <= v0_723 & ~maskExt_723 | maskExt_723 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hB5)
        v0_724 <= v0_724 & ~maskExt_724 | maskExt_724 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hB5)
        v0_725 <= v0_725 & ~maskExt_725 | maskExt_725 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hB5)
        v0_726 <= v0_726 & ~maskExt_726 | maskExt_726 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hB5)
        v0_727 <= v0_727 & ~maskExt_727 | maskExt_727 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hB6)
        v0_728 <= v0_728 & ~maskExt_728 | maskExt_728 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hB6)
        v0_729 <= v0_729 & ~maskExt_729 | maskExt_729 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hB6)
        v0_730 <= v0_730 & ~maskExt_730 | maskExt_730 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hB6)
        v0_731 <= v0_731 & ~maskExt_731 | maskExt_731 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hB7)
        v0_732 <= v0_732 & ~maskExt_732 | maskExt_732 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hB7)
        v0_733 <= v0_733 & ~maskExt_733 | maskExt_733 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hB7)
        v0_734 <= v0_734 & ~maskExt_734 | maskExt_734 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hB7)
        v0_735 <= v0_735 & ~maskExt_735 | maskExt_735 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hB8)
        v0_736 <= v0_736 & ~maskExt_736 | maskExt_736 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hB8)
        v0_737 <= v0_737 & ~maskExt_737 | maskExt_737 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hB8)
        v0_738 <= v0_738 & ~maskExt_738 | maskExt_738 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hB8)
        v0_739 <= v0_739 & ~maskExt_739 | maskExt_739 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hB9)
        v0_740 <= v0_740 & ~maskExt_740 | maskExt_740 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hB9)
        v0_741 <= v0_741 & ~maskExt_741 | maskExt_741 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hB9)
        v0_742 <= v0_742 & ~maskExt_742 | maskExt_742 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hB9)
        v0_743 <= v0_743 & ~maskExt_743 | maskExt_743 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hBA)
        v0_744 <= v0_744 & ~maskExt_744 | maskExt_744 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hBA)
        v0_745 <= v0_745 & ~maskExt_745 | maskExt_745 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hBA)
        v0_746 <= v0_746 & ~maskExt_746 | maskExt_746 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hBA)
        v0_747 <= v0_747 & ~maskExt_747 | maskExt_747 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hBB)
        v0_748 <= v0_748 & ~maskExt_748 | maskExt_748 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hBB)
        v0_749 <= v0_749 & ~maskExt_749 | maskExt_749 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hBB)
        v0_750 <= v0_750 & ~maskExt_750 | maskExt_750 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hBB)
        v0_751 <= v0_751 & ~maskExt_751 | maskExt_751 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hBC)
        v0_752 <= v0_752 & ~maskExt_752 | maskExt_752 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hBC)
        v0_753 <= v0_753 & ~maskExt_753 | maskExt_753 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hBC)
        v0_754 <= v0_754 & ~maskExt_754 | maskExt_754 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hBC)
        v0_755 <= v0_755 & ~maskExt_755 | maskExt_755 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hBD)
        v0_756 <= v0_756 & ~maskExt_756 | maskExt_756 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hBD)
        v0_757 <= v0_757 & ~maskExt_757 | maskExt_757 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hBD)
        v0_758 <= v0_758 & ~maskExt_758 | maskExt_758 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hBD)
        v0_759 <= v0_759 & ~maskExt_759 | maskExt_759 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hBE)
        v0_760 <= v0_760 & ~maskExt_760 | maskExt_760 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hBE)
        v0_761 <= v0_761 & ~maskExt_761 | maskExt_761 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hBE)
        v0_762 <= v0_762 & ~maskExt_762 | maskExt_762 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hBE)
        v0_763 <= v0_763 & ~maskExt_763 | maskExt_763 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hBF)
        v0_764 <= v0_764 & ~maskExt_764 | maskExt_764 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hBF)
        v0_765 <= v0_765 & ~maskExt_765 | maskExt_765 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hBF)
        v0_766 <= v0_766 & ~maskExt_766 | maskExt_766 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hBF)
        v0_767 <= v0_767 & ~maskExt_767 | maskExt_767 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hC0)
        v0_768 <= v0_768 & ~maskExt_768 | maskExt_768 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hC0)
        v0_769 <= v0_769 & ~maskExt_769 | maskExt_769 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hC0)
        v0_770 <= v0_770 & ~maskExt_770 | maskExt_770 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hC0)
        v0_771 <= v0_771 & ~maskExt_771 | maskExt_771 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hC1)
        v0_772 <= v0_772 & ~maskExt_772 | maskExt_772 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hC1)
        v0_773 <= v0_773 & ~maskExt_773 | maskExt_773 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hC1)
        v0_774 <= v0_774 & ~maskExt_774 | maskExt_774 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hC1)
        v0_775 <= v0_775 & ~maskExt_775 | maskExt_775 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hC2)
        v0_776 <= v0_776 & ~maskExt_776 | maskExt_776 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hC2)
        v0_777 <= v0_777 & ~maskExt_777 | maskExt_777 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hC2)
        v0_778 <= v0_778 & ~maskExt_778 | maskExt_778 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hC2)
        v0_779 <= v0_779 & ~maskExt_779 | maskExt_779 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hC3)
        v0_780 <= v0_780 & ~maskExt_780 | maskExt_780 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hC3)
        v0_781 <= v0_781 & ~maskExt_781 | maskExt_781 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hC3)
        v0_782 <= v0_782 & ~maskExt_782 | maskExt_782 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hC3)
        v0_783 <= v0_783 & ~maskExt_783 | maskExt_783 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hC4)
        v0_784 <= v0_784 & ~maskExt_784 | maskExt_784 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hC4)
        v0_785 <= v0_785 & ~maskExt_785 | maskExt_785 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hC4)
        v0_786 <= v0_786 & ~maskExt_786 | maskExt_786 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hC4)
        v0_787 <= v0_787 & ~maskExt_787 | maskExt_787 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hC5)
        v0_788 <= v0_788 & ~maskExt_788 | maskExt_788 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hC5)
        v0_789 <= v0_789 & ~maskExt_789 | maskExt_789 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hC5)
        v0_790 <= v0_790 & ~maskExt_790 | maskExt_790 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hC5)
        v0_791 <= v0_791 & ~maskExt_791 | maskExt_791 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hC6)
        v0_792 <= v0_792 & ~maskExt_792 | maskExt_792 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hC6)
        v0_793 <= v0_793 & ~maskExt_793 | maskExt_793 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hC6)
        v0_794 <= v0_794 & ~maskExt_794 | maskExt_794 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hC6)
        v0_795 <= v0_795 & ~maskExt_795 | maskExt_795 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hC7)
        v0_796 <= v0_796 & ~maskExt_796 | maskExt_796 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hC7)
        v0_797 <= v0_797 & ~maskExt_797 | maskExt_797 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hC7)
        v0_798 <= v0_798 & ~maskExt_798 | maskExt_798 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hC7)
        v0_799 <= v0_799 & ~maskExt_799 | maskExt_799 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hC8)
        v0_800 <= v0_800 & ~maskExt_800 | maskExt_800 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hC8)
        v0_801 <= v0_801 & ~maskExt_801 | maskExt_801 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hC8)
        v0_802 <= v0_802 & ~maskExt_802 | maskExt_802 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hC8)
        v0_803 <= v0_803 & ~maskExt_803 | maskExt_803 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hC9)
        v0_804 <= v0_804 & ~maskExt_804 | maskExt_804 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hC9)
        v0_805 <= v0_805 & ~maskExt_805 | maskExt_805 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hC9)
        v0_806 <= v0_806 & ~maskExt_806 | maskExt_806 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hC9)
        v0_807 <= v0_807 & ~maskExt_807 | maskExt_807 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hCA)
        v0_808 <= v0_808 & ~maskExt_808 | maskExt_808 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hCA)
        v0_809 <= v0_809 & ~maskExt_809 | maskExt_809 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hCA)
        v0_810 <= v0_810 & ~maskExt_810 | maskExt_810 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hCA)
        v0_811 <= v0_811 & ~maskExt_811 | maskExt_811 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hCB)
        v0_812 <= v0_812 & ~maskExt_812 | maskExt_812 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hCB)
        v0_813 <= v0_813 & ~maskExt_813 | maskExt_813 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hCB)
        v0_814 <= v0_814 & ~maskExt_814 | maskExt_814 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hCB)
        v0_815 <= v0_815 & ~maskExt_815 | maskExt_815 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hCC)
        v0_816 <= v0_816 & ~maskExt_816 | maskExt_816 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hCC)
        v0_817 <= v0_817 & ~maskExt_817 | maskExt_817 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hCC)
        v0_818 <= v0_818 & ~maskExt_818 | maskExt_818 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hCC)
        v0_819 <= v0_819 & ~maskExt_819 | maskExt_819 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hCD)
        v0_820 <= v0_820 & ~maskExt_820 | maskExt_820 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hCD)
        v0_821 <= v0_821 & ~maskExt_821 | maskExt_821 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hCD)
        v0_822 <= v0_822 & ~maskExt_822 | maskExt_822 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hCD)
        v0_823 <= v0_823 & ~maskExt_823 | maskExt_823 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hCE)
        v0_824 <= v0_824 & ~maskExt_824 | maskExt_824 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hCE)
        v0_825 <= v0_825 & ~maskExt_825 | maskExt_825 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hCE)
        v0_826 <= v0_826 & ~maskExt_826 | maskExt_826 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hCE)
        v0_827 <= v0_827 & ~maskExt_827 | maskExt_827 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hCF)
        v0_828 <= v0_828 & ~maskExt_828 | maskExt_828 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hCF)
        v0_829 <= v0_829 & ~maskExt_829 | maskExt_829 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hCF)
        v0_830 <= v0_830 & ~maskExt_830 | maskExt_830 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hCF)
        v0_831 <= v0_831 & ~maskExt_831 | maskExt_831 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hD0)
        v0_832 <= v0_832 & ~maskExt_832 | maskExt_832 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hD0)
        v0_833 <= v0_833 & ~maskExt_833 | maskExt_833 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hD0)
        v0_834 <= v0_834 & ~maskExt_834 | maskExt_834 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hD0)
        v0_835 <= v0_835 & ~maskExt_835 | maskExt_835 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hD1)
        v0_836 <= v0_836 & ~maskExt_836 | maskExt_836 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hD1)
        v0_837 <= v0_837 & ~maskExt_837 | maskExt_837 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hD1)
        v0_838 <= v0_838 & ~maskExt_838 | maskExt_838 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hD1)
        v0_839 <= v0_839 & ~maskExt_839 | maskExt_839 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hD2)
        v0_840 <= v0_840 & ~maskExt_840 | maskExt_840 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hD2)
        v0_841 <= v0_841 & ~maskExt_841 | maskExt_841 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hD2)
        v0_842 <= v0_842 & ~maskExt_842 | maskExt_842 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hD2)
        v0_843 <= v0_843 & ~maskExt_843 | maskExt_843 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hD3)
        v0_844 <= v0_844 & ~maskExt_844 | maskExt_844 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hD3)
        v0_845 <= v0_845 & ~maskExt_845 | maskExt_845 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hD3)
        v0_846 <= v0_846 & ~maskExt_846 | maskExt_846 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hD3)
        v0_847 <= v0_847 & ~maskExt_847 | maskExt_847 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hD4)
        v0_848 <= v0_848 & ~maskExt_848 | maskExt_848 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hD4)
        v0_849 <= v0_849 & ~maskExt_849 | maskExt_849 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hD4)
        v0_850 <= v0_850 & ~maskExt_850 | maskExt_850 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hD4)
        v0_851 <= v0_851 & ~maskExt_851 | maskExt_851 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hD5)
        v0_852 <= v0_852 & ~maskExt_852 | maskExt_852 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hD5)
        v0_853 <= v0_853 & ~maskExt_853 | maskExt_853 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hD5)
        v0_854 <= v0_854 & ~maskExt_854 | maskExt_854 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hD5)
        v0_855 <= v0_855 & ~maskExt_855 | maskExt_855 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hD6)
        v0_856 <= v0_856 & ~maskExt_856 | maskExt_856 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hD6)
        v0_857 <= v0_857 & ~maskExt_857 | maskExt_857 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hD6)
        v0_858 <= v0_858 & ~maskExt_858 | maskExt_858 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hD6)
        v0_859 <= v0_859 & ~maskExt_859 | maskExt_859 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hD7)
        v0_860 <= v0_860 & ~maskExt_860 | maskExt_860 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hD7)
        v0_861 <= v0_861 & ~maskExt_861 | maskExt_861 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hD7)
        v0_862 <= v0_862 & ~maskExt_862 | maskExt_862 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hD7)
        v0_863 <= v0_863 & ~maskExt_863 | maskExt_863 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hD8)
        v0_864 <= v0_864 & ~maskExt_864 | maskExt_864 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hD8)
        v0_865 <= v0_865 & ~maskExt_865 | maskExt_865 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hD8)
        v0_866 <= v0_866 & ~maskExt_866 | maskExt_866 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hD8)
        v0_867 <= v0_867 & ~maskExt_867 | maskExt_867 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hD9)
        v0_868 <= v0_868 & ~maskExt_868 | maskExt_868 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hD9)
        v0_869 <= v0_869 & ~maskExt_869 | maskExt_869 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hD9)
        v0_870 <= v0_870 & ~maskExt_870 | maskExt_870 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hD9)
        v0_871 <= v0_871 & ~maskExt_871 | maskExt_871 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hDA)
        v0_872 <= v0_872 & ~maskExt_872 | maskExt_872 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hDA)
        v0_873 <= v0_873 & ~maskExt_873 | maskExt_873 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hDA)
        v0_874 <= v0_874 & ~maskExt_874 | maskExt_874 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hDA)
        v0_875 <= v0_875 & ~maskExt_875 | maskExt_875 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hDB)
        v0_876 <= v0_876 & ~maskExt_876 | maskExt_876 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hDB)
        v0_877 <= v0_877 & ~maskExt_877 | maskExt_877 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hDB)
        v0_878 <= v0_878 & ~maskExt_878 | maskExt_878 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hDB)
        v0_879 <= v0_879 & ~maskExt_879 | maskExt_879 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hDC)
        v0_880 <= v0_880 & ~maskExt_880 | maskExt_880 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hDC)
        v0_881 <= v0_881 & ~maskExt_881 | maskExt_881 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hDC)
        v0_882 <= v0_882 & ~maskExt_882 | maskExt_882 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hDC)
        v0_883 <= v0_883 & ~maskExt_883 | maskExt_883 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hDD)
        v0_884 <= v0_884 & ~maskExt_884 | maskExt_884 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hDD)
        v0_885 <= v0_885 & ~maskExt_885 | maskExt_885 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hDD)
        v0_886 <= v0_886 & ~maskExt_886 | maskExt_886 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hDD)
        v0_887 <= v0_887 & ~maskExt_887 | maskExt_887 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hDE)
        v0_888 <= v0_888 & ~maskExt_888 | maskExt_888 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hDE)
        v0_889 <= v0_889 & ~maskExt_889 | maskExt_889 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hDE)
        v0_890 <= v0_890 & ~maskExt_890 | maskExt_890 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hDE)
        v0_891 <= v0_891 & ~maskExt_891 | maskExt_891 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hDF)
        v0_892 <= v0_892 & ~maskExt_892 | maskExt_892 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hDF)
        v0_893 <= v0_893 & ~maskExt_893 | maskExt_893 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hDF)
        v0_894 <= v0_894 & ~maskExt_894 | maskExt_894 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hDF)
        v0_895 <= v0_895 & ~maskExt_895 | maskExt_895 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hE0)
        v0_896 <= v0_896 & ~maskExt_896 | maskExt_896 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hE0)
        v0_897 <= v0_897 & ~maskExt_897 | maskExt_897 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hE0)
        v0_898 <= v0_898 & ~maskExt_898 | maskExt_898 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hE0)
        v0_899 <= v0_899 & ~maskExt_899 | maskExt_899 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hE1)
        v0_900 <= v0_900 & ~maskExt_900 | maskExt_900 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hE1)
        v0_901 <= v0_901 & ~maskExt_901 | maskExt_901 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hE1)
        v0_902 <= v0_902 & ~maskExt_902 | maskExt_902 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hE1)
        v0_903 <= v0_903 & ~maskExt_903 | maskExt_903 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hE2)
        v0_904 <= v0_904 & ~maskExt_904 | maskExt_904 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hE2)
        v0_905 <= v0_905 & ~maskExt_905 | maskExt_905 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hE2)
        v0_906 <= v0_906 & ~maskExt_906 | maskExt_906 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hE2)
        v0_907 <= v0_907 & ~maskExt_907 | maskExt_907 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hE3)
        v0_908 <= v0_908 & ~maskExt_908 | maskExt_908 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hE3)
        v0_909 <= v0_909 & ~maskExt_909 | maskExt_909 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hE3)
        v0_910 <= v0_910 & ~maskExt_910 | maskExt_910 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hE3)
        v0_911 <= v0_911 & ~maskExt_911 | maskExt_911 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hE4)
        v0_912 <= v0_912 & ~maskExt_912 | maskExt_912 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hE4)
        v0_913 <= v0_913 & ~maskExt_913 | maskExt_913 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hE4)
        v0_914 <= v0_914 & ~maskExt_914 | maskExt_914 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hE4)
        v0_915 <= v0_915 & ~maskExt_915 | maskExt_915 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hE5)
        v0_916 <= v0_916 & ~maskExt_916 | maskExt_916 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hE5)
        v0_917 <= v0_917 & ~maskExt_917 | maskExt_917 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hE5)
        v0_918 <= v0_918 & ~maskExt_918 | maskExt_918 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hE5)
        v0_919 <= v0_919 & ~maskExt_919 | maskExt_919 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hE6)
        v0_920 <= v0_920 & ~maskExt_920 | maskExt_920 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hE6)
        v0_921 <= v0_921 & ~maskExt_921 | maskExt_921 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hE6)
        v0_922 <= v0_922 & ~maskExt_922 | maskExt_922 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hE6)
        v0_923 <= v0_923 & ~maskExt_923 | maskExt_923 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hE7)
        v0_924 <= v0_924 & ~maskExt_924 | maskExt_924 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hE7)
        v0_925 <= v0_925 & ~maskExt_925 | maskExt_925 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hE7)
        v0_926 <= v0_926 & ~maskExt_926 | maskExt_926 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hE7)
        v0_927 <= v0_927 & ~maskExt_927 | maskExt_927 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hE8)
        v0_928 <= v0_928 & ~maskExt_928 | maskExt_928 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hE8)
        v0_929 <= v0_929 & ~maskExt_929 | maskExt_929 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hE8)
        v0_930 <= v0_930 & ~maskExt_930 | maskExt_930 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hE8)
        v0_931 <= v0_931 & ~maskExt_931 | maskExt_931 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hE9)
        v0_932 <= v0_932 & ~maskExt_932 | maskExt_932 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hE9)
        v0_933 <= v0_933 & ~maskExt_933 | maskExt_933 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hE9)
        v0_934 <= v0_934 & ~maskExt_934 | maskExt_934 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hE9)
        v0_935 <= v0_935 & ~maskExt_935 | maskExt_935 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hEA)
        v0_936 <= v0_936 & ~maskExt_936 | maskExt_936 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hEA)
        v0_937 <= v0_937 & ~maskExt_937 | maskExt_937 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hEA)
        v0_938 <= v0_938 & ~maskExt_938 | maskExt_938 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hEA)
        v0_939 <= v0_939 & ~maskExt_939 | maskExt_939 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hEB)
        v0_940 <= v0_940 & ~maskExt_940 | maskExt_940 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hEB)
        v0_941 <= v0_941 & ~maskExt_941 | maskExt_941 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hEB)
        v0_942 <= v0_942 & ~maskExt_942 | maskExt_942 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hEB)
        v0_943 <= v0_943 & ~maskExt_943 | maskExt_943 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hEC)
        v0_944 <= v0_944 & ~maskExt_944 | maskExt_944 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hEC)
        v0_945 <= v0_945 & ~maskExt_945 | maskExt_945 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hEC)
        v0_946 <= v0_946 & ~maskExt_946 | maskExt_946 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hEC)
        v0_947 <= v0_947 & ~maskExt_947 | maskExt_947 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hED)
        v0_948 <= v0_948 & ~maskExt_948 | maskExt_948 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hED)
        v0_949 <= v0_949 & ~maskExt_949 | maskExt_949 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hED)
        v0_950 <= v0_950 & ~maskExt_950 | maskExt_950 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hED)
        v0_951 <= v0_951 & ~maskExt_951 | maskExt_951 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hEE)
        v0_952 <= v0_952 & ~maskExt_952 | maskExt_952 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hEE)
        v0_953 <= v0_953 & ~maskExt_953 | maskExt_953 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hEE)
        v0_954 <= v0_954 & ~maskExt_954 | maskExt_954 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hEE)
        v0_955 <= v0_955 & ~maskExt_955 | maskExt_955 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hEF)
        v0_956 <= v0_956 & ~maskExt_956 | maskExt_956 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hEF)
        v0_957 <= v0_957 & ~maskExt_957 | maskExt_957 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hEF)
        v0_958 <= v0_958 & ~maskExt_958 | maskExt_958 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hEF)
        v0_959 <= v0_959 & ~maskExt_959 | maskExt_959 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hF0)
        v0_960 <= v0_960 & ~maskExt_960 | maskExt_960 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hF0)
        v0_961 <= v0_961 & ~maskExt_961 | maskExt_961 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hF0)
        v0_962 <= v0_962 & ~maskExt_962 | maskExt_962 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hF0)
        v0_963 <= v0_963 & ~maskExt_963 | maskExt_963 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hF1)
        v0_964 <= v0_964 & ~maskExt_964 | maskExt_964 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hF1)
        v0_965 <= v0_965 & ~maskExt_965 | maskExt_965 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hF1)
        v0_966 <= v0_966 & ~maskExt_966 | maskExt_966 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hF1)
        v0_967 <= v0_967 & ~maskExt_967 | maskExt_967 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hF2)
        v0_968 <= v0_968 & ~maskExt_968 | maskExt_968 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hF2)
        v0_969 <= v0_969 & ~maskExt_969 | maskExt_969 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hF2)
        v0_970 <= v0_970 & ~maskExt_970 | maskExt_970 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hF2)
        v0_971 <= v0_971 & ~maskExt_971 | maskExt_971 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hF3)
        v0_972 <= v0_972 & ~maskExt_972 | maskExt_972 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hF3)
        v0_973 <= v0_973 & ~maskExt_973 | maskExt_973 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hF3)
        v0_974 <= v0_974 & ~maskExt_974 | maskExt_974 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hF3)
        v0_975 <= v0_975 & ~maskExt_975 | maskExt_975 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hF4)
        v0_976 <= v0_976 & ~maskExt_976 | maskExt_976 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hF4)
        v0_977 <= v0_977 & ~maskExt_977 | maskExt_977 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hF4)
        v0_978 <= v0_978 & ~maskExt_978 | maskExt_978 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hF4)
        v0_979 <= v0_979 & ~maskExt_979 | maskExt_979 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hF5)
        v0_980 <= v0_980 & ~maskExt_980 | maskExt_980 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hF5)
        v0_981 <= v0_981 & ~maskExt_981 | maskExt_981 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hF5)
        v0_982 <= v0_982 & ~maskExt_982 | maskExt_982 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hF5)
        v0_983 <= v0_983 & ~maskExt_983 | maskExt_983 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hF6)
        v0_984 <= v0_984 & ~maskExt_984 | maskExt_984 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hF6)
        v0_985 <= v0_985 & ~maskExt_985 | maskExt_985 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hF6)
        v0_986 <= v0_986 & ~maskExt_986 | maskExt_986 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hF6)
        v0_987 <= v0_987 & ~maskExt_987 | maskExt_987 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hF7)
        v0_988 <= v0_988 & ~maskExt_988 | maskExt_988 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hF7)
        v0_989 <= v0_989 & ~maskExt_989 | maskExt_989 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hF7)
        v0_990 <= v0_990 & ~maskExt_990 | maskExt_990 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hF7)
        v0_991 <= v0_991 & ~maskExt_991 | maskExt_991 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hF8)
        v0_992 <= v0_992 & ~maskExt_992 | maskExt_992 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hF8)
        v0_993 <= v0_993 & ~maskExt_993 | maskExt_993 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hF8)
        v0_994 <= v0_994 & ~maskExt_994 | maskExt_994 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hF8)
        v0_995 <= v0_995 & ~maskExt_995 | maskExt_995 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hF9)
        v0_996 <= v0_996 & ~maskExt_996 | maskExt_996 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hF9)
        v0_997 <= v0_997 & ~maskExt_997 | maskExt_997 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hF9)
        v0_998 <= v0_998 & ~maskExt_998 | maskExt_998 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hF9)
        v0_999 <= v0_999 & ~maskExt_999 | maskExt_999 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hFA)
        v0_1000 <= v0_1000 & ~maskExt_1000 | maskExt_1000 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hFA)
        v0_1001 <= v0_1001 & ~maskExt_1001 | maskExt_1001 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hFA)
        v0_1002 <= v0_1002 & ~maskExt_1002 | maskExt_1002 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hFA)
        v0_1003 <= v0_1003 & ~maskExt_1003 | maskExt_1003 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hFB)
        v0_1004 <= v0_1004 & ~maskExt_1004 | maskExt_1004 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hFB)
        v0_1005 <= v0_1005 & ~maskExt_1005 | maskExt_1005 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hFB)
        v0_1006 <= v0_1006 & ~maskExt_1006 | maskExt_1006 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hFB)
        v0_1007 <= v0_1007 & ~maskExt_1007 | maskExt_1007 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hFC)
        v0_1008 <= v0_1008 & ~maskExt_1008 | maskExt_1008 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hFC)
        v0_1009 <= v0_1009 & ~maskExt_1009 | maskExt_1009 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hFC)
        v0_1010 <= v0_1010 & ~maskExt_1010 | maskExt_1010 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hFC)
        v0_1011 <= v0_1011 & ~maskExt_1011 | maskExt_1011 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hFD)
        v0_1012 <= v0_1012 & ~maskExt_1012 | maskExt_1012 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hFD)
        v0_1013 <= v0_1013 & ~maskExt_1013 | maskExt_1013 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hFD)
        v0_1014 <= v0_1014 & ~maskExt_1014 | maskExt_1014 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hFD)
        v0_1015 <= v0_1015 & ~maskExt_1015 | maskExt_1015 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hFE)
        v0_1016 <= v0_1016 & ~maskExt_1016 | maskExt_1016 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hFE)
        v0_1017 <= v0_1017 & ~maskExt_1017 | maskExt_1017 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hFE)
        v0_1018 <= v0_1018 & ~maskExt_1018 | maskExt_1018 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hFE)
        v0_1019 <= v0_1019 & ~maskExt_1019 | maskExt_1019 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'hFF)
        v0_1020 <= v0_1020 & ~maskExt_1020 | maskExt_1020 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'hFF)
        v0_1021 <= v0_1021 & ~maskExt_1021 | maskExt_1021 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'hFF)
        v0_1022 <= v0_1022 & ~maskExt_1022 | maskExt_1022 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'hFF)
        v0_1023 <= v0_1023 & ~maskExt_1023 | maskExt_1023 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h100)
        v0_1024 <= v0_1024 & ~maskExt_1024 | maskExt_1024 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h100)
        v0_1025 <= v0_1025 & ~maskExt_1025 | maskExt_1025 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h100)
        v0_1026 <= v0_1026 & ~maskExt_1026 | maskExt_1026 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h100)
        v0_1027 <= v0_1027 & ~maskExt_1027 | maskExt_1027 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h101)
        v0_1028 <= v0_1028 & ~maskExt_1028 | maskExt_1028 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h101)
        v0_1029 <= v0_1029 & ~maskExt_1029 | maskExt_1029 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h101)
        v0_1030 <= v0_1030 & ~maskExt_1030 | maskExt_1030 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h101)
        v0_1031 <= v0_1031 & ~maskExt_1031 | maskExt_1031 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h102)
        v0_1032 <= v0_1032 & ~maskExt_1032 | maskExt_1032 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h102)
        v0_1033 <= v0_1033 & ~maskExt_1033 | maskExt_1033 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h102)
        v0_1034 <= v0_1034 & ~maskExt_1034 | maskExt_1034 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h102)
        v0_1035 <= v0_1035 & ~maskExt_1035 | maskExt_1035 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h103)
        v0_1036 <= v0_1036 & ~maskExt_1036 | maskExt_1036 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h103)
        v0_1037 <= v0_1037 & ~maskExt_1037 | maskExt_1037 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h103)
        v0_1038 <= v0_1038 & ~maskExt_1038 | maskExt_1038 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h103)
        v0_1039 <= v0_1039 & ~maskExt_1039 | maskExt_1039 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h104)
        v0_1040 <= v0_1040 & ~maskExt_1040 | maskExt_1040 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h104)
        v0_1041 <= v0_1041 & ~maskExt_1041 | maskExt_1041 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h104)
        v0_1042 <= v0_1042 & ~maskExt_1042 | maskExt_1042 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h104)
        v0_1043 <= v0_1043 & ~maskExt_1043 | maskExt_1043 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h105)
        v0_1044 <= v0_1044 & ~maskExt_1044 | maskExt_1044 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h105)
        v0_1045 <= v0_1045 & ~maskExt_1045 | maskExt_1045 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h105)
        v0_1046 <= v0_1046 & ~maskExt_1046 | maskExt_1046 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h105)
        v0_1047 <= v0_1047 & ~maskExt_1047 | maskExt_1047 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h106)
        v0_1048 <= v0_1048 & ~maskExt_1048 | maskExt_1048 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h106)
        v0_1049 <= v0_1049 & ~maskExt_1049 | maskExt_1049 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h106)
        v0_1050 <= v0_1050 & ~maskExt_1050 | maskExt_1050 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h106)
        v0_1051 <= v0_1051 & ~maskExt_1051 | maskExt_1051 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h107)
        v0_1052 <= v0_1052 & ~maskExt_1052 | maskExt_1052 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h107)
        v0_1053 <= v0_1053 & ~maskExt_1053 | maskExt_1053 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h107)
        v0_1054 <= v0_1054 & ~maskExt_1054 | maskExt_1054 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h107)
        v0_1055 <= v0_1055 & ~maskExt_1055 | maskExt_1055 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h108)
        v0_1056 <= v0_1056 & ~maskExt_1056 | maskExt_1056 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h108)
        v0_1057 <= v0_1057 & ~maskExt_1057 | maskExt_1057 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h108)
        v0_1058 <= v0_1058 & ~maskExt_1058 | maskExt_1058 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h108)
        v0_1059 <= v0_1059 & ~maskExt_1059 | maskExt_1059 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h109)
        v0_1060 <= v0_1060 & ~maskExt_1060 | maskExt_1060 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h109)
        v0_1061 <= v0_1061 & ~maskExt_1061 | maskExt_1061 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h109)
        v0_1062 <= v0_1062 & ~maskExt_1062 | maskExt_1062 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h109)
        v0_1063 <= v0_1063 & ~maskExt_1063 | maskExt_1063 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h10A)
        v0_1064 <= v0_1064 & ~maskExt_1064 | maskExt_1064 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h10A)
        v0_1065 <= v0_1065 & ~maskExt_1065 | maskExt_1065 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h10A)
        v0_1066 <= v0_1066 & ~maskExt_1066 | maskExt_1066 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h10A)
        v0_1067 <= v0_1067 & ~maskExt_1067 | maskExt_1067 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h10B)
        v0_1068 <= v0_1068 & ~maskExt_1068 | maskExt_1068 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h10B)
        v0_1069 <= v0_1069 & ~maskExt_1069 | maskExt_1069 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h10B)
        v0_1070 <= v0_1070 & ~maskExt_1070 | maskExt_1070 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h10B)
        v0_1071 <= v0_1071 & ~maskExt_1071 | maskExt_1071 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h10C)
        v0_1072 <= v0_1072 & ~maskExt_1072 | maskExt_1072 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h10C)
        v0_1073 <= v0_1073 & ~maskExt_1073 | maskExt_1073 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h10C)
        v0_1074 <= v0_1074 & ~maskExt_1074 | maskExt_1074 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h10C)
        v0_1075 <= v0_1075 & ~maskExt_1075 | maskExt_1075 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h10D)
        v0_1076 <= v0_1076 & ~maskExt_1076 | maskExt_1076 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h10D)
        v0_1077 <= v0_1077 & ~maskExt_1077 | maskExt_1077 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h10D)
        v0_1078 <= v0_1078 & ~maskExt_1078 | maskExt_1078 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h10D)
        v0_1079 <= v0_1079 & ~maskExt_1079 | maskExt_1079 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h10E)
        v0_1080 <= v0_1080 & ~maskExt_1080 | maskExt_1080 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h10E)
        v0_1081 <= v0_1081 & ~maskExt_1081 | maskExt_1081 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h10E)
        v0_1082 <= v0_1082 & ~maskExt_1082 | maskExt_1082 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h10E)
        v0_1083 <= v0_1083 & ~maskExt_1083 | maskExt_1083 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h10F)
        v0_1084 <= v0_1084 & ~maskExt_1084 | maskExt_1084 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h10F)
        v0_1085 <= v0_1085 & ~maskExt_1085 | maskExt_1085 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h10F)
        v0_1086 <= v0_1086 & ~maskExt_1086 | maskExt_1086 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h10F)
        v0_1087 <= v0_1087 & ~maskExt_1087 | maskExt_1087 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h110)
        v0_1088 <= v0_1088 & ~maskExt_1088 | maskExt_1088 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h110)
        v0_1089 <= v0_1089 & ~maskExt_1089 | maskExt_1089 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h110)
        v0_1090 <= v0_1090 & ~maskExt_1090 | maskExt_1090 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h110)
        v0_1091 <= v0_1091 & ~maskExt_1091 | maskExt_1091 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h111)
        v0_1092 <= v0_1092 & ~maskExt_1092 | maskExt_1092 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h111)
        v0_1093 <= v0_1093 & ~maskExt_1093 | maskExt_1093 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h111)
        v0_1094 <= v0_1094 & ~maskExt_1094 | maskExt_1094 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h111)
        v0_1095 <= v0_1095 & ~maskExt_1095 | maskExt_1095 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h112)
        v0_1096 <= v0_1096 & ~maskExt_1096 | maskExt_1096 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h112)
        v0_1097 <= v0_1097 & ~maskExt_1097 | maskExt_1097 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h112)
        v0_1098 <= v0_1098 & ~maskExt_1098 | maskExt_1098 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h112)
        v0_1099 <= v0_1099 & ~maskExt_1099 | maskExt_1099 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h113)
        v0_1100 <= v0_1100 & ~maskExt_1100 | maskExt_1100 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h113)
        v0_1101 <= v0_1101 & ~maskExt_1101 | maskExt_1101 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h113)
        v0_1102 <= v0_1102 & ~maskExt_1102 | maskExt_1102 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h113)
        v0_1103 <= v0_1103 & ~maskExt_1103 | maskExt_1103 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h114)
        v0_1104 <= v0_1104 & ~maskExt_1104 | maskExt_1104 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h114)
        v0_1105 <= v0_1105 & ~maskExt_1105 | maskExt_1105 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h114)
        v0_1106 <= v0_1106 & ~maskExt_1106 | maskExt_1106 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h114)
        v0_1107 <= v0_1107 & ~maskExt_1107 | maskExt_1107 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h115)
        v0_1108 <= v0_1108 & ~maskExt_1108 | maskExt_1108 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h115)
        v0_1109 <= v0_1109 & ~maskExt_1109 | maskExt_1109 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h115)
        v0_1110 <= v0_1110 & ~maskExt_1110 | maskExt_1110 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h115)
        v0_1111 <= v0_1111 & ~maskExt_1111 | maskExt_1111 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h116)
        v0_1112 <= v0_1112 & ~maskExt_1112 | maskExt_1112 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h116)
        v0_1113 <= v0_1113 & ~maskExt_1113 | maskExt_1113 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h116)
        v0_1114 <= v0_1114 & ~maskExt_1114 | maskExt_1114 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h116)
        v0_1115 <= v0_1115 & ~maskExt_1115 | maskExt_1115 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h117)
        v0_1116 <= v0_1116 & ~maskExt_1116 | maskExt_1116 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h117)
        v0_1117 <= v0_1117 & ~maskExt_1117 | maskExt_1117 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h117)
        v0_1118 <= v0_1118 & ~maskExt_1118 | maskExt_1118 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h117)
        v0_1119 <= v0_1119 & ~maskExt_1119 | maskExt_1119 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h118)
        v0_1120 <= v0_1120 & ~maskExt_1120 | maskExt_1120 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h118)
        v0_1121 <= v0_1121 & ~maskExt_1121 | maskExt_1121 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h118)
        v0_1122 <= v0_1122 & ~maskExt_1122 | maskExt_1122 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h118)
        v0_1123 <= v0_1123 & ~maskExt_1123 | maskExt_1123 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h119)
        v0_1124 <= v0_1124 & ~maskExt_1124 | maskExt_1124 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h119)
        v0_1125 <= v0_1125 & ~maskExt_1125 | maskExt_1125 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h119)
        v0_1126 <= v0_1126 & ~maskExt_1126 | maskExt_1126 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h119)
        v0_1127 <= v0_1127 & ~maskExt_1127 | maskExt_1127 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h11A)
        v0_1128 <= v0_1128 & ~maskExt_1128 | maskExt_1128 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h11A)
        v0_1129 <= v0_1129 & ~maskExt_1129 | maskExt_1129 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h11A)
        v0_1130 <= v0_1130 & ~maskExt_1130 | maskExt_1130 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h11A)
        v0_1131 <= v0_1131 & ~maskExt_1131 | maskExt_1131 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h11B)
        v0_1132 <= v0_1132 & ~maskExt_1132 | maskExt_1132 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h11B)
        v0_1133 <= v0_1133 & ~maskExt_1133 | maskExt_1133 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h11B)
        v0_1134 <= v0_1134 & ~maskExt_1134 | maskExt_1134 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h11B)
        v0_1135 <= v0_1135 & ~maskExt_1135 | maskExt_1135 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h11C)
        v0_1136 <= v0_1136 & ~maskExt_1136 | maskExt_1136 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h11C)
        v0_1137 <= v0_1137 & ~maskExt_1137 | maskExt_1137 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h11C)
        v0_1138 <= v0_1138 & ~maskExt_1138 | maskExt_1138 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h11C)
        v0_1139 <= v0_1139 & ~maskExt_1139 | maskExt_1139 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h11D)
        v0_1140 <= v0_1140 & ~maskExt_1140 | maskExt_1140 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h11D)
        v0_1141 <= v0_1141 & ~maskExt_1141 | maskExt_1141 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h11D)
        v0_1142 <= v0_1142 & ~maskExt_1142 | maskExt_1142 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h11D)
        v0_1143 <= v0_1143 & ~maskExt_1143 | maskExt_1143 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h11E)
        v0_1144 <= v0_1144 & ~maskExt_1144 | maskExt_1144 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h11E)
        v0_1145 <= v0_1145 & ~maskExt_1145 | maskExt_1145 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h11E)
        v0_1146 <= v0_1146 & ~maskExt_1146 | maskExt_1146 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h11E)
        v0_1147 <= v0_1147 & ~maskExt_1147 | maskExt_1147 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h11F)
        v0_1148 <= v0_1148 & ~maskExt_1148 | maskExt_1148 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h11F)
        v0_1149 <= v0_1149 & ~maskExt_1149 | maskExt_1149 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h11F)
        v0_1150 <= v0_1150 & ~maskExt_1150 | maskExt_1150 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h11F)
        v0_1151 <= v0_1151 & ~maskExt_1151 | maskExt_1151 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h120)
        v0_1152 <= v0_1152 & ~maskExt_1152 | maskExt_1152 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h120)
        v0_1153 <= v0_1153 & ~maskExt_1153 | maskExt_1153 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h120)
        v0_1154 <= v0_1154 & ~maskExt_1154 | maskExt_1154 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h120)
        v0_1155 <= v0_1155 & ~maskExt_1155 | maskExt_1155 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h121)
        v0_1156 <= v0_1156 & ~maskExt_1156 | maskExt_1156 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h121)
        v0_1157 <= v0_1157 & ~maskExt_1157 | maskExt_1157 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h121)
        v0_1158 <= v0_1158 & ~maskExt_1158 | maskExt_1158 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h121)
        v0_1159 <= v0_1159 & ~maskExt_1159 | maskExt_1159 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h122)
        v0_1160 <= v0_1160 & ~maskExt_1160 | maskExt_1160 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h122)
        v0_1161 <= v0_1161 & ~maskExt_1161 | maskExt_1161 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h122)
        v0_1162 <= v0_1162 & ~maskExt_1162 | maskExt_1162 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h122)
        v0_1163 <= v0_1163 & ~maskExt_1163 | maskExt_1163 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h123)
        v0_1164 <= v0_1164 & ~maskExt_1164 | maskExt_1164 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h123)
        v0_1165 <= v0_1165 & ~maskExt_1165 | maskExt_1165 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h123)
        v0_1166 <= v0_1166 & ~maskExt_1166 | maskExt_1166 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h123)
        v0_1167 <= v0_1167 & ~maskExt_1167 | maskExt_1167 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h124)
        v0_1168 <= v0_1168 & ~maskExt_1168 | maskExt_1168 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h124)
        v0_1169 <= v0_1169 & ~maskExt_1169 | maskExt_1169 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h124)
        v0_1170 <= v0_1170 & ~maskExt_1170 | maskExt_1170 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h124)
        v0_1171 <= v0_1171 & ~maskExt_1171 | maskExt_1171 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h125)
        v0_1172 <= v0_1172 & ~maskExt_1172 | maskExt_1172 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h125)
        v0_1173 <= v0_1173 & ~maskExt_1173 | maskExt_1173 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h125)
        v0_1174 <= v0_1174 & ~maskExt_1174 | maskExt_1174 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h125)
        v0_1175 <= v0_1175 & ~maskExt_1175 | maskExt_1175 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h126)
        v0_1176 <= v0_1176 & ~maskExt_1176 | maskExt_1176 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h126)
        v0_1177 <= v0_1177 & ~maskExt_1177 | maskExt_1177 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h126)
        v0_1178 <= v0_1178 & ~maskExt_1178 | maskExt_1178 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h126)
        v0_1179 <= v0_1179 & ~maskExt_1179 | maskExt_1179 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h127)
        v0_1180 <= v0_1180 & ~maskExt_1180 | maskExt_1180 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h127)
        v0_1181 <= v0_1181 & ~maskExt_1181 | maskExt_1181 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h127)
        v0_1182 <= v0_1182 & ~maskExt_1182 | maskExt_1182 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h127)
        v0_1183 <= v0_1183 & ~maskExt_1183 | maskExt_1183 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h128)
        v0_1184 <= v0_1184 & ~maskExt_1184 | maskExt_1184 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h128)
        v0_1185 <= v0_1185 & ~maskExt_1185 | maskExt_1185 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h128)
        v0_1186 <= v0_1186 & ~maskExt_1186 | maskExt_1186 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h128)
        v0_1187 <= v0_1187 & ~maskExt_1187 | maskExt_1187 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h129)
        v0_1188 <= v0_1188 & ~maskExt_1188 | maskExt_1188 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h129)
        v0_1189 <= v0_1189 & ~maskExt_1189 | maskExt_1189 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h129)
        v0_1190 <= v0_1190 & ~maskExt_1190 | maskExt_1190 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h129)
        v0_1191 <= v0_1191 & ~maskExt_1191 | maskExt_1191 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h12A)
        v0_1192 <= v0_1192 & ~maskExt_1192 | maskExt_1192 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h12A)
        v0_1193 <= v0_1193 & ~maskExt_1193 | maskExt_1193 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h12A)
        v0_1194 <= v0_1194 & ~maskExt_1194 | maskExt_1194 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h12A)
        v0_1195 <= v0_1195 & ~maskExt_1195 | maskExt_1195 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h12B)
        v0_1196 <= v0_1196 & ~maskExt_1196 | maskExt_1196 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h12B)
        v0_1197 <= v0_1197 & ~maskExt_1197 | maskExt_1197 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h12B)
        v0_1198 <= v0_1198 & ~maskExt_1198 | maskExt_1198 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h12B)
        v0_1199 <= v0_1199 & ~maskExt_1199 | maskExt_1199 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h12C)
        v0_1200 <= v0_1200 & ~maskExt_1200 | maskExt_1200 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h12C)
        v0_1201 <= v0_1201 & ~maskExt_1201 | maskExt_1201 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h12C)
        v0_1202 <= v0_1202 & ~maskExt_1202 | maskExt_1202 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h12C)
        v0_1203 <= v0_1203 & ~maskExt_1203 | maskExt_1203 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h12D)
        v0_1204 <= v0_1204 & ~maskExt_1204 | maskExt_1204 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h12D)
        v0_1205 <= v0_1205 & ~maskExt_1205 | maskExt_1205 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h12D)
        v0_1206 <= v0_1206 & ~maskExt_1206 | maskExt_1206 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h12D)
        v0_1207 <= v0_1207 & ~maskExt_1207 | maskExt_1207 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h12E)
        v0_1208 <= v0_1208 & ~maskExt_1208 | maskExt_1208 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h12E)
        v0_1209 <= v0_1209 & ~maskExt_1209 | maskExt_1209 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h12E)
        v0_1210 <= v0_1210 & ~maskExt_1210 | maskExt_1210 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h12E)
        v0_1211 <= v0_1211 & ~maskExt_1211 | maskExt_1211 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h12F)
        v0_1212 <= v0_1212 & ~maskExt_1212 | maskExt_1212 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h12F)
        v0_1213 <= v0_1213 & ~maskExt_1213 | maskExt_1213 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h12F)
        v0_1214 <= v0_1214 & ~maskExt_1214 | maskExt_1214 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h12F)
        v0_1215 <= v0_1215 & ~maskExt_1215 | maskExt_1215 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h130)
        v0_1216 <= v0_1216 & ~maskExt_1216 | maskExt_1216 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h130)
        v0_1217 <= v0_1217 & ~maskExt_1217 | maskExt_1217 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h130)
        v0_1218 <= v0_1218 & ~maskExt_1218 | maskExt_1218 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h130)
        v0_1219 <= v0_1219 & ~maskExt_1219 | maskExt_1219 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h131)
        v0_1220 <= v0_1220 & ~maskExt_1220 | maskExt_1220 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h131)
        v0_1221 <= v0_1221 & ~maskExt_1221 | maskExt_1221 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h131)
        v0_1222 <= v0_1222 & ~maskExt_1222 | maskExt_1222 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h131)
        v0_1223 <= v0_1223 & ~maskExt_1223 | maskExt_1223 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h132)
        v0_1224 <= v0_1224 & ~maskExt_1224 | maskExt_1224 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h132)
        v0_1225 <= v0_1225 & ~maskExt_1225 | maskExt_1225 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h132)
        v0_1226 <= v0_1226 & ~maskExt_1226 | maskExt_1226 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h132)
        v0_1227 <= v0_1227 & ~maskExt_1227 | maskExt_1227 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h133)
        v0_1228 <= v0_1228 & ~maskExt_1228 | maskExt_1228 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h133)
        v0_1229 <= v0_1229 & ~maskExt_1229 | maskExt_1229 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h133)
        v0_1230 <= v0_1230 & ~maskExt_1230 | maskExt_1230 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h133)
        v0_1231 <= v0_1231 & ~maskExt_1231 | maskExt_1231 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h134)
        v0_1232 <= v0_1232 & ~maskExt_1232 | maskExt_1232 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h134)
        v0_1233 <= v0_1233 & ~maskExt_1233 | maskExt_1233 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h134)
        v0_1234 <= v0_1234 & ~maskExt_1234 | maskExt_1234 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h134)
        v0_1235 <= v0_1235 & ~maskExt_1235 | maskExt_1235 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h135)
        v0_1236 <= v0_1236 & ~maskExt_1236 | maskExt_1236 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h135)
        v0_1237 <= v0_1237 & ~maskExt_1237 | maskExt_1237 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h135)
        v0_1238 <= v0_1238 & ~maskExt_1238 | maskExt_1238 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h135)
        v0_1239 <= v0_1239 & ~maskExt_1239 | maskExt_1239 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h136)
        v0_1240 <= v0_1240 & ~maskExt_1240 | maskExt_1240 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h136)
        v0_1241 <= v0_1241 & ~maskExt_1241 | maskExt_1241 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h136)
        v0_1242 <= v0_1242 & ~maskExt_1242 | maskExt_1242 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h136)
        v0_1243 <= v0_1243 & ~maskExt_1243 | maskExt_1243 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h137)
        v0_1244 <= v0_1244 & ~maskExt_1244 | maskExt_1244 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h137)
        v0_1245 <= v0_1245 & ~maskExt_1245 | maskExt_1245 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h137)
        v0_1246 <= v0_1246 & ~maskExt_1246 | maskExt_1246 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h137)
        v0_1247 <= v0_1247 & ~maskExt_1247 | maskExt_1247 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h138)
        v0_1248 <= v0_1248 & ~maskExt_1248 | maskExt_1248 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h138)
        v0_1249 <= v0_1249 & ~maskExt_1249 | maskExt_1249 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h138)
        v0_1250 <= v0_1250 & ~maskExt_1250 | maskExt_1250 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h138)
        v0_1251 <= v0_1251 & ~maskExt_1251 | maskExt_1251 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h139)
        v0_1252 <= v0_1252 & ~maskExt_1252 | maskExt_1252 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h139)
        v0_1253 <= v0_1253 & ~maskExt_1253 | maskExt_1253 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h139)
        v0_1254 <= v0_1254 & ~maskExt_1254 | maskExt_1254 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h139)
        v0_1255 <= v0_1255 & ~maskExt_1255 | maskExt_1255 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h13A)
        v0_1256 <= v0_1256 & ~maskExt_1256 | maskExt_1256 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h13A)
        v0_1257 <= v0_1257 & ~maskExt_1257 | maskExt_1257 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h13A)
        v0_1258 <= v0_1258 & ~maskExt_1258 | maskExt_1258 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h13A)
        v0_1259 <= v0_1259 & ~maskExt_1259 | maskExt_1259 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h13B)
        v0_1260 <= v0_1260 & ~maskExt_1260 | maskExt_1260 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h13B)
        v0_1261 <= v0_1261 & ~maskExt_1261 | maskExt_1261 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h13B)
        v0_1262 <= v0_1262 & ~maskExt_1262 | maskExt_1262 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h13B)
        v0_1263 <= v0_1263 & ~maskExt_1263 | maskExt_1263 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h13C)
        v0_1264 <= v0_1264 & ~maskExt_1264 | maskExt_1264 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h13C)
        v0_1265 <= v0_1265 & ~maskExt_1265 | maskExt_1265 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h13C)
        v0_1266 <= v0_1266 & ~maskExt_1266 | maskExt_1266 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h13C)
        v0_1267 <= v0_1267 & ~maskExt_1267 | maskExt_1267 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h13D)
        v0_1268 <= v0_1268 & ~maskExt_1268 | maskExt_1268 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h13D)
        v0_1269 <= v0_1269 & ~maskExt_1269 | maskExt_1269 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h13D)
        v0_1270 <= v0_1270 & ~maskExt_1270 | maskExt_1270 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h13D)
        v0_1271 <= v0_1271 & ~maskExt_1271 | maskExt_1271 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h13E)
        v0_1272 <= v0_1272 & ~maskExt_1272 | maskExt_1272 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h13E)
        v0_1273 <= v0_1273 & ~maskExt_1273 | maskExt_1273 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h13E)
        v0_1274 <= v0_1274 & ~maskExt_1274 | maskExt_1274 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h13E)
        v0_1275 <= v0_1275 & ~maskExt_1275 | maskExt_1275 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h13F)
        v0_1276 <= v0_1276 & ~maskExt_1276 | maskExt_1276 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h13F)
        v0_1277 <= v0_1277 & ~maskExt_1277 | maskExt_1277 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h13F)
        v0_1278 <= v0_1278 & ~maskExt_1278 | maskExt_1278 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h13F)
        v0_1279 <= v0_1279 & ~maskExt_1279 | maskExt_1279 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h140)
        v0_1280 <= v0_1280 & ~maskExt_1280 | maskExt_1280 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h140)
        v0_1281 <= v0_1281 & ~maskExt_1281 | maskExt_1281 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h140)
        v0_1282 <= v0_1282 & ~maskExt_1282 | maskExt_1282 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h140)
        v0_1283 <= v0_1283 & ~maskExt_1283 | maskExt_1283 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h141)
        v0_1284 <= v0_1284 & ~maskExt_1284 | maskExt_1284 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h141)
        v0_1285 <= v0_1285 & ~maskExt_1285 | maskExt_1285 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h141)
        v0_1286 <= v0_1286 & ~maskExt_1286 | maskExt_1286 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h141)
        v0_1287 <= v0_1287 & ~maskExt_1287 | maskExt_1287 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h142)
        v0_1288 <= v0_1288 & ~maskExt_1288 | maskExt_1288 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h142)
        v0_1289 <= v0_1289 & ~maskExt_1289 | maskExt_1289 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h142)
        v0_1290 <= v0_1290 & ~maskExt_1290 | maskExt_1290 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h142)
        v0_1291 <= v0_1291 & ~maskExt_1291 | maskExt_1291 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h143)
        v0_1292 <= v0_1292 & ~maskExt_1292 | maskExt_1292 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h143)
        v0_1293 <= v0_1293 & ~maskExt_1293 | maskExt_1293 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h143)
        v0_1294 <= v0_1294 & ~maskExt_1294 | maskExt_1294 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h143)
        v0_1295 <= v0_1295 & ~maskExt_1295 | maskExt_1295 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h144)
        v0_1296 <= v0_1296 & ~maskExt_1296 | maskExt_1296 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h144)
        v0_1297 <= v0_1297 & ~maskExt_1297 | maskExt_1297 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h144)
        v0_1298 <= v0_1298 & ~maskExt_1298 | maskExt_1298 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h144)
        v0_1299 <= v0_1299 & ~maskExt_1299 | maskExt_1299 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h145)
        v0_1300 <= v0_1300 & ~maskExt_1300 | maskExt_1300 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h145)
        v0_1301 <= v0_1301 & ~maskExt_1301 | maskExt_1301 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h145)
        v0_1302 <= v0_1302 & ~maskExt_1302 | maskExt_1302 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h145)
        v0_1303 <= v0_1303 & ~maskExt_1303 | maskExt_1303 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h146)
        v0_1304 <= v0_1304 & ~maskExt_1304 | maskExt_1304 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h146)
        v0_1305 <= v0_1305 & ~maskExt_1305 | maskExt_1305 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h146)
        v0_1306 <= v0_1306 & ~maskExt_1306 | maskExt_1306 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h146)
        v0_1307 <= v0_1307 & ~maskExt_1307 | maskExt_1307 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h147)
        v0_1308 <= v0_1308 & ~maskExt_1308 | maskExt_1308 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h147)
        v0_1309 <= v0_1309 & ~maskExt_1309 | maskExt_1309 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h147)
        v0_1310 <= v0_1310 & ~maskExt_1310 | maskExt_1310 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h147)
        v0_1311 <= v0_1311 & ~maskExt_1311 | maskExt_1311 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h148)
        v0_1312 <= v0_1312 & ~maskExt_1312 | maskExt_1312 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h148)
        v0_1313 <= v0_1313 & ~maskExt_1313 | maskExt_1313 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h148)
        v0_1314 <= v0_1314 & ~maskExt_1314 | maskExt_1314 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h148)
        v0_1315 <= v0_1315 & ~maskExt_1315 | maskExt_1315 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h149)
        v0_1316 <= v0_1316 & ~maskExt_1316 | maskExt_1316 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h149)
        v0_1317 <= v0_1317 & ~maskExt_1317 | maskExt_1317 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h149)
        v0_1318 <= v0_1318 & ~maskExt_1318 | maskExt_1318 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h149)
        v0_1319 <= v0_1319 & ~maskExt_1319 | maskExt_1319 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h14A)
        v0_1320 <= v0_1320 & ~maskExt_1320 | maskExt_1320 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h14A)
        v0_1321 <= v0_1321 & ~maskExt_1321 | maskExt_1321 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h14A)
        v0_1322 <= v0_1322 & ~maskExt_1322 | maskExt_1322 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h14A)
        v0_1323 <= v0_1323 & ~maskExt_1323 | maskExt_1323 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h14B)
        v0_1324 <= v0_1324 & ~maskExt_1324 | maskExt_1324 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h14B)
        v0_1325 <= v0_1325 & ~maskExt_1325 | maskExt_1325 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h14B)
        v0_1326 <= v0_1326 & ~maskExt_1326 | maskExt_1326 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h14B)
        v0_1327 <= v0_1327 & ~maskExt_1327 | maskExt_1327 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h14C)
        v0_1328 <= v0_1328 & ~maskExt_1328 | maskExt_1328 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h14C)
        v0_1329 <= v0_1329 & ~maskExt_1329 | maskExt_1329 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h14C)
        v0_1330 <= v0_1330 & ~maskExt_1330 | maskExt_1330 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h14C)
        v0_1331 <= v0_1331 & ~maskExt_1331 | maskExt_1331 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h14D)
        v0_1332 <= v0_1332 & ~maskExt_1332 | maskExt_1332 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h14D)
        v0_1333 <= v0_1333 & ~maskExt_1333 | maskExt_1333 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h14D)
        v0_1334 <= v0_1334 & ~maskExt_1334 | maskExt_1334 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h14D)
        v0_1335 <= v0_1335 & ~maskExt_1335 | maskExt_1335 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h14E)
        v0_1336 <= v0_1336 & ~maskExt_1336 | maskExt_1336 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h14E)
        v0_1337 <= v0_1337 & ~maskExt_1337 | maskExt_1337 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h14E)
        v0_1338 <= v0_1338 & ~maskExt_1338 | maskExt_1338 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h14E)
        v0_1339 <= v0_1339 & ~maskExt_1339 | maskExt_1339 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h14F)
        v0_1340 <= v0_1340 & ~maskExt_1340 | maskExt_1340 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h14F)
        v0_1341 <= v0_1341 & ~maskExt_1341 | maskExt_1341 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h14F)
        v0_1342 <= v0_1342 & ~maskExt_1342 | maskExt_1342 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h14F)
        v0_1343 <= v0_1343 & ~maskExt_1343 | maskExt_1343 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h150)
        v0_1344 <= v0_1344 & ~maskExt_1344 | maskExt_1344 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h150)
        v0_1345 <= v0_1345 & ~maskExt_1345 | maskExt_1345 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h150)
        v0_1346 <= v0_1346 & ~maskExt_1346 | maskExt_1346 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h150)
        v0_1347 <= v0_1347 & ~maskExt_1347 | maskExt_1347 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h151)
        v0_1348 <= v0_1348 & ~maskExt_1348 | maskExt_1348 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h151)
        v0_1349 <= v0_1349 & ~maskExt_1349 | maskExt_1349 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h151)
        v0_1350 <= v0_1350 & ~maskExt_1350 | maskExt_1350 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h151)
        v0_1351 <= v0_1351 & ~maskExt_1351 | maskExt_1351 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h152)
        v0_1352 <= v0_1352 & ~maskExt_1352 | maskExt_1352 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h152)
        v0_1353 <= v0_1353 & ~maskExt_1353 | maskExt_1353 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h152)
        v0_1354 <= v0_1354 & ~maskExt_1354 | maskExt_1354 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h152)
        v0_1355 <= v0_1355 & ~maskExt_1355 | maskExt_1355 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h153)
        v0_1356 <= v0_1356 & ~maskExt_1356 | maskExt_1356 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h153)
        v0_1357 <= v0_1357 & ~maskExt_1357 | maskExt_1357 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h153)
        v0_1358 <= v0_1358 & ~maskExt_1358 | maskExt_1358 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h153)
        v0_1359 <= v0_1359 & ~maskExt_1359 | maskExt_1359 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h154)
        v0_1360 <= v0_1360 & ~maskExt_1360 | maskExt_1360 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h154)
        v0_1361 <= v0_1361 & ~maskExt_1361 | maskExt_1361 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h154)
        v0_1362 <= v0_1362 & ~maskExt_1362 | maskExt_1362 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h154)
        v0_1363 <= v0_1363 & ~maskExt_1363 | maskExt_1363 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h155)
        v0_1364 <= v0_1364 & ~maskExt_1364 | maskExt_1364 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h155)
        v0_1365 <= v0_1365 & ~maskExt_1365 | maskExt_1365 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h155)
        v0_1366 <= v0_1366 & ~maskExt_1366 | maskExt_1366 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h155)
        v0_1367 <= v0_1367 & ~maskExt_1367 | maskExt_1367 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h156)
        v0_1368 <= v0_1368 & ~maskExt_1368 | maskExt_1368 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h156)
        v0_1369 <= v0_1369 & ~maskExt_1369 | maskExt_1369 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h156)
        v0_1370 <= v0_1370 & ~maskExt_1370 | maskExt_1370 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h156)
        v0_1371 <= v0_1371 & ~maskExt_1371 | maskExt_1371 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h157)
        v0_1372 <= v0_1372 & ~maskExt_1372 | maskExt_1372 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h157)
        v0_1373 <= v0_1373 & ~maskExt_1373 | maskExt_1373 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h157)
        v0_1374 <= v0_1374 & ~maskExt_1374 | maskExt_1374 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h157)
        v0_1375 <= v0_1375 & ~maskExt_1375 | maskExt_1375 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h158)
        v0_1376 <= v0_1376 & ~maskExt_1376 | maskExt_1376 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h158)
        v0_1377 <= v0_1377 & ~maskExt_1377 | maskExt_1377 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h158)
        v0_1378 <= v0_1378 & ~maskExt_1378 | maskExt_1378 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h158)
        v0_1379 <= v0_1379 & ~maskExt_1379 | maskExt_1379 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h159)
        v0_1380 <= v0_1380 & ~maskExt_1380 | maskExt_1380 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h159)
        v0_1381 <= v0_1381 & ~maskExt_1381 | maskExt_1381 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h159)
        v0_1382 <= v0_1382 & ~maskExt_1382 | maskExt_1382 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h159)
        v0_1383 <= v0_1383 & ~maskExt_1383 | maskExt_1383 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h15A)
        v0_1384 <= v0_1384 & ~maskExt_1384 | maskExt_1384 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h15A)
        v0_1385 <= v0_1385 & ~maskExt_1385 | maskExt_1385 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h15A)
        v0_1386 <= v0_1386 & ~maskExt_1386 | maskExt_1386 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h15A)
        v0_1387 <= v0_1387 & ~maskExt_1387 | maskExt_1387 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h15B)
        v0_1388 <= v0_1388 & ~maskExt_1388 | maskExt_1388 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h15B)
        v0_1389 <= v0_1389 & ~maskExt_1389 | maskExt_1389 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h15B)
        v0_1390 <= v0_1390 & ~maskExt_1390 | maskExt_1390 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h15B)
        v0_1391 <= v0_1391 & ~maskExt_1391 | maskExt_1391 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h15C)
        v0_1392 <= v0_1392 & ~maskExt_1392 | maskExt_1392 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h15C)
        v0_1393 <= v0_1393 & ~maskExt_1393 | maskExt_1393 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h15C)
        v0_1394 <= v0_1394 & ~maskExt_1394 | maskExt_1394 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h15C)
        v0_1395 <= v0_1395 & ~maskExt_1395 | maskExt_1395 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h15D)
        v0_1396 <= v0_1396 & ~maskExt_1396 | maskExt_1396 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h15D)
        v0_1397 <= v0_1397 & ~maskExt_1397 | maskExt_1397 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h15D)
        v0_1398 <= v0_1398 & ~maskExt_1398 | maskExt_1398 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h15D)
        v0_1399 <= v0_1399 & ~maskExt_1399 | maskExt_1399 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h15E)
        v0_1400 <= v0_1400 & ~maskExt_1400 | maskExt_1400 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h15E)
        v0_1401 <= v0_1401 & ~maskExt_1401 | maskExt_1401 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h15E)
        v0_1402 <= v0_1402 & ~maskExt_1402 | maskExt_1402 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h15E)
        v0_1403 <= v0_1403 & ~maskExt_1403 | maskExt_1403 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h15F)
        v0_1404 <= v0_1404 & ~maskExt_1404 | maskExt_1404 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h15F)
        v0_1405 <= v0_1405 & ~maskExt_1405 | maskExt_1405 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h15F)
        v0_1406 <= v0_1406 & ~maskExt_1406 | maskExt_1406 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h15F)
        v0_1407 <= v0_1407 & ~maskExt_1407 | maskExt_1407 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h160)
        v0_1408 <= v0_1408 & ~maskExt_1408 | maskExt_1408 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h160)
        v0_1409 <= v0_1409 & ~maskExt_1409 | maskExt_1409 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h160)
        v0_1410 <= v0_1410 & ~maskExt_1410 | maskExt_1410 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h160)
        v0_1411 <= v0_1411 & ~maskExt_1411 | maskExt_1411 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h161)
        v0_1412 <= v0_1412 & ~maskExt_1412 | maskExt_1412 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h161)
        v0_1413 <= v0_1413 & ~maskExt_1413 | maskExt_1413 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h161)
        v0_1414 <= v0_1414 & ~maskExt_1414 | maskExt_1414 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h161)
        v0_1415 <= v0_1415 & ~maskExt_1415 | maskExt_1415 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h162)
        v0_1416 <= v0_1416 & ~maskExt_1416 | maskExt_1416 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h162)
        v0_1417 <= v0_1417 & ~maskExt_1417 | maskExt_1417 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h162)
        v0_1418 <= v0_1418 & ~maskExt_1418 | maskExt_1418 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h162)
        v0_1419 <= v0_1419 & ~maskExt_1419 | maskExt_1419 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h163)
        v0_1420 <= v0_1420 & ~maskExt_1420 | maskExt_1420 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h163)
        v0_1421 <= v0_1421 & ~maskExt_1421 | maskExt_1421 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h163)
        v0_1422 <= v0_1422 & ~maskExt_1422 | maskExt_1422 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h163)
        v0_1423 <= v0_1423 & ~maskExt_1423 | maskExt_1423 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h164)
        v0_1424 <= v0_1424 & ~maskExt_1424 | maskExt_1424 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h164)
        v0_1425 <= v0_1425 & ~maskExt_1425 | maskExt_1425 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h164)
        v0_1426 <= v0_1426 & ~maskExt_1426 | maskExt_1426 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h164)
        v0_1427 <= v0_1427 & ~maskExt_1427 | maskExt_1427 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h165)
        v0_1428 <= v0_1428 & ~maskExt_1428 | maskExt_1428 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h165)
        v0_1429 <= v0_1429 & ~maskExt_1429 | maskExt_1429 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h165)
        v0_1430 <= v0_1430 & ~maskExt_1430 | maskExt_1430 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h165)
        v0_1431 <= v0_1431 & ~maskExt_1431 | maskExt_1431 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h166)
        v0_1432 <= v0_1432 & ~maskExt_1432 | maskExt_1432 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h166)
        v0_1433 <= v0_1433 & ~maskExt_1433 | maskExt_1433 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h166)
        v0_1434 <= v0_1434 & ~maskExt_1434 | maskExt_1434 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h166)
        v0_1435 <= v0_1435 & ~maskExt_1435 | maskExt_1435 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h167)
        v0_1436 <= v0_1436 & ~maskExt_1436 | maskExt_1436 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h167)
        v0_1437 <= v0_1437 & ~maskExt_1437 | maskExt_1437 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h167)
        v0_1438 <= v0_1438 & ~maskExt_1438 | maskExt_1438 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h167)
        v0_1439 <= v0_1439 & ~maskExt_1439 | maskExt_1439 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h168)
        v0_1440 <= v0_1440 & ~maskExt_1440 | maskExt_1440 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h168)
        v0_1441 <= v0_1441 & ~maskExt_1441 | maskExt_1441 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h168)
        v0_1442 <= v0_1442 & ~maskExt_1442 | maskExt_1442 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h168)
        v0_1443 <= v0_1443 & ~maskExt_1443 | maskExt_1443 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h169)
        v0_1444 <= v0_1444 & ~maskExt_1444 | maskExt_1444 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h169)
        v0_1445 <= v0_1445 & ~maskExt_1445 | maskExt_1445 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h169)
        v0_1446 <= v0_1446 & ~maskExt_1446 | maskExt_1446 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h169)
        v0_1447 <= v0_1447 & ~maskExt_1447 | maskExt_1447 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h16A)
        v0_1448 <= v0_1448 & ~maskExt_1448 | maskExt_1448 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h16A)
        v0_1449 <= v0_1449 & ~maskExt_1449 | maskExt_1449 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h16A)
        v0_1450 <= v0_1450 & ~maskExt_1450 | maskExt_1450 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h16A)
        v0_1451 <= v0_1451 & ~maskExt_1451 | maskExt_1451 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h16B)
        v0_1452 <= v0_1452 & ~maskExt_1452 | maskExt_1452 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h16B)
        v0_1453 <= v0_1453 & ~maskExt_1453 | maskExt_1453 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h16B)
        v0_1454 <= v0_1454 & ~maskExt_1454 | maskExt_1454 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h16B)
        v0_1455 <= v0_1455 & ~maskExt_1455 | maskExt_1455 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h16C)
        v0_1456 <= v0_1456 & ~maskExt_1456 | maskExt_1456 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h16C)
        v0_1457 <= v0_1457 & ~maskExt_1457 | maskExt_1457 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h16C)
        v0_1458 <= v0_1458 & ~maskExt_1458 | maskExt_1458 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h16C)
        v0_1459 <= v0_1459 & ~maskExt_1459 | maskExt_1459 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h16D)
        v0_1460 <= v0_1460 & ~maskExt_1460 | maskExt_1460 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h16D)
        v0_1461 <= v0_1461 & ~maskExt_1461 | maskExt_1461 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h16D)
        v0_1462 <= v0_1462 & ~maskExt_1462 | maskExt_1462 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h16D)
        v0_1463 <= v0_1463 & ~maskExt_1463 | maskExt_1463 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h16E)
        v0_1464 <= v0_1464 & ~maskExt_1464 | maskExt_1464 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h16E)
        v0_1465 <= v0_1465 & ~maskExt_1465 | maskExt_1465 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h16E)
        v0_1466 <= v0_1466 & ~maskExt_1466 | maskExt_1466 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h16E)
        v0_1467 <= v0_1467 & ~maskExt_1467 | maskExt_1467 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h16F)
        v0_1468 <= v0_1468 & ~maskExt_1468 | maskExt_1468 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h16F)
        v0_1469 <= v0_1469 & ~maskExt_1469 | maskExt_1469 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h16F)
        v0_1470 <= v0_1470 & ~maskExt_1470 | maskExt_1470 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h16F)
        v0_1471 <= v0_1471 & ~maskExt_1471 | maskExt_1471 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h170)
        v0_1472 <= v0_1472 & ~maskExt_1472 | maskExt_1472 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h170)
        v0_1473 <= v0_1473 & ~maskExt_1473 | maskExt_1473 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h170)
        v0_1474 <= v0_1474 & ~maskExt_1474 | maskExt_1474 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h170)
        v0_1475 <= v0_1475 & ~maskExt_1475 | maskExt_1475 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h171)
        v0_1476 <= v0_1476 & ~maskExt_1476 | maskExt_1476 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h171)
        v0_1477 <= v0_1477 & ~maskExt_1477 | maskExt_1477 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h171)
        v0_1478 <= v0_1478 & ~maskExt_1478 | maskExt_1478 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h171)
        v0_1479 <= v0_1479 & ~maskExt_1479 | maskExt_1479 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h172)
        v0_1480 <= v0_1480 & ~maskExt_1480 | maskExt_1480 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h172)
        v0_1481 <= v0_1481 & ~maskExt_1481 | maskExt_1481 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h172)
        v0_1482 <= v0_1482 & ~maskExt_1482 | maskExt_1482 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h172)
        v0_1483 <= v0_1483 & ~maskExt_1483 | maskExt_1483 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h173)
        v0_1484 <= v0_1484 & ~maskExt_1484 | maskExt_1484 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h173)
        v0_1485 <= v0_1485 & ~maskExt_1485 | maskExt_1485 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h173)
        v0_1486 <= v0_1486 & ~maskExt_1486 | maskExt_1486 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h173)
        v0_1487 <= v0_1487 & ~maskExt_1487 | maskExt_1487 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h174)
        v0_1488 <= v0_1488 & ~maskExt_1488 | maskExt_1488 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h174)
        v0_1489 <= v0_1489 & ~maskExt_1489 | maskExt_1489 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h174)
        v0_1490 <= v0_1490 & ~maskExt_1490 | maskExt_1490 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h174)
        v0_1491 <= v0_1491 & ~maskExt_1491 | maskExt_1491 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h175)
        v0_1492 <= v0_1492 & ~maskExt_1492 | maskExt_1492 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h175)
        v0_1493 <= v0_1493 & ~maskExt_1493 | maskExt_1493 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h175)
        v0_1494 <= v0_1494 & ~maskExt_1494 | maskExt_1494 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h175)
        v0_1495 <= v0_1495 & ~maskExt_1495 | maskExt_1495 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h176)
        v0_1496 <= v0_1496 & ~maskExt_1496 | maskExt_1496 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h176)
        v0_1497 <= v0_1497 & ~maskExt_1497 | maskExt_1497 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h176)
        v0_1498 <= v0_1498 & ~maskExt_1498 | maskExt_1498 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h176)
        v0_1499 <= v0_1499 & ~maskExt_1499 | maskExt_1499 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h177)
        v0_1500 <= v0_1500 & ~maskExt_1500 | maskExt_1500 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h177)
        v0_1501 <= v0_1501 & ~maskExt_1501 | maskExt_1501 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h177)
        v0_1502 <= v0_1502 & ~maskExt_1502 | maskExt_1502 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h177)
        v0_1503 <= v0_1503 & ~maskExt_1503 | maskExt_1503 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h178)
        v0_1504 <= v0_1504 & ~maskExt_1504 | maskExt_1504 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h178)
        v0_1505 <= v0_1505 & ~maskExt_1505 | maskExt_1505 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h178)
        v0_1506 <= v0_1506 & ~maskExt_1506 | maskExt_1506 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h178)
        v0_1507 <= v0_1507 & ~maskExt_1507 | maskExt_1507 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h179)
        v0_1508 <= v0_1508 & ~maskExt_1508 | maskExt_1508 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h179)
        v0_1509 <= v0_1509 & ~maskExt_1509 | maskExt_1509 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h179)
        v0_1510 <= v0_1510 & ~maskExt_1510 | maskExt_1510 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h179)
        v0_1511 <= v0_1511 & ~maskExt_1511 | maskExt_1511 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h17A)
        v0_1512 <= v0_1512 & ~maskExt_1512 | maskExt_1512 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h17A)
        v0_1513 <= v0_1513 & ~maskExt_1513 | maskExt_1513 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h17A)
        v0_1514 <= v0_1514 & ~maskExt_1514 | maskExt_1514 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h17A)
        v0_1515 <= v0_1515 & ~maskExt_1515 | maskExt_1515 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h17B)
        v0_1516 <= v0_1516 & ~maskExt_1516 | maskExt_1516 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h17B)
        v0_1517 <= v0_1517 & ~maskExt_1517 | maskExt_1517 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h17B)
        v0_1518 <= v0_1518 & ~maskExt_1518 | maskExt_1518 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h17B)
        v0_1519 <= v0_1519 & ~maskExt_1519 | maskExt_1519 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h17C)
        v0_1520 <= v0_1520 & ~maskExt_1520 | maskExt_1520 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h17C)
        v0_1521 <= v0_1521 & ~maskExt_1521 | maskExt_1521 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h17C)
        v0_1522 <= v0_1522 & ~maskExt_1522 | maskExt_1522 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h17C)
        v0_1523 <= v0_1523 & ~maskExt_1523 | maskExt_1523 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h17D)
        v0_1524 <= v0_1524 & ~maskExt_1524 | maskExt_1524 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h17D)
        v0_1525 <= v0_1525 & ~maskExt_1525 | maskExt_1525 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h17D)
        v0_1526 <= v0_1526 & ~maskExt_1526 | maskExt_1526 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h17D)
        v0_1527 <= v0_1527 & ~maskExt_1527 | maskExt_1527 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h17E)
        v0_1528 <= v0_1528 & ~maskExt_1528 | maskExt_1528 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h17E)
        v0_1529 <= v0_1529 & ~maskExt_1529 | maskExt_1529 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h17E)
        v0_1530 <= v0_1530 & ~maskExt_1530 | maskExt_1530 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h17E)
        v0_1531 <= v0_1531 & ~maskExt_1531 | maskExt_1531 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h17F)
        v0_1532 <= v0_1532 & ~maskExt_1532 | maskExt_1532 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h17F)
        v0_1533 <= v0_1533 & ~maskExt_1533 | maskExt_1533 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h17F)
        v0_1534 <= v0_1534 & ~maskExt_1534 | maskExt_1534 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h17F)
        v0_1535 <= v0_1535 & ~maskExt_1535 | maskExt_1535 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h180)
        v0_1536 <= v0_1536 & ~maskExt_1536 | maskExt_1536 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h180)
        v0_1537 <= v0_1537 & ~maskExt_1537 | maskExt_1537 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h180)
        v0_1538 <= v0_1538 & ~maskExt_1538 | maskExt_1538 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h180)
        v0_1539 <= v0_1539 & ~maskExt_1539 | maskExt_1539 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h181)
        v0_1540 <= v0_1540 & ~maskExt_1540 | maskExt_1540 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h181)
        v0_1541 <= v0_1541 & ~maskExt_1541 | maskExt_1541 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h181)
        v0_1542 <= v0_1542 & ~maskExt_1542 | maskExt_1542 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h181)
        v0_1543 <= v0_1543 & ~maskExt_1543 | maskExt_1543 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h182)
        v0_1544 <= v0_1544 & ~maskExt_1544 | maskExt_1544 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h182)
        v0_1545 <= v0_1545 & ~maskExt_1545 | maskExt_1545 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h182)
        v0_1546 <= v0_1546 & ~maskExt_1546 | maskExt_1546 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h182)
        v0_1547 <= v0_1547 & ~maskExt_1547 | maskExt_1547 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h183)
        v0_1548 <= v0_1548 & ~maskExt_1548 | maskExt_1548 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h183)
        v0_1549 <= v0_1549 & ~maskExt_1549 | maskExt_1549 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h183)
        v0_1550 <= v0_1550 & ~maskExt_1550 | maskExt_1550 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h183)
        v0_1551 <= v0_1551 & ~maskExt_1551 | maskExt_1551 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h184)
        v0_1552 <= v0_1552 & ~maskExt_1552 | maskExt_1552 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h184)
        v0_1553 <= v0_1553 & ~maskExt_1553 | maskExt_1553 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h184)
        v0_1554 <= v0_1554 & ~maskExt_1554 | maskExt_1554 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h184)
        v0_1555 <= v0_1555 & ~maskExt_1555 | maskExt_1555 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h185)
        v0_1556 <= v0_1556 & ~maskExt_1556 | maskExt_1556 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h185)
        v0_1557 <= v0_1557 & ~maskExt_1557 | maskExt_1557 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h185)
        v0_1558 <= v0_1558 & ~maskExt_1558 | maskExt_1558 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h185)
        v0_1559 <= v0_1559 & ~maskExt_1559 | maskExt_1559 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h186)
        v0_1560 <= v0_1560 & ~maskExt_1560 | maskExt_1560 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h186)
        v0_1561 <= v0_1561 & ~maskExt_1561 | maskExt_1561 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h186)
        v0_1562 <= v0_1562 & ~maskExt_1562 | maskExt_1562 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h186)
        v0_1563 <= v0_1563 & ~maskExt_1563 | maskExt_1563 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h187)
        v0_1564 <= v0_1564 & ~maskExt_1564 | maskExt_1564 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h187)
        v0_1565 <= v0_1565 & ~maskExt_1565 | maskExt_1565 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h187)
        v0_1566 <= v0_1566 & ~maskExt_1566 | maskExt_1566 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h187)
        v0_1567 <= v0_1567 & ~maskExt_1567 | maskExt_1567 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h188)
        v0_1568 <= v0_1568 & ~maskExt_1568 | maskExt_1568 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h188)
        v0_1569 <= v0_1569 & ~maskExt_1569 | maskExt_1569 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h188)
        v0_1570 <= v0_1570 & ~maskExt_1570 | maskExt_1570 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h188)
        v0_1571 <= v0_1571 & ~maskExt_1571 | maskExt_1571 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h189)
        v0_1572 <= v0_1572 & ~maskExt_1572 | maskExt_1572 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h189)
        v0_1573 <= v0_1573 & ~maskExt_1573 | maskExt_1573 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h189)
        v0_1574 <= v0_1574 & ~maskExt_1574 | maskExt_1574 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h189)
        v0_1575 <= v0_1575 & ~maskExt_1575 | maskExt_1575 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h18A)
        v0_1576 <= v0_1576 & ~maskExt_1576 | maskExt_1576 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h18A)
        v0_1577 <= v0_1577 & ~maskExt_1577 | maskExt_1577 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h18A)
        v0_1578 <= v0_1578 & ~maskExt_1578 | maskExt_1578 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h18A)
        v0_1579 <= v0_1579 & ~maskExt_1579 | maskExt_1579 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h18B)
        v0_1580 <= v0_1580 & ~maskExt_1580 | maskExt_1580 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h18B)
        v0_1581 <= v0_1581 & ~maskExt_1581 | maskExt_1581 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h18B)
        v0_1582 <= v0_1582 & ~maskExt_1582 | maskExt_1582 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h18B)
        v0_1583 <= v0_1583 & ~maskExt_1583 | maskExt_1583 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h18C)
        v0_1584 <= v0_1584 & ~maskExt_1584 | maskExt_1584 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h18C)
        v0_1585 <= v0_1585 & ~maskExt_1585 | maskExt_1585 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h18C)
        v0_1586 <= v0_1586 & ~maskExt_1586 | maskExt_1586 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h18C)
        v0_1587 <= v0_1587 & ~maskExt_1587 | maskExt_1587 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h18D)
        v0_1588 <= v0_1588 & ~maskExt_1588 | maskExt_1588 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h18D)
        v0_1589 <= v0_1589 & ~maskExt_1589 | maskExt_1589 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h18D)
        v0_1590 <= v0_1590 & ~maskExt_1590 | maskExt_1590 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h18D)
        v0_1591 <= v0_1591 & ~maskExt_1591 | maskExt_1591 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h18E)
        v0_1592 <= v0_1592 & ~maskExt_1592 | maskExt_1592 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h18E)
        v0_1593 <= v0_1593 & ~maskExt_1593 | maskExt_1593 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h18E)
        v0_1594 <= v0_1594 & ~maskExt_1594 | maskExt_1594 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h18E)
        v0_1595 <= v0_1595 & ~maskExt_1595 | maskExt_1595 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h18F)
        v0_1596 <= v0_1596 & ~maskExt_1596 | maskExt_1596 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h18F)
        v0_1597 <= v0_1597 & ~maskExt_1597 | maskExt_1597 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h18F)
        v0_1598 <= v0_1598 & ~maskExt_1598 | maskExt_1598 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h18F)
        v0_1599 <= v0_1599 & ~maskExt_1599 | maskExt_1599 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h190)
        v0_1600 <= v0_1600 & ~maskExt_1600 | maskExt_1600 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h190)
        v0_1601 <= v0_1601 & ~maskExt_1601 | maskExt_1601 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h190)
        v0_1602 <= v0_1602 & ~maskExt_1602 | maskExt_1602 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h190)
        v0_1603 <= v0_1603 & ~maskExt_1603 | maskExt_1603 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h191)
        v0_1604 <= v0_1604 & ~maskExt_1604 | maskExt_1604 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h191)
        v0_1605 <= v0_1605 & ~maskExt_1605 | maskExt_1605 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h191)
        v0_1606 <= v0_1606 & ~maskExt_1606 | maskExt_1606 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h191)
        v0_1607 <= v0_1607 & ~maskExt_1607 | maskExt_1607 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h192)
        v0_1608 <= v0_1608 & ~maskExt_1608 | maskExt_1608 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h192)
        v0_1609 <= v0_1609 & ~maskExt_1609 | maskExt_1609 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h192)
        v0_1610 <= v0_1610 & ~maskExt_1610 | maskExt_1610 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h192)
        v0_1611 <= v0_1611 & ~maskExt_1611 | maskExt_1611 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h193)
        v0_1612 <= v0_1612 & ~maskExt_1612 | maskExt_1612 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h193)
        v0_1613 <= v0_1613 & ~maskExt_1613 | maskExt_1613 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h193)
        v0_1614 <= v0_1614 & ~maskExt_1614 | maskExt_1614 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h193)
        v0_1615 <= v0_1615 & ~maskExt_1615 | maskExt_1615 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h194)
        v0_1616 <= v0_1616 & ~maskExt_1616 | maskExt_1616 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h194)
        v0_1617 <= v0_1617 & ~maskExt_1617 | maskExt_1617 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h194)
        v0_1618 <= v0_1618 & ~maskExt_1618 | maskExt_1618 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h194)
        v0_1619 <= v0_1619 & ~maskExt_1619 | maskExt_1619 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h195)
        v0_1620 <= v0_1620 & ~maskExt_1620 | maskExt_1620 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h195)
        v0_1621 <= v0_1621 & ~maskExt_1621 | maskExt_1621 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h195)
        v0_1622 <= v0_1622 & ~maskExt_1622 | maskExt_1622 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h195)
        v0_1623 <= v0_1623 & ~maskExt_1623 | maskExt_1623 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h196)
        v0_1624 <= v0_1624 & ~maskExt_1624 | maskExt_1624 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h196)
        v0_1625 <= v0_1625 & ~maskExt_1625 | maskExt_1625 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h196)
        v0_1626 <= v0_1626 & ~maskExt_1626 | maskExt_1626 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h196)
        v0_1627 <= v0_1627 & ~maskExt_1627 | maskExt_1627 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h197)
        v0_1628 <= v0_1628 & ~maskExt_1628 | maskExt_1628 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h197)
        v0_1629 <= v0_1629 & ~maskExt_1629 | maskExt_1629 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h197)
        v0_1630 <= v0_1630 & ~maskExt_1630 | maskExt_1630 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h197)
        v0_1631 <= v0_1631 & ~maskExt_1631 | maskExt_1631 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h198)
        v0_1632 <= v0_1632 & ~maskExt_1632 | maskExt_1632 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h198)
        v0_1633 <= v0_1633 & ~maskExt_1633 | maskExt_1633 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h198)
        v0_1634 <= v0_1634 & ~maskExt_1634 | maskExt_1634 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h198)
        v0_1635 <= v0_1635 & ~maskExt_1635 | maskExt_1635 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h199)
        v0_1636 <= v0_1636 & ~maskExt_1636 | maskExt_1636 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h199)
        v0_1637 <= v0_1637 & ~maskExt_1637 | maskExt_1637 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h199)
        v0_1638 <= v0_1638 & ~maskExt_1638 | maskExt_1638 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h199)
        v0_1639 <= v0_1639 & ~maskExt_1639 | maskExt_1639 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h19A)
        v0_1640 <= v0_1640 & ~maskExt_1640 | maskExt_1640 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h19A)
        v0_1641 <= v0_1641 & ~maskExt_1641 | maskExt_1641 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h19A)
        v0_1642 <= v0_1642 & ~maskExt_1642 | maskExt_1642 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h19A)
        v0_1643 <= v0_1643 & ~maskExt_1643 | maskExt_1643 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h19B)
        v0_1644 <= v0_1644 & ~maskExt_1644 | maskExt_1644 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h19B)
        v0_1645 <= v0_1645 & ~maskExt_1645 | maskExt_1645 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h19B)
        v0_1646 <= v0_1646 & ~maskExt_1646 | maskExt_1646 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h19B)
        v0_1647 <= v0_1647 & ~maskExt_1647 | maskExt_1647 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h19C)
        v0_1648 <= v0_1648 & ~maskExt_1648 | maskExt_1648 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h19C)
        v0_1649 <= v0_1649 & ~maskExt_1649 | maskExt_1649 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h19C)
        v0_1650 <= v0_1650 & ~maskExt_1650 | maskExt_1650 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h19C)
        v0_1651 <= v0_1651 & ~maskExt_1651 | maskExt_1651 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h19D)
        v0_1652 <= v0_1652 & ~maskExt_1652 | maskExt_1652 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h19D)
        v0_1653 <= v0_1653 & ~maskExt_1653 | maskExt_1653 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h19D)
        v0_1654 <= v0_1654 & ~maskExt_1654 | maskExt_1654 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h19D)
        v0_1655 <= v0_1655 & ~maskExt_1655 | maskExt_1655 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h19E)
        v0_1656 <= v0_1656 & ~maskExt_1656 | maskExt_1656 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h19E)
        v0_1657 <= v0_1657 & ~maskExt_1657 | maskExt_1657 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h19E)
        v0_1658 <= v0_1658 & ~maskExt_1658 | maskExt_1658 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h19E)
        v0_1659 <= v0_1659 & ~maskExt_1659 | maskExt_1659 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h19F)
        v0_1660 <= v0_1660 & ~maskExt_1660 | maskExt_1660 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h19F)
        v0_1661 <= v0_1661 & ~maskExt_1661 | maskExt_1661 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h19F)
        v0_1662 <= v0_1662 & ~maskExt_1662 | maskExt_1662 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h19F)
        v0_1663 <= v0_1663 & ~maskExt_1663 | maskExt_1663 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1A0)
        v0_1664 <= v0_1664 & ~maskExt_1664 | maskExt_1664 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1A0)
        v0_1665 <= v0_1665 & ~maskExt_1665 | maskExt_1665 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1A0)
        v0_1666 <= v0_1666 & ~maskExt_1666 | maskExt_1666 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1A0)
        v0_1667 <= v0_1667 & ~maskExt_1667 | maskExt_1667 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1A1)
        v0_1668 <= v0_1668 & ~maskExt_1668 | maskExt_1668 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1A1)
        v0_1669 <= v0_1669 & ~maskExt_1669 | maskExt_1669 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1A1)
        v0_1670 <= v0_1670 & ~maskExt_1670 | maskExt_1670 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1A1)
        v0_1671 <= v0_1671 & ~maskExt_1671 | maskExt_1671 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1A2)
        v0_1672 <= v0_1672 & ~maskExt_1672 | maskExt_1672 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1A2)
        v0_1673 <= v0_1673 & ~maskExt_1673 | maskExt_1673 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1A2)
        v0_1674 <= v0_1674 & ~maskExt_1674 | maskExt_1674 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1A2)
        v0_1675 <= v0_1675 & ~maskExt_1675 | maskExt_1675 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1A3)
        v0_1676 <= v0_1676 & ~maskExt_1676 | maskExt_1676 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1A3)
        v0_1677 <= v0_1677 & ~maskExt_1677 | maskExt_1677 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1A3)
        v0_1678 <= v0_1678 & ~maskExt_1678 | maskExt_1678 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1A3)
        v0_1679 <= v0_1679 & ~maskExt_1679 | maskExt_1679 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1A4)
        v0_1680 <= v0_1680 & ~maskExt_1680 | maskExt_1680 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1A4)
        v0_1681 <= v0_1681 & ~maskExt_1681 | maskExt_1681 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1A4)
        v0_1682 <= v0_1682 & ~maskExt_1682 | maskExt_1682 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1A4)
        v0_1683 <= v0_1683 & ~maskExt_1683 | maskExt_1683 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1A5)
        v0_1684 <= v0_1684 & ~maskExt_1684 | maskExt_1684 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1A5)
        v0_1685 <= v0_1685 & ~maskExt_1685 | maskExt_1685 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1A5)
        v0_1686 <= v0_1686 & ~maskExt_1686 | maskExt_1686 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1A5)
        v0_1687 <= v0_1687 & ~maskExt_1687 | maskExt_1687 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1A6)
        v0_1688 <= v0_1688 & ~maskExt_1688 | maskExt_1688 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1A6)
        v0_1689 <= v0_1689 & ~maskExt_1689 | maskExt_1689 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1A6)
        v0_1690 <= v0_1690 & ~maskExt_1690 | maskExt_1690 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1A6)
        v0_1691 <= v0_1691 & ~maskExt_1691 | maskExt_1691 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1A7)
        v0_1692 <= v0_1692 & ~maskExt_1692 | maskExt_1692 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1A7)
        v0_1693 <= v0_1693 & ~maskExt_1693 | maskExt_1693 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1A7)
        v0_1694 <= v0_1694 & ~maskExt_1694 | maskExt_1694 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1A7)
        v0_1695 <= v0_1695 & ~maskExt_1695 | maskExt_1695 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1A8)
        v0_1696 <= v0_1696 & ~maskExt_1696 | maskExt_1696 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1A8)
        v0_1697 <= v0_1697 & ~maskExt_1697 | maskExt_1697 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1A8)
        v0_1698 <= v0_1698 & ~maskExt_1698 | maskExt_1698 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1A8)
        v0_1699 <= v0_1699 & ~maskExt_1699 | maskExt_1699 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1A9)
        v0_1700 <= v0_1700 & ~maskExt_1700 | maskExt_1700 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1A9)
        v0_1701 <= v0_1701 & ~maskExt_1701 | maskExt_1701 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1A9)
        v0_1702 <= v0_1702 & ~maskExt_1702 | maskExt_1702 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1A9)
        v0_1703 <= v0_1703 & ~maskExt_1703 | maskExt_1703 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1AA)
        v0_1704 <= v0_1704 & ~maskExt_1704 | maskExt_1704 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1AA)
        v0_1705 <= v0_1705 & ~maskExt_1705 | maskExt_1705 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1AA)
        v0_1706 <= v0_1706 & ~maskExt_1706 | maskExt_1706 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1AA)
        v0_1707 <= v0_1707 & ~maskExt_1707 | maskExt_1707 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1AB)
        v0_1708 <= v0_1708 & ~maskExt_1708 | maskExt_1708 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1AB)
        v0_1709 <= v0_1709 & ~maskExt_1709 | maskExt_1709 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1AB)
        v0_1710 <= v0_1710 & ~maskExt_1710 | maskExt_1710 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1AB)
        v0_1711 <= v0_1711 & ~maskExt_1711 | maskExt_1711 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1AC)
        v0_1712 <= v0_1712 & ~maskExt_1712 | maskExt_1712 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1AC)
        v0_1713 <= v0_1713 & ~maskExt_1713 | maskExt_1713 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1AC)
        v0_1714 <= v0_1714 & ~maskExt_1714 | maskExt_1714 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1AC)
        v0_1715 <= v0_1715 & ~maskExt_1715 | maskExt_1715 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1AD)
        v0_1716 <= v0_1716 & ~maskExt_1716 | maskExt_1716 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1AD)
        v0_1717 <= v0_1717 & ~maskExt_1717 | maskExt_1717 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1AD)
        v0_1718 <= v0_1718 & ~maskExt_1718 | maskExt_1718 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1AD)
        v0_1719 <= v0_1719 & ~maskExt_1719 | maskExt_1719 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1AE)
        v0_1720 <= v0_1720 & ~maskExt_1720 | maskExt_1720 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1AE)
        v0_1721 <= v0_1721 & ~maskExt_1721 | maskExt_1721 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1AE)
        v0_1722 <= v0_1722 & ~maskExt_1722 | maskExt_1722 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1AE)
        v0_1723 <= v0_1723 & ~maskExt_1723 | maskExt_1723 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1AF)
        v0_1724 <= v0_1724 & ~maskExt_1724 | maskExt_1724 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1AF)
        v0_1725 <= v0_1725 & ~maskExt_1725 | maskExt_1725 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1AF)
        v0_1726 <= v0_1726 & ~maskExt_1726 | maskExt_1726 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1AF)
        v0_1727 <= v0_1727 & ~maskExt_1727 | maskExt_1727 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1B0)
        v0_1728 <= v0_1728 & ~maskExt_1728 | maskExt_1728 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1B0)
        v0_1729 <= v0_1729 & ~maskExt_1729 | maskExt_1729 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1B0)
        v0_1730 <= v0_1730 & ~maskExt_1730 | maskExt_1730 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1B0)
        v0_1731 <= v0_1731 & ~maskExt_1731 | maskExt_1731 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1B1)
        v0_1732 <= v0_1732 & ~maskExt_1732 | maskExt_1732 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1B1)
        v0_1733 <= v0_1733 & ~maskExt_1733 | maskExt_1733 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1B1)
        v0_1734 <= v0_1734 & ~maskExt_1734 | maskExt_1734 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1B1)
        v0_1735 <= v0_1735 & ~maskExt_1735 | maskExt_1735 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1B2)
        v0_1736 <= v0_1736 & ~maskExt_1736 | maskExt_1736 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1B2)
        v0_1737 <= v0_1737 & ~maskExt_1737 | maskExt_1737 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1B2)
        v0_1738 <= v0_1738 & ~maskExt_1738 | maskExt_1738 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1B2)
        v0_1739 <= v0_1739 & ~maskExt_1739 | maskExt_1739 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1B3)
        v0_1740 <= v0_1740 & ~maskExt_1740 | maskExt_1740 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1B3)
        v0_1741 <= v0_1741 & ~maskExt_1741 | maskExt_1741 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1B3)
        v0_1742 <= v0_1742 & ~maskExt_1742 | maskExt_1742 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1B3)
        v0_1743 <= v0_1743 & ~maskExt_1743 | maskExt_1743 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1B4)
        v0_1744 <= v0_1744 & ~maskExt_1744 | maskExt_1744 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1B4)
        v0_1745 <= v0_1745 & ~maskExt_1745 | maskExt_1745 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1B4)
        v0_1746 <= v0_1746 & ~maskExt_1746 | maskExt_1746 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1B4)
        v0_1747 <= v0_1747 & ~maskExt_1747 | maskExt_1747 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1B5)
        v0_1748 <= v0_1748 & ~maskExt_1748 | maskExt_1748 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1B5)
        v0_1749 <= v0_1749 & ~maskExt_1749 | maskExt_1749 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1B5)
        v0_1750 <= v0_1750 & ~maskExt_1750 | maskExt_1750 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1B5)
        v0_1751 <= v0_1751 & ~maskExt_1751 | maskExt_1751 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1B6)
        v0_1752 <= v0_1752 & ~maskExt_1752 | maskExt_1752 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1B6)
        v0_1753 <= v0_1753 & ~maskExt_1753 | maskExt_1753 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1B6)
        v0_1754 <= v0_1754 & ~maskExt_1754 | maskExt_1754 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1B6)
        v0_1755 <= v0_1755 & ~maskExt_1755 | maskExt_1755 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1B7)
        v0_1756 <= v0_1756 & ~maskExt_1756 | maskExt_1756 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1B7)
        v0_1757 <= v0_1757 & ~maskExt_1757 | maskExt_1757 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1B7)
        v0_1758 <= v0_1758 & ~maskExt_1758 | maskExt_1758 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1B7)
        v0_1759 <= v0_1759 & ~maskExt_1759 | maskExt_1759 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1B8)
        v0_1760 <= v0_1760 & ~maskExt_1760 | maskExt_1760 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1B8)
        v0_1761 <= v0_1761 & ~maskExt_1761 | maskExt_1761 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1B8)
        v0_1762 <= v0_1762 & ~maskExt_1762 | maskExt_1762 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1B8)
        v0_1763 <= v0_1763 & ~maskExt_1763 | maskExt_1763 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1B9)
        v0_1764 <= v0_1764 & ~maskExt_1764 | maskExt_1764 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1B9)
        v0_1765 <= v0_1765 & ~maskExt_1765 | maskExt_1765 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1B9)
        v0_1766 <= v0_1766 & ~maskExt_1766 | maskExt_1766 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1B9)
        v0_1767 <= v0_1767 & ~maskExt_1767 | maskExt_1767 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1BA)
        v0_1768 <= v0_1768 & ~maskExt_1768 | maskExt_1768 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1BA)
        v0_1769 <= v0_1769 & ~maskExt_1769 | maskExt_1769 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1BA)
        v0_1770 <= v0_1770 & ~maskExt_1770 | maskExt_1770 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1BA)
        v0_1771 <= v0_1771 & ~maskExt_1771 | maskExt_1771 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1BB)
        v0_1772 <= v0_1772 & ~maskExt_1772 | maskExt_1772 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1BB)
        v0_1773 <= v0_1773 & ~maskExt_1773 | maskExt_1773 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1BB)
        v0_1774 <= v0_1774 & ~maskExt_1774 | maskExt_1774 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1BB)
        v0_1775 <= v0_1775 & ~maskExt_1775 | maskExt_1775 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1BC)
        v0_1776 <= v0_1776 & ~maskExt_1776 | maskExt_1776 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1BC)
        v0_1777 <= v0_1777 & ~maskExt_1777 | maskExt_1777 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1BC)
        v0_1778 <= v0_1778 & ~maskExt_1778 | maskExt_1778 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1BC)
        v0_1779 <= v0_1779 & ~maskExt_1779 | maskExt_1779 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1BD)
        v0_1780 <= v0_1780 & ~maskExt_1780 | maskExt_1780 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1BD)
        v0_1781 <= v0_1781 & ~maskExt_1781 | maskExt_1781 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1BD)
        v0_1782 <= v0_1782 & ~maskExt_1782 | maskExt_1782 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1BD)
        v0_1783 <= v0_1783 & ~maskExt_1783 | maskExt_1783 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1BE)
        v0_1784 <= v0_1784 & ~maskExt_1784 | maskExt_1784 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1BE)
        v0_1785 <= v0_1785 & ~maskExt_1785 | maskExt_1785 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1BE)
        v0_1786 <= v0_1786 & ~maskExt_1786 | maskExt_1786 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1BE)
        v0_1787 <= v0_1787 & ~maskExt_1787 | maskExt_1787 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1BF)
        v0_1788 <= v0_1788 & ~maskExt_1788 | maskExt_1788 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1BF)
        v0_1789 <= v0_1789 & ~maskExt_1789 | maskExt_1789 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1BF)
        v0_1790 <= v0_1790 & ~maskExt_1790 | maskExt_1790 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1BF)
        v0_1791 <= v0_1791 & ~maskExt_1791 | maskExt_1791 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1C0)
        v0_1792 <= v0_1792 & ~maskExt_1792 | maskExt_1792 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1C0)
        v0_1793 <= v0_1793 & ~maskExt_1793 | maskExt_1793 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1C0)
        v0_1794 <= v0_1794 & ~maskExt_1794 | maskExt_1794 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1C0)
        v0_1795 <= v0_1795 & ~maskExt_1795 | maskExt_1795 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1C1)
        v0_1796 <= v0_1796 & ~maskExt_1796 | maskExt_1796 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1C1)
        v0_1797 <= v0_1797 & ~maskExt_1797 | maskExt_1797 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1C1)
        v0_1798 <= v0_1798 & ~maskExt_1798 | maskExt_1798 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1C1)
        v0_1799 <= v0_1799 & ~maskExt_1799 | maskExt_1799 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1C2)
        v0_1800 <= v0_1800 & ~maskExt_1800 | maskExt_1800 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1C2)
        v0_1801 <= v0_1801 & ~maskExt_1801 | maskExt_1801 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1C2)
        v0_1802 <= v0_1802 & ~maskExt_1802 | maskExt_1802 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1C2)
        v0_1803 <= v0_1803 & ~maskExt_1803 | maskExt_1803 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1C3)
        v0_1804 <= v0_1804 & ~maskExt_1804 | maskExt_1804 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1C3)
        v0_1805 <= v0_1805 & ~maskExt_1805 | maskExt_1805 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1C3)
        v0_1806 <= v0_1806 & ~maskExt_1806 | maskExt_1806 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1C3)
        v0_1807 <= v0_1807 & ~maskExt_1807 | maskExt_1807 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1C4)
        v0_1808 <= v0_1808 & ~maskExt_1808 | maskExt_1808 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1C4)
        v0_1809 <= v0_1809 & ~maskExt_1809 | maskExt_1809 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1C4)
        v0_1810 <= v0_1810 & ~maskExt_1810 | maskExt_1810 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1C4)
        v0_1811 <= v0_1811 & ~maskExt_1811 | maskExt_1811 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1C5)
        v0_1812 <= v0_1812 & ~maskExt_1812 | maskExt_1812 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1C5)
        v0_1813 <= v0_1813 & ~maskExt_1813 | maskExt_1813 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1C5)
        v0_1814 <= v0_1814 & ~maskExt_1814 | maskExt_1814 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1C5)
        v0_1815 <= v0_1815 & ~maskExt_1815 | maskExt_1815 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1C6)
        v0_1816 <= v0_1816 & ~maskExt_1816 | maskExt_1816 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1C6)
        v0_1817 <= v0_1817 & ~maskExt_1817 | maskExt_1817 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1C6)
        v0_1818 <= v0_1818 & ~maskExt_1818 | maskExt_1818 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1C6)
        v0_1819 <= v0_1819 & ~maskExt_1819 | maskExt_1819 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1C7)
        v0_1820 <= v0_1820 & ~maskExt_1820 | maskExt_1820 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1C7)
        v0_1821 <= v0_1821 & ~maskExt_1821 | maskExt_1821 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1C7)
        v0_1822 <= v0_1822 & ~maskExt_1822 | maskExt_1822 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1C7)
        v0_1823 <= v0_1823 & ~maskExt_1823 | maskExt_1823 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1C8)
        v0_1824 <= v0_1824 & ~maskExt_1824 | maskExt_1824 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1C8)
        v0_1825 <= v0_1825 & ~maskExt_1825 | maskExt_1825 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1C8)
        v0_1826 <= v0_1826 & ~maskExt_1826 | maskExt_1826 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1C8)
        v0_1827 <= v0_1827 & ~maskExt_1827 | maskExt_1827 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1C9)
        v0_1828 <= v0_1828 & ~maskExt_1828 | maskExt_1828 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1C9)
        v0_1829 <= v0_1829 & ~maskExt_1829 | maskExt_1829 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1C9)
        v0_1830 <= v0_1830 & ~maskExt_1830 | maskExt_1830 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1C9)
        v0_1831 <= v0_1831 & ~maskExt_1831 | maskExt_1831 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1CA)
        v0_1832 <= v0_1832 & ~maskExt_1832 | maskExt_1832 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1CA)
        v0_1833 <= v0_1833 & ~maskExt_1833 | maskExt_1833 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1CA)
        v0_1834 <= v0_1834 & ~maskExt_1834 | maskExt_1834 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1CA)
        v0_1835 <= v0_1835 & ~maskExt_1835 | maskExt_1835 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1CB)
        v0_1836 <= v0_1836 & ~maskExt_1836 | maskExt_1836 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1CB)
        v0_1837 <= v0_1837 & ~maskExt_1837 | maskExt_1837 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1CB)
        v0_1838 <= v0_1838 & ~maskExt_1838 | maskExt_1838 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1CB)
        v0_1839 <= v0_1839 & ~maskExt_1839 | maskExt_1839 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1CC)
        v0_1840 <= v0_1840 & ~maskExt_1840 | maskExt_1840 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1CC)
        v0_1841 <= v0_1841 & ~maskExt_1841 | maskExt_1841 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1CC)
        v0_1842 <= v0_1842 & ~maskExt_1842 | maskExt_1842 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1CC)
        v0_1843 <= v0_1843 & ~maskExt_1843 | maskExt_1843 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1CD)
        v0_1844 <= v0_1844 & ~maskExt_1844 | maskExt_1844 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1CD)
        v0_1845 <= v0_1845 & ~maskExt_1845 | maskExt_1845 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1CD)
        v0_1846 <= v0_1846 & ~maskExt_1846 | maskExt_1846 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1CD)
        v0_1847 <= v0_1847 & ~maskExt_1847 | maskExt_1847 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1CE)
        v0_1848 <= v0_1848 & ~maskExt_1848 | maskExt_1848 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1CE)
        v0_1849 <= v0_1849 & ~maskExt_1849 | maskExt_1849 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1CE)
        v0_1850 <= v0_1850 & ~maskExt_1850 | maskExt_1850 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1CE)
        v0_1851 <= v0_1851 & ~maskExt_1851 | maskExt_1851 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1CF)
        v0_1852 <= v0_1852 & ~maskExt_1852 | maskExt_1852 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1CF)
        v0_1853 <= v0_1853 & ~maskExt_1853 | maskExt_1853 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1CF)
        v0_1854 <= v0_1854 & ~maskExt_1854 | maskExt_1854 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1CF)
        v0_1855 <= v0_1855 & ~maskExt_1855 | maskExt_1855 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1D0)
        v0_1856 <= v0_1856 & ~maskExt_1856 | maskExt_1856 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1D0)
        v0_1857 <= v0_1857 & ~maskExt_1857 | maskExt_1857 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1D0)
        v0_1858 <= v0_1858 & ~maskExt_1858 | maskExt_1858 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1D0)
        v0_1859 <= v0_1859 & ~maskExt_1859 | maskExt_1859 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1D1)
        v0_1860 <= v0_1860 & ~maskExt_1860 | maskExt_1860 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1D1)
        v0_1861 <= v0_1861 & ~maskExt_1861 | maskExt_1861 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1D1)
        v0_1862 <= v0_1862 & ~maskExt_1862 | maskExt_1862 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1D1)
        v0_1863 <= v0_1863 & ~maskExt_1863 | maskExt_1863 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1D2)
        v0_1864 <= v0_1864 & ~maskExt_1864 | maskExt_1864 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1D2)
        v0_1865 <= v0_1865 & ~maskExt_1865 | maskExt_1865 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1D2)
        v0_1866 <= v0_1866 & ~maskExt_1866 | maskExt_1866 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1D2)
        v0_1867 <= v0_1867 & ~maskExt_1867 | maskExt_1867 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1D3)
        v0_1868 <= v0_1868 & ~maskExt_1868 | maskExt_1868 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1D3)
        v0_1869 <= v0_1869 & ~maskExt_1869 | maskExt_1869 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1D3)
        v0_1870 <= v0_1870 & ~maskExt_1870 | maskExt_1870 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1D3)
        v0_1871 <= v0_1871 & ~maskExt_1871 | maskExt_1871 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1D4)
        v0_1872 <= v0_1872 & ~maskExt_1872 | maskExt_1872 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1D4)
        v0_1873 <= v0_1873 & ~maskExt_1873 | maskExt_1873 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1D4)
        v0_1874 <= v0_1874 & ~maskExt_1874 | maskExt_1874 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1D4)
        v0_1875 <= v0_1875 & ~maskExt_1875 | maskExt_1875 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1D5)
        v0_1876 <= v0_1876 & ~maskExt_1876 | maskExt_1876 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1D5)
        v0_1877 <= v0_1877 & ~maskExt_1877 | maskExt_1877 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1D5)
        v0_1878 <= v0_1878 & ~maskExt_1878 | maskExt_1878 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1D5)
        v0_1879 <= v0_1879 & ~maskExt_1879 | maskExt_1879 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1D6)
        v0_1880 <= v0_1880 & ~maskExt_1880 | maskExt_1880 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1D6)
        v0_1881 <= v0_1881 & ~maskExt_1881 | maskExt_1881 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1D6)
        v0_1882 <= v0_1882 & ~maskExt_1882 | maskExt_1882 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1D6)
        v0_1883 <= v0_1883 & ~maskExt_1883 | maskExt_1883 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1D7)
        v0_1884 <= v0_1884 & ~maskExt_1884 | maskExt_1884 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1D7)
        v0_1885 <= v0_1885 & ~maskExt_1885 | maskExt_1885 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1D7)
        v0_1886 <= v0_1886 & ~maskExt_1886 | maskExt_1886 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1D7)
        v0_1887 <= v0_1887 & ~maskExt_1887 | maskExt_1887 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1D8)
        v0_1888 <= v0_1888 & ~maskExt_1888 | maskExt_1888 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1D8)
        v0_1889 <= v0_1889 & ~maskExt_1889 | maskExt_1889 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1D8)
        v0_1890 <= v0_1890 & ~maskExt_1890 | maskExt_1890 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1D8)
        v0_1891 <= v0_1891 & ~maskExt_1891 | maskExt_1891 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1D9)
        v0_1892 <= v0_1892 & ~maskExt_1892 | maskExt_1892 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1D9)
        v0_1893 <= v0_1893 & ~maskExt_1893 | maskExt_1893 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1D9)
        v0_1894 <= v0_1894 & ~maskExt_1894 | maskExt_1894 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1D9)
        v0_1895 <= v0_1895 & ~maskExt_1895 | maskExt_1895 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1DA)
        v0_1896 <= v0_1896 & ~maskExt_1896 | maskExt_1896 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1DA)
        v0_1897 <= v0_1897 & ~maskExt_1897 | maskExt_1897 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1DA)
        v0_1898 <= v0_1898 & ~maskExt_1898 | maskExt_1898 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1DA)
        v0_1899 <= v0_1899 & ~maskExt_1899 | maskExt_1899 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1DB)
        v0_1900 <= v0_1900 & ~maskExt_1900 | maskExt_1900 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1DB)
        v0_1901 <= v0_1901 & ~maskExt_1901 | maskExt_1901 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1DB)
        v0_1902 <= v0_1902 & ~maskExt_1902 | maskExt_1902 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1DB)
        v0_1903 <= v0_1903 & ~maskExt_1903 | maskExt_1903 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1DC)
        v0_1904 <= v0_1904 & ~maskExt_1904 | maskExt_1904 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1DC)
        v0_1905 <= v0_1905 & ~maskExt_1905 | maskExt_1905 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1DC)
        v0_1906 <= v0_1906 & ~maskExt_1906 | maskExt_1906 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1DC)
        v0_1907 <= v0_1907 & ~maskExt_1907 | maskExt_1907 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1DD)
        v0_1908 <= v0_1908 & ~maskExt_1908 | maskExt_1908 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1DD)
        v0_1909 <= v0_1909 & ~maskExt_1909 | maskExt_1909 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1DD)
        v0_1910 <= v0_1910 & ~maskExt_1910 | maskExt_1910 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1DD)
        v0_1911 <= v0_1911 & ~maskExt_1911 | maskExt_1911 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1DE)
        v0_1912 <= v0_1912 & ~maskExt_1912 | maskExt_1912 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1DE)
        v0_1913 <= v0_1913 & ~maskExt_1913 | maskExt_1913 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1DE)
        v0_1914 <= v0_1914 & ~maskExt_1914 | maskExt_1914 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1DE)
        v0_1915 <= v0_1915 & ~maskExt_1915 | maskExt_1915 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1DF)
        v0_1916 <= v0_1916 & ~maskExt_1916 | maskExt_1916 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1DF)
        v0_1917 <= v0_1917 & ~maskExt_1917 | maskExt_1917 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1DF)
        v0_1918 <= v0_1918 & ~maskExt_1918 | maskExt_1918 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1DF)
        v0_1919 <= v0_1919 & ~maskExt_1919 | maskExt_1919 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1E0)
        v0_1920 <= v0_1920 & ~maskExt_1920 | maskExt_1920 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1E0)
        v0_1921 <= v0_1921 & ~maskExt_1921 | maskExt_1921 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1E0)
        v0_1922 <= v0_1922 & ~maskExt_1922 | maskExt_1922 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1E0)
        v0_1923 <= v0_1923 & ~maskExt_1923 | maskExt_1923 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1E1)
        v0_1924 <= v0_1924 & ~maskExt_1924 | maskExt_1924 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1E1)
        v0_1925 <= v0_1925 & ~maskExt_1925 | maskExt_1925 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1E1)
        v0_1926 <= v0_1926 & ~maskExt_1926 | maskExt_1926 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1E1)
        v0_1927 <= v0_1927 & ~maskExt_1927 | maskExt_1927 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1E2)
        v0_1928 <= v0_1928 & ~maskExt_1928 | maskExt_1928 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1E2)
        v0_1929 <= v0_1929 & ~maskExt_1929 | maskExt_1929 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1E2)
        v0_1930 <= v0_1930 & ~maskExt_1930 | maskExt_1930 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1E2)
        v0_1931 <= v0_1931 & ~maskExt_1931 | maskExt_1931 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1E3)
        v0_1932 <= v0_1932 & ~maskExt_1932 | maskExt_1932 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1E3)
        v0_1933 <= v0_1933 & ~maskExt_1933 | maskExt_1933 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1E3)
        v0_1934 <= v0_1934 & ~maskExt_1934 | maskExt_1934 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1E3)
        v0_1935 <= v0_1935 & ~maskExt_1935 | maskExt_1935 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1E4)
        v0_1936 <= v0_1936 & ~maskExt_1936 | maskExt_1936 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1E4)
        v0_1937 <= v0_1937 & ~maskExt_1937 | maskExt_1937 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1E4)
        v0_1938 <= v0_1938 & ~maskExt_1938 | maskExt_1938 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1E4)
        v0_1939 <= v0_1939 & ~maskExt_1939 | maskExt_1939 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1E5)
        v0_1940 <= v0_1940 & ~maskExt_1940 | maskExt_1940 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1E5)
        v0_1941 <= v0_1941 & ~maskExt_1941 | maskExt_1941 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1E5)
        v0_1942 <= v0_1942 & ~maskExt_1942 | maskExt_1942 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1E5)
        v0_1943 <= v0_1943 & ~maskExt_1943 | maskExt_1943 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1E6)
        v0_1944 <= v0_1944 & ~maskExt_1944 | maskExt_1944 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1E6)
        v0_1945 <= v0_1945 & ~maskExt_1945 | maskExt_1945 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1E6)
        v0_1946 <= v0_1946 & ~maskExt_1946 | maskExt_1946 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1E6)
        v0_1947 <= v0_1947 & ~maskExt_1947 | maskExt_1947 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1E7)
        v0_1948 <= v0_1948 & ~maskExt_1948 | maskExt_1948 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1E7)
        v0_1949 <= v0_1949 & ~maskExt_1949 | maskExt_1949 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1E7)
        v0_1950 <= v0_1950 & ~maskExt_1950 | maskExt_1950 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1E7)
        v0_1951 <= v0_1951 & ~maskExt_1951 | maskExt_1951 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1E8)
        v0_1952 <= v0_1952 & ~maskExt_1952 | maskExt_1952 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1E8)
        v0_1953 <= v0_1953 & ~maskExt_1953 | maskExt_1953 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1E8)
        v0_1954 <= v0_1954 & ~maskExt_1954 | maskExt_1954 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1E8)
        v0_1955 <= v0_1955 & ~maskExt_1955 | maskExt_1955 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1E9)
        v0_1956 <= v0_1956 & ~maskExt_1956 | maskExt_1956 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1E9)
        v0_1957 <= v0_1957 & ~maskExt_1957 | maskExt_1957 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1E9)
        v0_1958 <= v0_1958 & ~maskExt_1958 | maskExt_1958 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1E9)
        v0_1959 <= v0_1959 & ~maskExt_1959 | maskExt_1959 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1EA)
        v0_1960 <= v0_1960 & ~maskExt_1960 | maskExt_1960 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1EA)
        v0_1961 <= v0_1961 & ~maskExt_1961 | maskExt_1961 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1EA)
        v0_1962 <= v0_1962 & ~maskExt_1962 | maskExt_1962 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1EA)
        v0_1963 <= v0_1963 & ~maskExt_1963 | maskExt_1963 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1EB)
        v0_1964 <= v0_1964 & ~maskExt_1964 | maskExt_1964 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1EB)
        v0_1965 <= v0_1965 & ~maskExt_1965 | maskExt_1965 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1EB)
        v0_1966 <= v0_1966 & ~maskExt_1966 | maskExt_1966 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1EB)
        v0_1967 <= v0_1967 & ~maskExt_1967 | maskExt_1967 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1EC)
        v0_1968 <= v0_1968 & ~maskExt_1968 | maskExt_1968 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1EC)
        v0_1969 <= v0_1969 & ~maskExt_1969 | maskExt_1969 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1EC)
        v0_1970 <= v0_1970 & ~maskExt_1970 | maskExt_1970 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1EC)
        v0_1971 <= v0_1971 & ~maskExt_1971 | maskExt_1971 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1ED)
        v0_1972 <= v0_1972 & ~maskExt_1972 | maskExt_1972 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1ED)
        v0_1973 <= v0_1973 & ~maskExt_1973 | maskExt_1973 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1ED)
        v0_1974 <= v0_1974 & ~maskExt_1974 | maskExt_1974 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1ED)
        v0_1975 <= v0_1975 & ~maskExt_1975 | maskExt_1975 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1EE)
        v0_1976 <= v0_1976 & ~maskExt_1976 | maskExt_1976 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1EE)
        v0_1977 <= v0_1977 & ~maskExt_1977 | maskExt_1977 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1EE)
        v0_1978 <= v0_1978 & ~maskExt_1978 | maskExt_1978 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1EE)
        v0_1979 <= v0_1979 & ~maskExt_1979 | maskExt_1979 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1EF)
        v0_1980 <= v0_1980 & ~maskExt_1980 | maskExt_1980 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1EF)
        v0_1981 <= v0_1981 & ~maskExt_1981 | maskExt_1981 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1EF)
        v0_1982 <= v0_1982 & ~maskExt_1982 | maskExt_1982 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1EF)
        v0_1983 <= v0_1983 & ~maskExt_1983 | maskExt_1983 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1F0)
        v0_1984 <= v0_1984 & ~maskExt_1984 | maskExt_1984 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1F0)
        v0_1985 <= v0_1985 & ~maskExt_1985 | maskExt_1985 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1F0)
        v0_1986 <= v0_1986 & ~maskExt_1986 | maskExt_1986 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1F0)
        v0_1987 <= v0_1987 & ~maskExt_1987 | maskExt_1987 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1F1)
        v0_1988 <= v0_1988 & ~maskExt_1988 | maskExt_1988 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1F1)
        v0_1989 <= v0_1989 & ~maskExt_1989 | maskExt_1989 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1F1)
        v0_1990 <= v0_1990 & ~maskExt_1990 | maskExt_1990 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1F1)
        v0_1991 <= v0_1991 & ~maskExt_1991 | maskExt_1991 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1F2)
        v0_1992 <= v0_1992 & ~maskExt_1992 | maskExt_1992 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1F2)
        v0_1993 <= v0_1993 & ~maskExt_1993 | maskExt_1993 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1F2)
        v0_1994 <= v0_1994 & ~maskExt_1994 | maskExt_1994 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1F2)
        v0_1995 <= v0_1995 & ~maskExt_1995 | maskExt_1995 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1F3)
        v0_1996 <= v0_1996 & ~maskExt_1996 | maskExt_1996 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1F3)
        v0_1997 <= v0_1997 & ~maskExt_1997 | maskExt_1997 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1F3)
        v0_1998 <= v0_1998 & ~maskExt_1998 | maskExt_1998 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1F3)
        v0_1999 <= v0_1999 & ~maskExt_1999 | maskExt_1999 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1F4)
        v0_2000 <= v0_2000 & ~maskExt_2000 | maskExt_2000 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1F4)
        v0_2001 <= v0_2001 & ~maskExt_2001 | maskExt_2001 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1F4)
        v0_2002 <= v0_2002 & ~maskExt_2002 | maskExt_2002 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1F4)
        v0_2003 <= v0_2003 & ~maskExt_2003 | maskExt_2003 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1F5)
        v0_2004 <= v0_2004 & ~maskExt_2004 | maskExt_2004 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1F5)
        v0_2005 <= v0_2005 & ~maskExt_2005 | maskExt_2005 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1F5)
        v0_2006 <= v0_2006 & ~maskExt_2006 | maskExt_2006 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1F5)
        v0_2007 <= v0_2007 & ~maskExt_2007 | maskExt_2007 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1F6)
        v0_2008 <= v0_2008 & ~maskExt_2008 | maskExt_2008 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1F6)
        v0_2009 <= v0_2009 & ~maskExt_2009 | maskExt_2009 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1F6)
        v0_2010 <= v0_2010 & ~maskExt_2010 | maskExt_2010 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1F6)
        v0_2011 <= v0_2011 & ~maskExt_2011 | maskExt_2011 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1F7)
        v0_2012 <= v0_2012 & ~maskExt_2012 | maskExt_2012 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1F7)
        v0_2013 <= v0_2013 & ~maskExt_2013 | maskExt_2013 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1F7)
        v0_2014 <= v0_2014 & ~maskExt_2014 | maskExt_2014 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1F7)
        v0_2015 <= v0_2015 & ~maskExt_2015 | maskExt_2015 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1F8)
        v0_2016 <= v0_2016 & ~maskExt_2016 | maskExt_2016 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1F8)
        v0_2017 <= v0_2017 & ~maskExt_2017 | maskExt_2017 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1F8)
        v0_2018 <= v0_2018 & ~maskExt_2018 | maskExt_2018 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1F8)
        v0_2019 <= v0_2019 & ~maskExt_2019 | maskExt_2019 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1F9)
        v0_2020 <= v0_2020 & ~maskExt_2020 | maskExt_2020 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1F9)
        v0_2021 <= v0_2021 & ~maskExt_2021 | maskExt_2021 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1F9)
        v0_2022 <= v0_2022 & ~maskExt_2022 | maskExt_2022 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1F9)
        v0_2023 <= v0_2023 & ~maskExt_2023 | maskExt_2023 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1FA)
        v0_2024 <= v0_2024 & ~maskExt_2024 | maskExt_2024 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1FA)
        v0_2025 <= v0_2025 & ~maskExt_2025 | maskExt_2025 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1FA)
        v0_2026 <= v0_2026 & ~maskExt_2026 | maskExt_2026 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1FA)
        v0_2027 <= v0_2027 & ~maskExt_2027 | maskExt_2027 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1FB)
        v0_2028 <= v0_2028 & ~maskExt_2028 | maskExt_2028 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1FB)
        v0_2029 <= v0_2029 & ~maskExt_2029 | maskExt_2029 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1FB)
        v0_2030 <= v0_2030 & ~maskExt_2030 | maskExt_2030 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1FB)
        v0_2031 <= v0_2031 & ~maskExt_2031 | maskExt_2031 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1FC)
        v0_2032 <= v0_2032 & ~maskExt_2032 | maskExt_2032 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1FC)
        v0_2033 <= v0_2033 & ~maskExt_2033 | maskExt_2033 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1FC)
        v0_2034 <= v0_2034 & ~maskExt_2034 | maskExt_2034 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1FC)
        v0_2035 <= v0_2035 & ~maskExt_2035 | maskExt_2035 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1FD)
        v0_2036 <= v0_2036 & ~maskExt_2036 | maskExt_2036 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1FD)
        v0_2037 <= v0_2037 & ~maskExt_2037 | maskExt_2037 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1FD)
        v0_2038 <= v0_2038 & ~maskExt_2038 | maskExt_2038 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1FD)
        v0_2039 <= v0_2039 & ~maskExt_2039 | maskExt_2039 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 9'h1FE)
        v0_2040 <= v0_2040 & ~maskExt_2040 | maskExt_2040 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 9'h1FE)
        v0_2041 <= v0_2041 & ~maskExt_2041 | maskExt_2041 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 9'h1FE)
        v0_2042 <= v0_2042 & ~maskExt_2042 | maskExt_2042 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 9'h1FE)
        v0_2043 <= v0_2043 & ~maskExt_2043 | maskExt_2043 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & (&v0UpdateVec_0_bits_offset))
        v0_2044 <= v0_2044 & ~maskExt_2044 | maskExt_2044 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & (&v0UpdateVec_1_bits_offset))
        v0_2045 <= v0_2045 & ~maskExt_2045 | maskExt_2045 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & (&v0UpdateVec_2_bits_offset))
        v0_2046 <= v0_2046 & ~maskExt_2046 | maskExt_2046 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & (&v0UpdateVec_3_bits_offset))
        v0_2047 <= v0_2047 & ~maskExt_2047 | maskExt_2047 & v0UpdateVec_3_bits_data;
      if (queueEnq[0] ^ queueDeq[0])
        queueCount_0 <= queueCount_0 + counterUpdate;
      if (queueEnq[1] ^ queueDeq[1])
        queueCount_1 <= queueCount_1 + counterUpdate_1;
      if (queueEnq[2] ^ queueDeq[2])
        queueCount_2 <= queueCount_2 + counterUpdate_2;
      if (queueEnq[3] ^ queueDeq[3])
        queueCount_3 <= queueCount_3 + counterUpdate_3;
      if (queueEnq[4] ^ queueDeq[4])
        queueCount_4 <= queueCount_4 + counterUpdate_4;
      if (queueEnq[5] ^ queueDeq[5])
        queueCount_5 <= queueCount_5 + counterUpdate_5;
      if (queueEnq[6] ^ queueDeq[6])
        queueCount_6 <= queueCount_6 + counterUpdate_6;
      if (queueEnq[7] ^ queueDeq[7])
        queueCount_7 <= queueCount_7 + counterUpdate_7;
      if (queueEnq_1[0] ^ queueDeq_1[0])
        queueCount_0_1 <= queueCount_0_1 + counterUpdate_8;
      if (queueEnq_1[1] ^ queueDeq_1[1])
        queueCount_1_1 <= queueCount_1_1 + counterUpdate_9;
      if (queueEnq_1[2] ^ queueDeq_1[2])
        queueCount_2_1 <= queueCount_2_1 + counterUpdate_10;
      if (queueEnq_1[3] ^ queueDeq_1[3])
        queueCount_3_1 <= queueCount_3_1 + counterUpdate_11;
      if (queueEnq_1[4] ^ queueDeq_1[4])
        queueCount_4_1 <= queueCount_4_1 + counterUpdate_12;
      if (queueEnq_1[5] ^ queueDeq_1[5])
        queueCount_5_1 <= queueCount_5_1 + counterUpdate_13;
      if (queueEnq_1[6] ^ queueDeq_1[6])
        queueCount_6_1 <= queueCount_6_1 + counterUpdate_14;
      if (queueEnq_1[7] ^ queueDeq_1[7])
        queueCount_7_1 <= queueCount_7_1 + counterUpdate_15;
      if (queueEnq_2[0] ^ queueDeq_2[0])
        queueCount_0_2 <= queueCount_0_2 + counterUpdate_16;
      if (queueEnq_2[1] ^ queueDeq_2[1])
        queueCount_1_2 <= queueCount_1_2 + counterUpdate_17;
      if (queueEnq_2[2] ^ queueDeq_2[2])
        queueCount_2_2 <= queueCount_2_2 + counterUpdate_18;
      if (queueEnq_2[3] ^ queueDeq_2[3])
        queueCount_3_2 <= queueCount_3_2 + counterUpdate_19;
      if (queueEnq_2[4] ^ queueDeq_2[4])
        queueCount_4_2 <= queueCount_4_2 + counterUpdate_20;
      if (queueEnq_2[5] ^ queueDeq_2[5])
        queueCount_5_2 <= queueCount_5_2 + counterUpdate_21;
      if (queueEnq_2[6] ^ queueDeq_2[6])
        queueCount_6_2 <= queueCount_6_2 + counterUpdate_22;
      if (queueEnq_2[7] ^ queueDeq_2[7])
        queueCount_7_2 <= queueCount_7_2 + counterUpdate_23;
      if (queueEnq_3[0] ^ queueDeq_3[0])
        queueCount_0_3 <= queueCount_0_3 + counterUpdate_24;
      if (queueEnq_3[1] ^ queueDeq_3[1])
        queueCount_1_3 <= queueCount_1_3 + counterUpdate_25;
      if (queueEnq_3[2] ^ queueDeq_3[2])
        queueCount_2_3 <= queueCount_2_3 + counterUpdate_26;
      if (queueEnq_3[3] ^ queueDeq_3[3])
        queueCount_3_3 <= queueCount_3_3 + counterUpdate_27;
      if (queueEnq_3[4] ^ queueDeq_3[4])
        queueCount_4_3 <= queueCount_4_3 + counterUpdate_28;
      if (queueEnq_3[5] ^ queueDeq_3[5])
        queueCount_5_3 <= queueCount_5_3 + counterUpdate_29;
      if (queueEnq_3[6] ^ queueDeq_3[6])
        queueCount_6_3 <= queueCount_6_3 + counterUpdate_30;
      if (queueEnq_3[7] ^ queueDeq_3[7])
        queueCount_7_3 <= queueCount_7_3 + counterUpdate_31;
    end
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:2054];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [11:0] i = 12'h0; i < 12'h807; i += 12'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        v0_0 = _RANDOM[12'h0];
        v0_1 = _RANDOM[12'h1];
        v0_2 = _RANDOM[12'h2];
        v0_3 = _RANDOM[12'h3];
        v0_4 = _RANDOM[12'h4];
        v0_5 = _RANDOM[12'h5];
        v0_6 = _RANDOM[12'h6];
        v0_7 = _RANDOM[12'h7];
        v0_8 = _RANDOM[12'h8];
        v0_9 = _RANDOM[12'h9];
        v0_10 = _RANDOM[12'hA];
        v0_11 = _RANDOM[12'hB];
        v0_12 = _RANDOM[12'hC];
        v0_13 = _RANDOM[12'hD];
        v0_14 = _RANDOM[12'hE];
        v0_15 = _RANDOM[12'hF];
        v0_16 = _RANDOM[12'h10];
        v0_17 = _RANDOM[12'h11];
        v0_18 = _RANDOM[12'h12];
        v0_19 = _RANDOM[12'h13];
        v0_20 = _RANDOM[12'h14];
        v0_21 = _RANDOM[12'h15];
        v0_22 = _RANDOM[12'h16];
        v0_23 = _RANDOM[12'h17];
        v0_24 = _RANDOM[12'h18];
        v0_25 = _RANDOM[12'h19];
        v0_26 = _RANDOM[12'h1A];
        v0_27 = _RANDOM[12'h1B];
        v0_28 = _RANDOM[12'h1C];
        v0_29 = _RANDOM[12'h1D];
        v0_30 = _RANDOM[12'h1E];
        v0_31 = _RANDOM[12'h1F];
        v0_32 = _RANDOM[12'h20];
        v0_33 = _RANDOM[12'h21];
        v0_34 = _RANDOM[12'h22];
        v0_35 = _RANDOM[12'h23];
        v0_36 = _RANDOM[12'h24];
        v0_37 = _RANDOM[12'h25];
        v0_38 = _RANDOM[12'h26];
        v0_39 = _RANDOM[12'h27];
        v0_40 = _RANDOM[12'h28];
        v0_41 = _RANDOM[12'h29];
        v0_42 = _RANDOM[12'h2A];
        v0_43 = _RANDOM[12'h2B];
        v0_44 = _RANDOM[12'h2C];
        v0_45 = _RANDOM[12'h2D];
        v0_46 = _RANDOM[12'h2E];
        v0_47 = _RANDOM[12'h2F];
        v0_48 = _RANDOM[12'h30];
        v0_49 = _RANDOM[12'h31];
        v0_50 = _RANDOM[12'h32];
        v0_51 = _RANDOM[12'h33];
        v0_52 = _RANDOM[12'h34];
        v0_53 = _RANDOM[12'h35];
        v0_54 = _RANDOM[12'h36];
        v0_55 = _RANDOM[12'h37];
        v0_56 = _RANDOM[12'h38];
        v0_57 = _RANDOM[12'h39];
        v0_58 = _RANDOM[12'h3A];
        v0_59 = _RANDOM[12'h3B];
        v0_60 = _RANDOM[12'h3C];
        v0_61 = _RANDOM[12'h3D];
        v0_62 = _RANDOM[12'h3E];
        v0_63 = _RANDOM[12'h3F];
        v0_64 = _RANDOM[12'h40];
        v0_65 = _RANDOM[12'h41];
        v0_66 = _RANDOM[12'h42];
        v0_67 = _RANDOM[12'h43];
        v0_68 = _RANDOM[12'h44];
        v0_69 = _RANDOM[12'h45];
        v0_70 = _RANDOM[12'h46];
        v0_71 = _RANDOM[12'h47];
        v0_72 = _RANDOM[12'h48];
        v0_73 = _RANDOM[12'h49];
        v0_74 = _RANDOM[12'h4A];
        v0_75 = _RANDOM[12'h4B];
        v0_76 = _RANDOM[12'h4C];
        v0_77 = _RANDOM[12'h4D];
        v0_78 = _RANDOM[12'h4E];
        v0_79 = _RANDOM[12'h4F];
        v0_80 = _RANDOM[12'h50];
        v0_81 = _RANDOM[12'h51];
        v0_82 = _RANDOM[12'h52];
        v0_83 = _RANDOM[12'h53];
        v0_84 = _RANDOM[12'h54];
        v0_85 = _RANDOM[12'h55];
        v0_86 = _RANDOM[12'h56];
        v0_87 = _RANDOM[12'h57];
        v0_88 = _RANDOM[12'h58];
        v0_89 = _RANDOM[12'h59];
        v0_90 = _RANDOM[12'h5A];
        v0_91 = _RANDOM[12'h5B];
        v0_92 = _RANDOM[12'h5C];
        v0_93 = _RANDOM[12'h5D];
        v0_94 = _RANDOM[12'h5E];
        v0_95 = _RANDOM[12'h5F];
        v0_96 = _RANDOM[12'h60];
        v0_97 = _RANDOM[12'h61];
        v0_98 = _RANDOM[12'h62];
        v0_99 = _RANDOM[12'h63];
        v0_100 = _RANDOM[12'h64];
        v0_101 = _RANDOM[12'h65];
        v0_102 = _RANDOM[12'h66];
        v0_103 = _RANDOM[12'h67];
        v0_104 = _RANDOM[12'h68];
        v0_105 = _RANDOM[12'h69];
        v0_106 = _RANDOM[12'h6A];
        v0_107 = _RANDOM[12'h6B];
        v0_108 = _RANDOM[12'h6C];
        v0_109 = _RANDOM[12'h6D];
        v0_110 = _RANDOM[12'h6E];
        v0_111 = _RANDOM[12'h6F];
        v0_112 = _RANDOM[12'h70];
        v0_113 = _RANDOM[12'h71];
        v0_114 = _RANDOM[12'h72];
        v0_115 = _RANDOM[12'h73];
        v0_116 = _RANDOM[12'h74];
        v0_117 = _RANDOM[12'h75];
        v0_118 = _RANDOM[12'h76];
        v0_119 = _RANDOM[12'h77];
        v0_120 = _RANDOM[12'h78];
        v0_121 = _RANDOM[12'h79];
        v0_122 = _RANDOM[12'h7A];
        v0_123 = _RANDOM[12'h7B];
        v0_124 = _RANDOM[12'h7C];
        v0_125 = _RANDOM[12'h7D];
        v0_126 = _RANDOM[12'h7E];
        v0_127 = _RANDOM[12'h7F];
        v0_128 = _RANDOM[12'h80];
        v0_129 = _RANDOM[12'h81];
        v0_130 = _RANDOM[12'h82];
        v0_131 = _RANDOM[12'h83];
        v0_132 = _RANDOM[12'h84];
        v0_133 = _RANDOM[12'h85];
        v0_134 = _RANDOM[12'h86];
        v0_135 = _RANDOM[12'h87];
        v0_136 = _RANDOM[12'h88];
        v0_137 = _RANDOM[12'h89];
        v0_138 = _RANDOM[12'h8A];
        v0_139 = _RANDOM[12'h8B];
        v0_140 = _RANDOM[12'h8C];
        v0_141 = _RANDOM[12'h8D];
        v0_142 = _RANDOM[12'h8E];
        v0_143 = _RANDOM[12'h8F];
        v0_144 = _RANDOM[12'h90];
        v0_145 = _RANDOM[12'h91];
        v0_146 = _RANDOM[12'h92];
        v0_147 = _RANDOM[12'h93];
        v0_148 = _RANDOM[12'h94];
        v0_149 = _RANDOM[12'h95];
        v0_150 = _RANDOM[12'h96];
        v0_151 = _RANDOM[12'h97];
        v0_152 = _RANDOM[12'h98];
        v0_153 = _RANDOM[12'h99];
        v0_154 = _RANDOM[12'h9A];
        v0_155 = _RANDOM[12'h9B];
        v0_156 = _RANDOM[12'h9C];
        v0_157 = _RANDOM[12'h9D];
        v0_158 = _RANDOM[12'h9E];
        v0_159 = _RANDOM[12'h9F];
        v0_160 = _RANDOM[12'hA0];
        v0_161 = _RANDOM[12'hA1];
        v0_162 = _RANDOM[12'hA2];
        v0_163 = _RANDOM[12'hA3];
        v0_164 = _RANDOM[12'hA4];
        v0_165 = _RANDOM[12'hA5];
        v0_166 = _RANDOM[12'hA6];
        v0_167 = _RANDOM[12'hA7];
        v0_168 = _RANDOM[12'hA8];
        v0_169 = _RANDOM[12'hA9];
        v0_170 = _RANDOM[12'hAA];
        v0_171 = _RANDOM[12'hAB];
        v0_172 = _RANDOM[12'hAC];
        v0_173 = _RANDOM[12'hAD];
        v0_174 = _RANDOM[12'hAE];
        v0_175 = _RANDOM[12'hAF];
        v0_176 = _RANDOM[12'hB0];
        v0_177 = _RANDOM[12'hB1];
        v0_178 = _RANDOM[12'hB2];
        v0_179 = _RANDOM[12'hB3];
        v0_180 = _RANDOM[12'hB4];
        v0_181 = _RANDOM[12'hB5];
        v0_182 = _RANDOM[12'hB6];
        v0_183 = _RANDOM[12'hB7];
        v0_184 = _RANDOM[12'hB8];
        v0_185 = _RANDOM[12'hB9];
        v0_186 = _RANDOM[12'hBA];
        v0_187 = _RANDOM[12'hBB];
        v0_188 = _RANDOM[12'hBC];
        v0_189 = _RANDOM[12'hBD];
        v0_190 = _RANDOM[12'hBE];
        v0_191 = _RANDOM[12'hBF];
        v0_192 = _RANDOM[12'hC0];
        v0_193 = _RANDOM[12'hC1];
        v0_194 = _RANDOM[12'hC2];
        v0_195 = _RANDOM[12'hC3];
        v0_196 = _RANDOM[12'hC4];
        v0_197 = _RANDOM[12'hC5];
        v0_198 = _RANDOM[12'hC6];
        v0_199 = _RANDOM[12'hC7];
        v0_200 = _RANDOM[12'hC8];
        v0_201 = _RANDOM[12'hC9];
        v0_202 = _RANDOM[12'hCA];
        v0_203 = _RANDOM[12'hCB];
        v0_204 = _RANDOM[12'hCC];
        v0_205 = _RANDOM[12'hCD];
        v0_206 = _RANDOM[12'hCE];
        v0_207 = _RANDOM[12'hCF];
        v0_208 = _RANDOM[12'hD0];
        v0_209 = _RANDOM[12'hD1];
        v0_210 = _RANDOM[12'hD2];
        v0_211 = _RANDOM[12'hD3];
        v0_212 = _RANDOM[12'hD4];
        v0_213 = _RANDOM[12'hD5];
        v0_214 = _RANDOM[12'hD6];
        v0_215 = _RANDOM[12'hD7];
        v0_216 = _RANDOM[12'hD8];
        v0_217 = _RANDOM[12'hD9];
        v0_218 = _RANDOM[12'hDA];
        v0_219 = _RANDOM[12'hDB];
        v0_220 = _RANDOM[12'hDC];
        v0_221 = _RANDOM[12'hDD];
        v0_222 = _RANDOM[12'hDE];
        v0_223 = _RANDOM[12'hDF];
        v0_224 = _RANDOM[12'hE0];
        v0_225 = _RANDOM[12'hE1];
        v0_226 = _RANDOM[12'hE2];
        v0_227 = _RANDOM[12'hE3];
        v0_228 = _RANDOM[12'hE4];
        v0_229 = _RANDOM[12'hE5];
        v0_230 = _RANDOM[12'hE6];
        v0_231 = _RANDOM[12'hE7];
        v0_232 = _RANDOM[12'hE8];
        v0_233 = _RANDOM[12'hE9];
        v0_234 = _RANDOM[12'hEA];
        v0_235 = _RANDOM[12'hEB];
        v0_236 = _RANDOM[12'hEC];
        v0_237 = _RANDOM[12'hED];
        v0_238 = _RANDOM[12'hEE];
        v0_239 = _RANDOM[12'hEF];
        v0_240 = _RANDOM[12'hF0];
        v0_241 = _RANDOM[12'hF1];
        v0_242 = _RANDOM[12'hF2];
        v0_243 = _RANDOM[12'hF3];
        v0_244 = _RANDOM[12'hF4];
        v0_245 = _RANDOM[12'hF5];
        v0_246 = _RANDOM[12'hF6];
        v0_247 = _RANDOM[12'hF7];
        v0_248 = _RANDOM[12'hF8];
        v0_249 = _RANDOM[12'hF9];
        v0_250 = _RANDOM[12'hFA];
        v0_251 = _RANDOM[12'hFB];
        v0_252 = _RANDOM[12'hFC];
        v0_253 = _RANDOM[12'hFD];
        v0_254 = _RANDOM[12'hFE];
        v0_255 = _RANDOM[12'hFF];
        v0_256 = _RANDOM[12'h100];
        v0_257 = _RANDOM[12'h101];
        v0_258 = _RANDOM[12'h102];
        v0_259 = _RANDOM[12'h103];
        v0_260 = _RANDOM[12'h104];
        v0_261 = _RANDOM[12'h105];
        v0_262 = _RANDOM[12'h106];
        v0_263 = _RANDOM[12'h107];
        v0_264 = _RANDOM[12'h108];
        v0_265 = _RANDOM[12'h109];
        v0_266 = _RANDOM[12'h10A];
        v0_267 = _RANDOM[12'h10B];
        v0_268 = _RANDOM[12'h10C];
        v0_269 = _RANDOM[12'h10D];
        v0_270 = _RANDOM[12'h10E];
        v0_271 = _RANDOM[12'h10F];
        v0_272 = _RANDOM[12'h110];
        v0_273 = _RANDOM[12'h111];
        v0_274 = _RANDOM[12'h112];
        v0_275 = _RANDOM[12'h113];
        v0_276 = _RANDOM[12'h114];
        v0_277 = _RANDOM[12'h115];
        v0_278 = _RANDOM[12'h116];
        v0_279 = _RANDOM[12'h117];
        v0_280 = _RANDOM[12'h118];
        v0_281 = _RANDOM[12'h119];
        v0_282 = _RANDOM[12'h11A];
        v0_283 = _RANDOM[12'h11B];
        v0_284 = _RANDOM[12'h11C];
        v0_285 = _RANDOM[12'h11D];
        v0_286 = _RANDOM[12'h11E];
        v0_287 = _RANDOM[12'h11F];
        v0_288 = _RANDOM[12'h120];
        v0_289 = _RANDOM[12'h121];
        v0_290 = _RANDOM[12'h122];
        v0_291 = _RANDOM[12'h123];
        v0_292 = _RANDOM[12'h124];
        v0_293 = _RANDOM[12'h125];
        v0_294 = _RANDOM[12'h126];
        v0_295 = _RANDOM[12'h127];
        v0_296 = _RANDOM[12'h128];
        v0_297 = _RANDOM[12'h129];
        v0_298 = _RANDOM[12'h12A];
        v0_299 = _RANDOM[12'h12B];
        v0_300 = _RANDOM[12'h12C];
        v0_301 = _RANDOM[12'h12D];
        v0_302 = _RANDOM[12'h12E];
        v0_303 = _RANDOM[12'h12F];
        v0_304 = _RANDOM[12'h130];
        v0_305 = _RANDOM[12'h131];
        v0_306 = _RANDOM[12'h132];
        v0_307 = _RANDOM[12'h133];
        v0_308 = _RANDOM[12'h134];
        v0_309 = _RANDOM[12'h135];
        v0_310 = _RANDOM[12'h136];
        v0_311 = _RANDOM[12'h137];
        v0_312 = _RANDOM[12'h138];
        v0_313 = _RANDOM[12'h139];
        v0_314 = _RANDOM[12'h13A];
        v0_315 = _RANDOM[12'h13B];
        v0_316 = _RANDOM[12'h13C];
        v0_317 = _RANDOM[12'h13D];
        v0_318 = _RANDOM[12'h13E];
        v0_319 = _RANDOM[12'h13F];
        v0_320 = _RANDOM[12'h140];
        v0_321 = _RANDOM[12'h141];
        v0_322 = _RANDOM[12'h142];
        v0_323 = _RANDOM[12'h143];
        v0_324 = _RANDOM[12'h144];
        v0_325 = _RANDOM[12'h145];
        v0_326 = _RANDOM[12'h146];
        v0_327 = _RANDOM[12'h147];
        v0_328 = _RANDOM[12'h148];
        v0_329 = _RANDOM[12'h149];
        v0_330 = _RANDOM[12'h14A];
        v0_331 = _RANDOM[12'h14B];
        v0_332 = _RANDOM[12'h14C];
        v0_333 = _RANDOM[12'h14D];
        v0_334 = _RANDOM[12'h14E];
        v0_335 = _RANDOM[12'h14F];
        v0_336 = _RANDOM[12'h150];
        v0_337 = _RANDOM[12'h151];
        v0_338 = _RANDOM[12'h152];
        v0_339 = _RANDOM[12'h153];
        v0_340 = _RANDOM[12'h154];
        v0_341 = _RANDOM[12'h155];
        v0_342 = _RANDOM[12'h156];
        v0_343 = _RANDOM[12'h157];
        v0_344 = _RANDOM[12'h158];
        v0_345 = _RANDOM[12'h159];
        v0_346 = _RANDOM[12'h15A];
        v0_347 = _RANDOM[12'h15B];
        v0_348 = _RANDOM[12'h15C];
        v0_349 = _RANDOM[12'h15D];
        v0_350 = _RANDOM[12'h15E];
        v0_351 = _RANDOM[12'h15F];
        v0_352 = _RANDOM[12'h160];
        v0_353 = _RANDOM[12'h161];
        v0_354 = _RANDOM[12'h162];
        v0_355 = _RANDOM[12'h163];
        v0_356 = _RANDOM[12'h164];
        v0_357 = _RANDOM[12'h165];
        v0_358 = _RANDOM[12'h166];
        v0_359 = _RANDOM[12'h167];
        v0_360 = _RANDOM[12'h168];
        v0_361 = _RANDOM[12'h169];
        v0_362 = _RANDOM[12'h16A];
        v0_363 = _RANDOM[12'h16B];
        v0_364 = _RANDOM[12'h16C];
        v0_365 = _RANDOM[12'h16D];
        v0_366 = _RANDOM[12'h16E];
        v0_367 = _RANDOM[12'h16F];
        v0_368 = _RANDOM[12'h170];
        v0_369 = _RANDOM[12'h171];
        v0_370 = _RANDOM[12'h172];
        v0_371 = _RANDOM[12'h173];
        v0_372 = _RANDOM[12'h174];
        v0_373 = _RANDOM[12'h175];
        v0_374 = _RANDOM[12'h176];
        v0_375 = _RANDOM[12'h177];
        v0_376 = _RANDOM[12'h178];
        v0_377 = _RANDOM[12'h179];
        v0_378 = _RANDOM[12'h17A];
        v0_379 = _RANDOM[12'h17B];
        v0_380 = _RANDOM[12'h17C];
        v0_381 = _RANDOM[12'h17D];
        v0_382 = _RANDOM[12'h17E];
        v0_383 = _RANDOM[12'h17F];
        v0_384 = _RANDOM[12'h180];
        v0_385 = _RANDOM[12'h181];
        v0_386 = _RANDOM[12'h182];
        v0_387 = _RANDOM[12'h183];
        v0_388 = _RANDOM[12'h184];
        v0_389 = _RANDOM[12'h185];
        v0_390 = _RANDOM[12'h186];
        v0_391 = _RANDOM[12'h187];
        v0_392 = _RANDOM[12'h188];
        v0_393 = _RANDOM[12'h189];
        v0_394 = _RANDOM[12'h18A];
        v0_395 = _RANDOM[12'h18B];
        v0_396 = _RANDOM[12'h18C];
        v0_397 = _RANDOM[12'h18D];
        v0_398 = _RANDOM[12'h18E];
        v0_399 = _RANDOM[12'h18F];
        v0_400 = _RANDOM[12'h190];
        v0_401 = _RANDOM[12'h191];
        v0_402 = _RANDOM[12'h192];
        v0_403 = _RANDOM[12'h193];
        v0_404 = _RANDOM[12'h194];
        v0_405 = _RANDOM[12'h195];
        v0_406 = _RANDOM[12'h196];
        v0_407 = _RANDOM[12'h197];
        v0_408 = _RANDOM[12'h198];
        v0_409 = _RANDOM[12'h199];
        v0_410 = _RANDOM[12'h19A];
        v0_411 = _RANDOM[12'h19B];
        v0_412 = _RANDOM[12'h19C];
        v0_413 = _RANDOM[12'h19D];
        v0_414 = _RANDOM[12'h19E];
        v0_415 = _RANDOM[12'h19F];
        v0_416 = _RANDOM[12'h1A0];
        v0_417 = _RANDOM[12'h1A1];
        v0_418 = _RANDOM[12'h1A2];
        v0_419 = _RANDOM[12'h1A3];
        v0_420 = _RANDOM[12'h1A4];
        v0_421 = _RANDOM[12'h1A5];
        v0_422 = _RANDOM[12'h1A6];
        v0_423 = _RANDOM[12'h1A7];
        v0_424 = _RANDOM[12'h1A8];
        v0_425 = _RANDOM[12'h1A9];
        v0_426 = _RANDOM[12'h1AA];
        v0_427 = _RANDOM[12'h1AB];
        v0_428 = _RANDOM[12'h1AC];
        v0_429 = _RANDOM[12'h1AD];
        v0_430 = _RANDOM[12'h1AE];
        v0_431 = _RANDOM[12'h1AF];
        v0_432 = _RANDOM[12'h1B0];
        v0_433 = _RANDOM[12'h1B1];
        v0_434 = _RANDOM[12'h1B2];
        v0_435 = _RANDOM[12'h1B3];
        v0_436 = _RANDOM[12'h1B4];
        v0_437 = _RANDOM[12'h1B5];
        v0_438 = _RANDOM[12'h1B6];
        v0_439 = _RANDOM[12'h1B7];
        v0_440 = _RANDOM[12'h1B8];
        v0_441 = _RANDOM[12'h1B9];
        v0_442 = _RANDOM[12'h1BA];
        v0_443 = _RANDOM[12'h1BB];
        v0_444 = _RANDOM[12'h1BC];
        v0_445 = _RANDOM[12'h1BD];
        v0_446 = _RANDOM[12'h1BE];
        v0_447 = _RANDOM[12'h1BF];
        v0_448 = _RANDOM[12'h1C0];
        v0_449 = _RANDOM[12'h1C1];
        v0_450 = _RANDOM[12'h1C2];
        v0_451 = _RANDOM[12'h1C3];
        v0_452 = _RANDOM[12'h1C4];
        v0_453 = _RANDOM[12'h1C5];
        v0_454 = _RANDOM[12'h1C6];
        v0_455 = _RANDOM[12'h1C7];
        v0_456 = _RANDOM[12'h1C8];
        v0_457 = _RANDOM[12'h1C9];
        v0_458 = _RANDOM[12'h1CA];
        v0_459 = _RANDOM[12'h1CB];
        v0_460 = _RANDOM[12'h1CC];
        v0_461 = _RANDOM[12'h1CD];
        v0_462 = _RANDOM[12'h1CE];
        v0_463 = _RANDOM[12'h1CF];
        v0_464 = _RANDOM[12'h1D0];
        v0_465 = _RANDOM[12'h1D1];
        v0_466 = _RANDOM[12'h1D2];
        v0_467 = _RANDOM[12'h1D3];
        v0_468 = _RANDOM[12'h1D4];
        v0_469 = _RANDOM[12'h1D5];
        v0_470 = _RANDOM[12'h1D6];
        v0_471 = _RANDOM[12'h1D7];
        v0_472 = _RANDOM[12'h1D8];
        v0_473 = _RANDOM[12'h1D9];
        v0_474 = _RANDOM[12'h1DA];
        v0_475 = _RANDOM[12'h1DB];
        v0_476 = _RANDOM[12'h1DC];
        v0_477 = _RANDOM[12'h1DD];
        v0_478 = _RANDOM[12'h1DE];
        v0_479 = _RANDOM[12'h1DF];
        v0_480 = _RANDOM[12'h1E0];
        v0_481 = _RANDOM[12'h1E1];
        v0_482 = _RANDOM[12'h1E2];
        v0_483 = _RANDOM[12'h1E3];
        v0_484 = _RANDOM[12'h1E4];
        v0_485 = _RANDOM[12'h1E5];
        v0_486 = _RANDOM[12'h1E6];
        v0_487 = _RANDOM[12'h1E7];
        v0_488 = _RANDOM[12'h1E8];
        v0_489 = _RANDOM[12'h1E9];
        v0_490 = _RANDOM[12'h1EA];
        v0_491 = _RANDOM[12'h1EB];
        v0_492 = _RANDOM[12'h1EC];
        v0_493 = _RANDOM[12'h1ED];
        v0_494 = _RANDOM[12'h1EE];
        v0_495 = _RANDOM[12'h1EF];
        v0_496 = _RANDOM[12'h1F0];
        v0_497 = _RANDOM[12'h1F1];
        v0_498 = _RANDOM[12'h1F2];
        v0_499 = _RANDOM[12'h1F3];
        v0_500 = _RANDOM[12'h1F4];
        v0_501 = _RANDOM[12'h1F5];
        v0_502 = _RANDOM[12'h1F6];
        v0_503 = _RANDOM[12'h1F7];
        v0_504 = _RANDOM[12'h1F8];
        v0_505 = _RANDOM[12'h1F9];
        v0_506 = _RANDOM[12'h1FA];
        v0_507 = _RANDOM[12'h1FB];
        v0_508 = _RANDOM[12'h1FC];
        v0_509 = _RANDOM[12'h1FD];
        v0_510 = _RANDOM[12'h1FE];
        v0_511 = _RANDOM[12'h1FF];
        v0_512 = _RANDOM[12'h200];
        v0_513 = _RANDOM[12'h201];
        v0_514 = _RANDOM[12'h202];
        v0_515 = _RANDOM[12'h203];
        v0_516 = _RANDOM[12'h204];
        v0_517 = _RANDOM[12'h205];
        v0_518 = _RANDOM[12'h206];
        v0_519 = _RANDOM[12'h207];
        v0_520 = _RANDOM[12'h208];
        v0_521 = _RANDOM[12'h209];
        v0_522 = _RANDOM[12'h20A];
        v0_523 = _RANDOM[12'h20B];
        v0_524 = _RANDOM[12'h20C];
        v0_525 = _RANDOM[12'h20D];
        v0_526 = _RANDOM[12'h20E];
        v0_527 = _RANDOM[12'h20F];
        v0_528 = _RANDOM[12'h210];
        v0_529 = _RANDOM[12'h211];
        v0_530 = _RANDOM[12'h212];
        v0_531 = _RANDOM[12'h213];
        v0_532 = _RANDOM[12'h214];
        v0_533 = _RANDOM[12'h215];
        v0_534 = _RANDOM[12'h216];
        v0_535 = _RANDOM[12'h217];
        v0_536 = _RANDOM[12'h218];
        v0_537 = _RANDOM[12'h219];
        v0_538 = _RANDOM[12'h21A];
        v0_539 = _RANDOM[12'h21B];
        v0_540 = _RANDOM[12'h21C];
        v0_541 = _RANDOM[12'h21D];
        v0_542 = _RANDOM[12'h21E];
        v0_543 = _RANDOM[12'h21F];
        v0_544 = _RANDOM[12'h220];
        v0_545 = _RANDOM[12'h221];
        v0_546 = _RANDOM[12'h222];
        v0_547 = _RANDOM[12'h223];
        v0_548 = _RANDOM[12'h224];
        v0_549 = _RANDOM[12'h225];
        v0_550 = _RANDOM[12'h226];
        v0_551 = _RANDOM[12'h227];
        v0_552 = _RANDOM[12'h228];
        v0_553 = _RANDOM[12'h229];
        v0_554 = _RANDOM[12'h22A];
        v0_555 = _RANDOM[12'h22B];
        v0_556 = _RANDOM[12'h22C];
        v0_557 = _RANDOM[12'h22D];
        v0_558 = _RANDOM[12'h22E];
        v0_559 = _RANDOM[12'h22F];
        v0_560 = _RANDOM[12'h230];
        v0_561 = _RANDOM[12'h231];
        v0_562 = _RANDOM[12'h232];
        v0_563 = _RANDOM[12'h233];
        v0_564 = _RANDOM[12'h234];
        v0_565 = _RANDOM[12'h235];
        v0_566 = _RANDOM[12'h236];
        v0_567 = _RANDOM[12'h237];
        v0_568 = _RANDOM[12'h238];
        v0_569 = _RANDOM[12'h239];
        v0_570 = _RANDOM[12'h23A];
        v0_571 = _RANDOM[12'h23B];
        v0_572 = _RANDOM[12'h23C];
        v0_573 = _RANDOM[12'h23D];
        v0_574 = _RANDOM[12'h23E];
        v0_575 = _RANDOM[12'h23F];
        v0_576 = _RANDOM[12'h240];
        v0_577 = _RANDOM[12'h241];
        v0_578 = _RANDOM[12'h242];
        v0_579 = _RANDOM[12'h243];
        v0_580 = _RANDOM[12'h244];
        v0_581 = _RANDOM[12'h245];
        v0_582 = _RANDOM[12'h246];
        v0_583 = _RANDOM[12'h247];
        v0_584 = _RANDOM[12'h248];
        v0_585 = _RANDOM[12'h249];
        v0_586 = _RANDOM[12'h24A];
        v0_587 = _RANDOM[12'h24B];
        v0_588 = _RANDOM[12'h24C];
        v0_589 = _RANDOM[12'h24D];
        v0_590 = _RANDOM[12'h24E];
        v0_591 = _RANDOM[12'h24F];
        v0_592 = _RANDOM[12'h250];
        v0_593 = _RANDOM[12'h251];
        v0_594 = _RANDOM[12'h252];
        v0_595 = _RANDOM[12'h253];
        v0_596 = _RANDOM[12'h254];
        v0_597 = _RANDOM[12'h255];
        v0_598 = _RANDOM[12'h256];
        v0_599 = _RANDOM[12'h257];
        v0_600 = _RANDOM[12'h258];
        v0_601 = _RANDOM[12'h259];
        v0_602 = _RANDOM[12'h25A];
        v0_603 = _RANDOM[12'h25B];
        v0_604 = _RANDOM[12'h25C];
        v0_605 = _RANDOM[12'h25D];
        v0_606 = _RANDOM[12'h25E];
        v0_607 = _RANDOM[12'h25F];
        v0_608 = _RANDOM[12'h260];
        v0_609 = _RANDOM[12'h261];
        v0_610 = _RANDOM[12'h262];
        v0_611 = _RANDOM[12'h263];
        v0_612 = _RANDOM[12'h264];
        v0_613 = _RANDOM[12'h265];
        v0_614 = _RANDOM[12'h266];
        v0_615 = _RANDOM[12'h267];
        v0_616 = _RANDOM[12'h268];
        v0_617 = _RANDOM[12'h269];
        v0_618 = _RANDOM[12'h26A];
        v0_619 = _RANDOM[12'h26B];
        v0_620 = _RANDOM[12'h26C];
        v0_621 = _RANDOM[12'h26D];
        v0_622 = _RANDOM[12'h26E];
        v0_623 = _RANDOM[12'h26F];
        v0_624 = _RANDOM[12'h270];
        v0_625 = _RANDOM[12'h271];
        v0_626 = _RANDOM[12'h272];
        v0_627 = _RANDOM[12'h273];
        v0_628 = _RANDOM[12'h274];
        v0_629 = _RANDOM[12'h275];
        v0_630 = _RANDOM[12'h276];
        v0_631 = _RANDOM[12'h277];
        v0_632 = _RANDOM[12'h278];
        v0_633 = _RANDOM[12'h279];
        v0_634 = _RANDOM[12'h27A];
        v0_635 = _RANDOM[12'h27B];
        v0_636 = _RANDOM[12'h27C];
        v0_637 = _RANDOM[12'h27D];
        v0_638 = _RANDOM[12'h27E];
        v0_639 = _RANDOM[12'h27F];
        v0_640 = _RANDOM[12'h280];
        v0_641 = _RANDOM[12'h281];
        v0_642 = _RANDOM[12'h282];
        v0_643 = _RANDOM[12'h283];
        v0_644 = _RANDOM[12'h284];
        v0_645 = _RANDOM[12'h285];
        v0_646 = _RANDOM[12'h286];
        v0_647 = _RANDOM[12'h287];
        v0_648 = _RANDOM[12'h288];
        v0_649 = _RANDOM[12'h289];
        v0_650 = _RANDOM[12'h28A];
        v0_651 = _RANDOM[12'h28B];
        v0_652 = _RANDOM[12'h28C];
        v0_653 = _RANDOM[12'h28D];
        v0_654 = _RANDOM[12'h28E];
        v0_655 = _RANDOM[12'h28F];
        v0_656 = _RANDOM[12'h290];
        v0_657 = _RANDOM[12'h291];
        v0_658 = _RANDOM[12'h292];
        v0_659 = _RANDOM[12'h293];
        v0_660 = _RANDOM[12'h294];
        v0_661 = _RANDOM[12'h295];
        v0_662 = _RANDOM[12'h296];
        v0_663 = _RANDOM[12'h297];
        v0_664 = _RANDOM[12'h298];
        v0_665 = _RANDOM[12'h299];
        v0_666 = _RANDOM[12'h29A];
        v0_667 = _RANDOM[12'h29B];
        v0_668 = _RANDOM[12'h29C];
        v0_669 = _RANDOM[12'h29D];
        v0_670 = _RANDOM[12'h29E];
        v0_671 = _RANDOM[12'h29F];
        v0_672 = _RANDOM[12'h2A0];
        v0_673 = _RANDOM[12'h2A1];
        v0_674 = _RANDOM[12'h2A2];
        v0_675 = _RANDOM[12'h2A3];
        v0_676 = _RANDOM[12'h2A4];
        v0_677 = _RANDOM[12'h2A5];
        v0_678 = _RANDOM[12'h2A6];
        v0_679 = _RANDOM[12'h2A7];
        v0_680 = _RANDOM[12'h2A8];
        v0_681 = _RANDOM[12'h2A9];
        v0_682 = _RANDOM[12'h2AA];
        v0_683 = _RANDOM[12'h2AB];
        v0_684 = _RANDOM[12'h2AC];
        v0_685 = _RANDOM[12'h2AD];
        v0_686 = _RANDOM[12'h2AE];
        v0_687 = _RANDOM[12'h2AF];
        v0_688 = _RANDOM[12'h2B0];
        v0_689 = _RANDOM[12'h2B1];
        v0_690 = _RANDOM[12'h2B2];
        v0_691 = _RANDOM[12'h2B3];
        v0_692 = _RANDOM[12'h2B4];
        v0_693 = _RANDOM[12'h2B5];
        v0_694 = _RANDOM[12'h2B6];
        v0_695 = _RANDOM[12'h2B7];
        v0_696 = _RANDOM[12'h2B8];
        v0_697 = _RANDOM[12'h2B9];
        v0_698 = _RANDOM[12'h2BA];
        v0_699 = _RANDOM[12'h2BB];
        v0_700 = _RANDOM[12'h2BC];
        v0_701 = _RANDOM[12'h2BD];
        v0_702 = _RANDOM[12'h2BE];
        v0_703 = _RANDOM[12'h2BF];
        v0_704 = _RANDOM[12'h2C0];
        v0_705 = _RANDOM[12'h2C1];
        v0_706 = _RANDOM[12'h2C2];
        v0_707 = _RANDOM[12'h2C3];
        v0_708 = _RANDOM[12'h2C4];
        v0_709 = _RANDOM[12'h2C5];
        v0_710 = _RANDOM[12'h2C6];
        v0_711 = _RANDOM[12'h2C7];
        v0_712 = _RANDOM[12'h2C8];
        v0_713 = _RANDOM[12'h2C9];
        v0_714 = _RANDOM[12'h2CA];
        v0_715 = _RANDOM[12'h2CB];
        v0_716 = _RANDOM[12'h2CC];
        v0_717 = _RANDOM[12'h2CD];
        v0_718 = _RANDOM[12'h2CE];
        v0_719 = _RANDOM[12'h2CF];
        v0_720 = _RANDOM[12'h2D0];
        v0_721 = _RANDOM[12'h2D1];
        v0_722 = _RANDOM[12'h2D2];
        v0_723 = _RANDOM[12'h2D3];
        v0_724 = _RANDOM[12'h2D4];
        v0_725 = _RANDOM[12'h2D5];
        v0_726 = _RANDOM[12'h2D6];
        v0_727 = _RANDOM[12'h2D7];
        v0_728 = _RANDOM[12'h2D8];
        v0_729 = _RANDOM[12'h2D9];
        v0_730 = _RANDOM[12'h2DA];
        v0_731 = _RANDOM[12'h2DB];
        v0_732 = _RANDOM[12'h2DC];
        v0_733 = _RANDOM[12'h2DD];
        v0_734 = _RANDOM[12'h2DE];
        v0_735 = _RANDOM[12'h2DF];
        v0_736 = _RANDOM[12'h2E0];
        v0_737 = _RANDOM[12'h2E1];
        v0_738 = _RANDOM[12'h2E2];
        v0_739 = _RANDOM[12'h2E3];
        v0_740 = _RANDOM[12'h2E4];
        v0_741 = _RANDOM[12'h2E5];
        v0_742 = _RANDOM[12'h2E6];
        v0_743 = _RANDOM[12'h2E7];
        v0_744 = _RANDOM[12'h2E8];
        v0_745 = _RANDOM[12'h2E9];
        v0_746 = _RANDOM[12'h2EA];
        v0_747 = _RANDOM[12'h2EB];
        v0_748 = _RANDOM[12'h2EC];
        v0_749 = _RANDOM[12'h2ED];
        v0_750 = _RANDOM[12'h2EE];
        v0_751 = _RANDOM[12'h2EF];
        v0_752 = _RANDOM[12'h2F0];
        v0_753 = _RANDOM[12'h2F1];
        v0_754 = _RANDOM[12'h2F2];
        v0_755 = _RANDOM[12'h2F3];
        v0_756 = _RANDOM[12'h2F4];
        v0_757 = _RANDOM[12'h2F5];
        v0_758 = _RANDOM[12'h2F6];
        v0_759 = _RANDOM[12'h2F7];
        v0_760 = _RANDOM[12'h2F8];
        v0_761 = _RANDOM[12'h2F9];
        v0_762 = _RANDOM[12'h2FA];
        v0_763 = _RANDOM[12'h2FB];
        v0_764 = _RANDOM[12'h2FC];
        v0_765 = _RANDOM[12'h2FD];
        v0_766 = _RANDOM[12'h2FE];
        v0_767 = _RANDOM[12'h2FF];
        v0_768 = _RANDOM[12'h300];
        v0_769 = _RANDOM[12'h301];
        v0_770 = _RANDOM[12'h302];
        v0_771 = _RANDOM[12'h303];
        v0_772 = _RANDOM[12'h304];
        v0_773 = _RANDOM[12'h305];
        v0_774 = _RANDOM[12'h306];
        v0_775 = _RANDOM[12'h307];
        v0_776 = _RANDOM[12'h308];
        v0_777 = _RANDOM[12'h309];
        v0_778 = _RANDOM[12'h30A];
        v0_779 = _RANDOM[12'h30B];
        v0_780 = _RANDOM[12'h30C];
        v0_781 = _RANDOM[12'h30D];
        v0_782 = _RANDOM[12'h30E];
        v0_783 = _RANDOM[12'h30F];
        v0_784 = _RANDOM[12'h310];
        v0_785 = _RANDOM[12'h311];
        v0_786 = _RANDOM[12'h312];
        v0_787 = _RANDOM[12'h313];
        v0_788 = _RANDOM[12'h314];
        v0_789 = _RANDOM[12'h315];
        v0_790 = _RANDOM[12'h316];
        v0_791 = _RANDOM[12'h317];
        v0_792 = _RANDOM[12'h318];
        v0_793 = _RANDOM[12'h319];
        v0_794 = _RANDOM[12'h31A];
        v0_795 = _RANDOM[12'h31B];
        v0_796 = _RANDOM[12'h31C];
        v0_797 = _RANDOM[12'h31D];
        v0_798 = _RANDOM[12'h31E];
        v0_799 = _RANDOM[12'h31F];
        v0_800 = _RANDOM[12'h320];
        v0_801 = _RANDOM[12'h321];
        v0_802 = _RANDOM[12'h322];
        v0_803 = _RANDOM[12'h323];
        v0_804 = _RANDOM[12'h324];
        v0_805 = _RANDOM[12'h325];
        v0_806 = _RANDOM[12'h326];
        v0_807 = _RANDOM[12'h327];
        v0_808 = _RANDOM[12'h328];
        v0_809 = _RANDOM[12'h329];
        v0_810 = _RANDOM[12'h32A];
        v0_811 = _RANDOM[12'h32B];
        v0_812 = _RANDOM[12'h32C];
        v0_813 = _RANDOM[12'h32D];
        v0_814 = _RANDOM[12'h32E];
        v0_815 = _RANDOM[12'h32F];
        v0_816 = _RANDOM[12'h330];
        v0_817 = _RANDOM[12'h331];
        v0_818 = _RANDOM[12'h332];
        v0_819 = _RANDOM[12'h333];
        v0_820 = _RANDOM[12'h334];
        v0_821 = _RANDOM[12'h335];
        v0_822 = _RANDOM[12'h336];
        v0_823 = _RANDOM[12'h337];
        v0_824 = _RANDOM[12'h338];
        v0_825 = _RANDOM[12'h339];
        v0_826 = _RANDOM[12'h33A];
        v0_827 = _RANDOM[12'h33B];
        v0_828 = _RANDOM[12'h33C];
        v0_829 = _RANDOM[12'h33D];
        v0_830 = _RANDOM[12'h33E];
        v0_831 = _RANDOM[12'h33F];
        v0_832 = _RANDOM[12'h340];
        v0_833 = _RANDOM[12'h341];
        v0_834 = _RANDOM[12'h342];
        v0_835 = _RANDOM[12'h343];
        v0_836 = _RANDOM[12'h344];
        v0_837 = _RANDOM[12'h345];
        v0_838 = _RANDOM[12'h346];
        v0_839 = _RANDOM[12'h347];
        v0_840 = _RANDOM[12'h348];
        v0_841 = _RANDOM[12'h349];
        v0_842 = _RANDOM[12'h34A];
        v0_843 = _RANDOM[12'h34B];
        v0_844 = _RANDOM[12'h34C];
        v0_845 = _RANDOM[12'h34D];
        v0_846 = _RANDOM[12'h34E];
        v0_847 = _RANDOM[12'h34F];
        v0_848 = _RANDOM[12'h350];
        v0_849 = _RANDOM[12'h351];
        v0_850 = _RANDOM[12'h352];
        v0_851 = _RANDOM[12'h353];
        v0_852 = _RANDOM[12'h354];
        v0_853 = _RANDOM[12'h355];
        v0_854 = _RANDOM[12'h356];
        v0_855 = _RANDOM[12'h357];
        v0_856 = _RANDOM[12'h358];
        v0_857 = _RANDOM[12'h359];
        v0_858 = _RANDOM[12'h35A];
        v0_859 = _RANDOM[12'h35B];
        v0_860 = _RANDOM[12'h35C];
        v0_861 = _RANDOM[12'h35D];
        v0_862 = _RANDOM[12'h35E];
        v0_863 = _RANDOM[12'h35F];
        v0_864 = _RANDOM[12'h360];
        v0_865 = _RANDOM[12'h361];
        v0_866 = _RANDOM[12'h362];
        v0_867 = _RANDOM[12'h363];
        v0_868 = _RANDOM[12'h364];
        v0_869 = _RANDOM[12'h365];
        v0_870 = _RANDOM[12'h366];
        v0_871 = _RANDOM[12'h367];
        v0_872 = _RANDOM[12'h368];
        v0_873 = _RANDOM[12'h369];
        v0_874 = _RANDOM[12'h36A];
        v0_875 = _RANDOM[12'h36B];
        v0_876 = _RANDOM[12'h36C];
        v0_877 = _RANDOM[12'h36D];
        v0_878 = _RANDOM[12'h36E];
        v0_879 = _RANDOM[12'h36F];
        v0_880 = _RANDOM[12'h370];
        v0_881 = _RANDOM[12'h371];
        v0_882 = _RANDOM[12'h372];
        v0_883 = _RANDOM[12'h373];
        v0_884 = _RANDOM[12'h374];
        v0_885 = _RANDOM[12'h375];
        v0_886 = _RANDOM[12'h376];
        v0_887 = _RANDOM[12'h377];
        v0_888 = _RANDOM[12'h378];
        v0_889 = _RANDOM[12'h379];
        v0_890 = _RANDOM[12'h37A];
        v0_891 = _RANDOM[12'h37B];
        v0_892 = _RANDOM[12'h37C];
        v0_893 = _RANDOM[12'h37D];
        v0_894 = _RANDOM[12'h37E];
        v0_895 = _RANDOM[12'h37F];
        v0_896 = _RANDOM[12'h380];
        v0_897 = _RANDOM[12'h381];
        v0_898 = _RANDOM[12'h382];
        v0_899 = _RANDOM[12'h383];
        v0_900 = _RANDOM[12'h384];
        v0_901 = _RANDOM[12'h385];
        v0_902 = _RANDOM[12'h386];
        v0_903 = _RANDOM[12'h387];
        v0_904 = _RANDOM[12'h388];
        v0_905 = _RANDOM[12'h389];
        v0_906 = _RANDOM[12'h38A];
        v0_907 = _RANDOM[12'h38B];
        v0_908 = _RANDOM[12'h38C];
        v0_909 = _RANDOM[12'h38D];
        v0_910 = _RANDOM[12'h38E];
        v0_911 = _RANDOM[12'h38F];
        v0_912 = _RANDOM[12'h390];
        v0_913 = _RANDOM[12'h391];
        v0_914 = _RANDOM[12'h392];
        v0_915 = _RANDOM[12'h393];
        v0_916 = _RANDOM[12'h394];
        v0_917 = _RANDOM[12'h395];
        v0_918 = _RANDOM[12'h396];
        v0_919 = _RANDOM[12'h397];
        v0_920 = _RANDOM[12'h398];
        v0_921 = _RANDOM[12'h399];
        v0_922 = _RANDOM[12'h39A];
        v0_923 = _RANDOM[12'h39B];
        v0_924 = _RANDOM[12'h39C];
        v0_925 = _RANDOM[12'h39D];
        v0_926 = _RANDOM[12'h39E];
        v0_927 = _RANDOM[12'h39F];
        v0_928 = _RANDOM[12'h3A0];
        v0_929 = _RANDOM[12'h3A1];
        v0_930 = _RANDOM[12'h3A2];
        v0_931 = _RANDOM[12'h3A3];
        v0_932 = _RANDOM[12'h3A4];
        v0_933 = _RANDOM[12'h3A5];
        v0_934 = _RANDOM[12'h3A6];
        v0_935 = _RANDOM[12'h3A7];
        v0_936 = _RANDOM[12'h3A8];
        v0_937 = _RANDOM[12'h3A9];
        v0_938 = _RANDOM[12'h3AA];
        v0_939 = _RANDOM[12'h3AB];
        v0_940 = _RANDOM[12'h3AC];
        v0_941 = _RANDOM[12'h3AD];
        v0_942 = _RANDOM[12'h3AE];
        v0_943 = _RANDOM[12'h3AF];
        v0_944 = _RANDOM[12'h3B0];
        v0_945 = _RANDOM[12'h3B1];
        v0_946 = _RANDOM[12'h3B2];
        v0_947 = _RANDOM[12'h3B3];
        v0_948 = _RANDOM[12'h3B4];
        v0_949 = _RANDOM[12'h3B5];
        v0_950 = _RANDOM[12'h3B6];
        v0_951 = _RANDOM[12'h3B7];
        v0_952 = _RANDOM[12'h3B8];
        v0_953 = _RANDOM[12'h3B9];
        v0_954 = _RANDOM[12'h3BA];
        v0_955 = _RANDOM[12'h3BB];
        v0_956 = _RANDOM[12'h3BC];
        v0_957 = _RANDOM[12'h3BD];
        v0_958 = _RANDOM[12'h3BE];
        v0_959 = _RANDOM[12'h3BF];
        v0_960 = _RANDOM[12'h3C0];
        v0_961 = _RANDOM[12'h3C1];
        v0_962 = _RANDOM[12'h3C2];
        v0_963 = _RANDOM[12'h3C3];
        v0_964 = _RANDOM[12'h3C4];
        v0_965 = _RANDOM[12'h3C5];
        v0_966 = _RANDOM[12'h3C6];
        v0_967 = _RANDOM[12'h3C7];
        v0_968 = _RANDOM[12'h3C8];
        v0_969 = _RANDOM[12'h3C9];
        v0_970 = _RANDOM[12'h3CA];
        v0_971 = _RANDOM[12'h3CB];
        v0_972 = _RANDOM[12'h3CC];
        v0_973 = _RANDOM[12'h3CD];
        v0_974 = _RANDOM[12'h3CE];
        v0_975 = _RANDOM[12'h3CF];
        v0_976 = _RANDOM[12'h3D0];
        v0_977 = _RANDOM[12'h3D1];
        v0_978 = _RANDOM[12'h3D2];
        v0_979 = _RANDOM[12'h3D3];
        v0_980 = _RANDOM[12'h3D4];
        v0_981 = _RANDOM[12'h3D5];
        v0_982 = _RANDOM[12'h3D6];
        v0_983 = _RANDOM[12'h3D7];
        v0_984 = _RANDOM[12'h3D8];
        v0_985 = _RANDOM[12'h3D9];
        v0_986 = _RANDOM[12'h3DA];
        v0_987 = _RANDOM[12'h3DB];
        v0_988 = _RANDOM[12'h3DC];
        v0_989 = _RANDOM[12'h3DD];
        v0_990 = _RANDOM[12'h3DE];
        v0_991 = _RANDOM[12'h3DF];
        v0_992 = _RANDOM[12'h3E0];
        v0_993 = _RANDOM[12'h3E1];
        v0_994 = _RANDOM[12'h3E2];
        v0_995 = _RANDOM[12'h3E3];
        v0_996 = _RANDOM[12'h3E4];
        v0_997 = _RANDOM[12'h3E5];
        v0_998 = _RANDOM[12'h3E6];
        v0_999 = _RANDOM[12'h3E7];
        v0_1000 = _RANDOM[12'h3E8];
        v0_1001 = _RANDOM[12'h3E9];
        v0_1002 = _RANDOM[12'h3EA];
        v0_1003 = _RANDOM[12'h3EB];
        v0_1004 = _RANDOM[12'h3EC];
        v0_1005 = _RANDOM[12'h3ED];
        v0_1006 = _RANDOM[12'h3EE];
        v0_1007 = _RANDOM[12'h3EF];
        v0_1008 = _RANDOM[12'h3F0];
        v0_1009 = _RANDOM[12'h3F1];
        v0_1010 = _RANDOM[12'h3F2];
        v0_1011 = _RANDOM[12'h3F3];
        v0_1012 = _RANDOM[12'h3F4];
        v0_1013 = _RANDOM[12'h3F5];
        v0_1014 = _RANDOM[12'h3F6];
        v0_1015 = _RANDOM[12'h3F7];
        v0_1016 = _RANDOM[12'h3F8];
        v0_1017 = _RANDOM[12'h3F9];
        v0_1018 = _RANDOM[12'h3FA];
        v0_1019 = _RANDOM[12'h3FB];
        v0_1020 = _RANDOM[12'h3FC];
        v0_1021 = _RANDOM[12'h3FD];
        v0_1022 = _RANDOM[12'h3FE];
        v0_1023 = _RANDOM[12'h3FF];
        v0_1024 = _RANDOM[12'h400];
        v0_1025 = _RANDOM[12'h401];
        v0_1026 = _RANDOM[12'h402];
        v0_1027 = _RANDOM[12'h403];
        v0_1028 = _RANDOM[12'h404];
        v0_1029 = _RANDOM[12'h405];
        v0_1030 = _RANDOM[12'h406];
        v0_1031 = _RANDOM[12'h407];
        v0_1032 = _RANDOM[12'h408];
        v0_1033 = _RANDOM[12'h409];
        v0_1034 = _RANDOM[12'h40A];
        v0_1035 = _RANDOM[12'h40B];
        v0_1036 = _RANDOM[12'h40C];
        v0_1037 = _RANDOM[12'h40D];
        v0_1038 = _RANDOM[12'h40E];
        v0_1039 = _RANDOM[12'h40F];
        v0_1040 = _RANDOM[12'h410];
        v0_1041 = _RANDOM[12'h411];
        v0_1042 = _RANDOM[12'h412];
        v0_1043 = _RANDOM[12'h413];
        v0_1044 = _RANDOM[12'h414];
        v0_1045 = _RANDOM[12'h415];
        v0_1046 = _RANDOM[12'h416];
        v0_1047 = _RANDOM[12'h417];
        v0_1048 = _RANDOM[12'h418];
        v0_1049 = _RANDOM[12'h419];
        v0_1050 = _RANDOM[12'h41A];
        v0_1051 = _RANDOM[12'h41B];
        v0_1052 = _RANDOM[12'h41C];
        v0_1053 = _RANDOM[12'h41D];
        v0_1054 = _RANDOM[12'h41E];
        v0_1055 = _RANDOM[12'h41F];
        v0_1056 = _RANDOM[12'h420];
        v0_1057 = _RANDOM[12'h421];
        v0_1058 = _RANDOM[12'h422];
        v0_1059 = _RANDOM[12'h423];
        v0_1060 = _RANDOM[12'h424];
        v0_1061 = _RANDOM[12'h425];
        v0_1062 = _RANDOM[12'h426];
        v0_1063 = _RANDOM[12'h427];
        v0_1064 = _RANDOM[12'h428];
        v0_1065 = _RANDOM[12'h429];
        v0_1066 = _RANDOM[12'h42A];
        v0_1067 = _RANDOM[12'h42B];
        v0_1068 = _RANDOM[12'h42C];
        v0_1069 = _RANDOM[12'h42D];
        v0_1070 = _RANDOM[12'h42E];
        v0_1071 = _RANDOM[12'h42F];
        v0_1072 = _RANDOM[12'h430];
        v0_1073 = _RANDOM[12'h431];
        v0_1074 = _RANDOM[12'h432];
        v0_1075 = _RANDOM[12'h433];
        v0_1076 = _RANDOM[12'h434];
        v0_1077 = _RANDOM[12'h435];
        v0_1078 = _RANDOM[12'h436];
        v0_1079 = _RANDOM[12'h437];
        v0_1080 = _RANDOM[12'h438];
        v0_1081 = _RANDOM[12'h439];
        v0_1082 = _RANDOM[12'h43A];
        v0_1083 = _RANDOM[12'h43B];
        v0_1084 = _RANDOM[12'h43C];
        v0_1085 = _RANDOM[12'h43D];
        v0_1086 = _RANDOM[12'h43E];
        v0_1087 = _RANDOM[12'h43F];
        v0_1088 = _RANDOM[12'h440];
        v0_1089 = _RANDOM[12'h441];
        v0_1090 = _RANDOM[12'h442];
        v0_1091 = _RANDOM[12'h443];
        v0_1092 = _RANDOM[12'h444];
        v0_1093 = _RANDOM[12'h445];
        v0_1094 = _RANDOM[12'h446];
        v0_1095 = _RANDOM[12'h447];
        v0_1096 = _RANDOM[12'h448];
        v0_1097 = _RANDOM[12'h449];
        v0_1098 = _RANDOM[12'h44A];
        v0_1099 = _RANDOM[12'h44B];
        v0_1100 = _RANDOM[12'h44C];
        v0_1101 = _RANDOM[12'h44D];
        v0_1102 = _RANDOM[12'h44E];
        v0_1103 = _RANDOM[12'h44F];
        v0_1104 = _RANDOM[12'h450];
        v0_1105 = _RANDOM[12'h451];
        v0_1106 = _RANDOM[12'h452];
        v0_1107 = _RANDOM[12'h453];
        v0_1108 = _RANDOM[12'h454];
        v0_1109 = _RANDOM[12'h455];
        v0_1110 = _RANDOM[12'h456];
        v0_1111 = _RANDOM[12'h457];
        v0_1112 = _RANDOM[12'h458];
        v0_1113 = _RANDOM[12'h459];
        v0_1114 = _RANDOM[12'h45A];
        v0_1115 = _RANDOM[12'h45B];
        v0_1116 = _RANDOM[12'h45C];
        v0_1117 = _RANDOM[12'h45D];
        v0_1118 = _RANDOM[12'h45E];
        v0_1119 = _RANDOM[12'h45F];
        v0_1120 = _RANDOM[12'h460];
        v0_1121 = _RANDOM[12'h461];
        v0_1122 = _RANDOM[12'h462];
        v0_1123 = _RANDOM[12'h463];
        v0_1124 = _RANDOM[12'h464];
        v0_1125 = _RANDOM[12'h465];
        v0_1126 = _RANDOM[12'h466];
        v0_1127 = _RANDOM[12'h467];
        v0_1128 = _RANDOM[12'h468];
        v0_1129 = _RANDOM[12'h469];
        v0_1130 = _RANDOM[12'h46A];
        v0_1131 = _RANDOM[12'h46B];
        v0_1132 = _RANDOM[12'h46C];
        v0_1133 = _RANDOM[12'h46D];
        v0_1134 = _RANDOM[12'h46E];
        v0_1135 = _RANDOM[12'h46F];
        v0_1136 = _RANDOM[12'h470];
        v0_1137 = _RANDOM[12'h471];
        v0_1138 = _RANDOM[12'h472];
        v0_1139 = _RANDOM[12'h473];
        v0_1140 = _RANDOM[12'h474];
        v0_1141 = _RANDOM[12'h475];
        v0_1142 = _RANDOM[12'h476];
        v0_1143 = _RANDOM[12'h477];
        v0_1144 = _RANDOM[12'h478];
        v0_1145 = _RANDOM[12'h479];
        v0_1146 = _RANDOM[12'h47A];
        v0_1147 = _RANDOM[12'h47B];
        v0_1148 = _RANDOM[12'h47C];
        v0_1149 = _RANDOM[12'h47D];
        v0_1150 = _RANDOM[12'h47E];
        v0_1151 = _RANDOM[12'h47F];
        v0_1152 = _RANDOM[12'h480];
        v0_1153 = _RANDOM[12'h481];
        v0_1154 = _RANDOM[12'h482];
        v0_1155 = _RANDOM[12'h483];
        v0_1156 = _RANDOM[12'h484];
        v0_1157 = _RANDOM[12'h485];
        v0_1158 = _RANDOM[12'h486];
        v0_1159 = _RANDOM[12'h487];
        v0_1160 = _RANDOM[12'h488];
        v0_1161 = _RANDOM[12'h489];
        v0_1162 = _RANDOM[12'h48A];
        v0_1163 = _RANDOM[12'h48B];
        v0_1164 = _RANDOM[12'h48C];
        v0_1165 = _RANDOM[12'h48D];
        v0_1166 = _RANDOM[12'h48E];
        v0_1167 = _RANDOM[12'h48F];
        v0_1168 = _RANDOM[12'h490];
        v0_1169 = _RANDOM[12'h491];
        v0_1170 = _RANDOM[12'h492];
        v0_1171 = _RANDOM[12'h493];
        v0_1172 = _RANDOM[12'h494];
        v0_1173 = _RANDOM[12'h495];
        v0_1174 = _RANDOM[12'h496];
        v0_1175 = _RANDOM[12'h497];
        v0_1176 = _RANDOM[12'h498];
        v0_1177 = _RANDOM[12'h499];
        v0_1178 = _RANDOM[12'h49A];
        v0_1179 = _RANDOM[12'h49B];
        v0_1180 = _RANDOM[12'h49C];
        v0_1181 = _RANDOM[12'h49D];
        v0_1182 = _RANDOM[12'h49E];
        v0_1183 = _RANDOM[12'h49F];
        v0_1184 = _RANDOM[12'h4A0];
        v0_1185 = _RANDOM[12'h4A1];
        v0_1186 = _RANDOM[12'h4A2];
        v0_1187 = _RANDOM[12'h4A3];
        v0_1188 = _RANDOM[12'h4A4];
        v0_1189 = _RANDOM[12'h4A5];
        v0_1190 = _RANDOM[12'h4A6];
        v0_1191 = _RANDOM[12'h4A7];
        v0_1192 = _RANDOM[12'h4A8];
        v0_1193 = _RANDOM[12'h4A9];
        v0_1194 = _RANDOM[12'h4AA];
        v0_1195 = _RANDOM[12'h4AB];
        v0_1196 = _RANDOM[12'h4AC];
        v0_1197 = _RANDOM[12'h4AD];
        v0_1198 = _RANDOM[12'h4AE];
        v0_1199 = _RANDOM[12'h4AF];
        v0_1200 = _RANDOM[12'h4B0];
        v0_1201 = _RANDOM[12'h4B1];
        v0_1202 = _RANDOM[12'h4B2];
        v0_1203 = _RANDOM[12'h4B3];
        v0_1204 = _RANDOM[12'h4B4];
        v0_1205 = _RANDOM[12'h4B5];
        v0_1206 = _RANDOM[12'h4B6];
        v0_1207 = _RANDOM[12'h4B7];
        v0_1208 = _RANDOM[12'h4B8];
        v0_1209 = _RANDOM[12'h4B9];
        v0_1210 = _RANDOM[12'h4BA];
        v0_1211 = _RANDOM[12'h4BB];
        v0_1212 = _RANDOM[12'h4BC];
        v0_1213 = _RANDOM[12'h4BD];
        v0_1214 = _RANDOM[12'h4BE];
        v0_1215 = _RANDOM[12'h4BF];
        v0_1216 = _RANDOM[12'h4C0];
        v0_1217 = _RANDOM[12'h4C1];
        v0_1218 = _RANDOM[12'h4C2];
        v0_1219 = _RANDOM[12'h4C3];
        v0_1220 = _RANDOM[12'h4C4];
        v0_1221 = _RANDOM[12'h4C5];
        v0_1222 = _RANDOM[12'h4C6];
        v0_1223 = _RANDOM[12'h4C7];
        v0_1224 = _RANDOM[12'h4C8];
        v0_1225 = _RANDOM[12'h4C9];
        v0_1226 = _RANDOM[12'h4CA];
        v0_1227 = _RANDOM[12'h4CB];
        v0_1228 = _RANDOM[12'h4CC];
        v0_1229 = _RANDOM[12'h4CD];
        v0_1230 = _RANDOM[12'h4CE];
        v0_1231 = _RANDOM[12'h4CF];
        v0_1232 = _RANDOM[12'h4D0];
        v0_1233 = _RANDOM[12'h4D1];
        v0_1234 = _RANDOM[12'h4D2];
        v0_1235 = _RANDOM[12'h4D3];
        v0_1236 = _RANDOM[12'h4D4];
        v0_1237 = _RANDOM[12'h4D5];
        v0_1238 = _RANDOM[12'h4D6];
        v0_1239 = _RANDOM[12'h4D7];
        v0_1240 = _RANDOM[12'h4D8];
        v0_1241 = _RANDOM[12'h4D9];
        v0_1242 = _RANDOM[12'h4DA];
        v0_1243 = _RANDOM[12'h4DB];
        v0_1244 = _RANDOM[12'h4DC];
        v0_1245 = _RANDOM[12'h4DD];
        v0_1246 = _RANDOM[12'h4DE];
        v0_1247 = _RANDOM[12'h4DF];
        v0_1248 = _RANDOM[12'h4E0];
        v0_1249 = _RANDOM[12'h4E1];
        v0_1250 = _RANDOM[12'h4E2];
        v0_1251 = _RANDOM[12'h4E3];
        v0_1252 = _RANDOM[12'h4E4];
        v0_1253 = _RANDOM[12'h4E5];
        v0_1254 = _RANDOM[12'h4E6];
        v0_1255 = _RANDOM[12'h4E7];
        v0_1256 = _RANDOM[12'h4E8];
        v0_1257 = _RANDOM[12'h4E9];
        v0_1258 = _RANDOM[12'h4EA];
        v0_1259 = _RANDOM[12'h4EB];
        v0_1260 = _RANDOM[12'h4EC];
        v0_1261 = _RANDOM[12'h4ED];
        v0_1262 = _RANDOM[12'h4EE];
        v0_1263 = _RANDOM[12'h4EF];
        v0_1264 = _RANDOM[12'h4F0];
        v0_1265 = _RANDOM[12'h4F1];
        v0_1266 = _RANDOM[12'h4F2];
        v0_1267 = _RANDOM[12'h4F3];
        v0_1268 = _RANDOM[12'h4F4];
        v0_1269 = _RANDOM[12'h4F5];
        v0_1270 = _RANDOM[12'h4F6];
        v0_1271 = _RANDOM[12'h4F7];
        v0_1272 = _RANDOM[12'h4F8];
        v0_1273 = _RANDOM[12'h4F9];
        v0_1274 = _RANDOM[12'h4FA];
        v0_1275 = _RANDOM[12'h4FB];
        v0_1276 = _RANDOM[12'h4FC];
        v0_1277 = _RANDOM[12'h4FD];
        v0_1278 = _RANDOM[12'h4FE];
        v0_1279 = _RANDOM[12'h4FF];
        v0_1280 = _RANDOM[12'h500];
        v0_1281 = _RANDOM[12'h501];
        v0_1282 = _RANDOM[12'h502];
        v0_1283 = _RANDOM[12'h503];
        v0_1284 = _RANDOM[12'h504];
        v0_1285 = _RANDOM[12'h505];
        v0_1286 = _RANDOM[12'h506];
        v0_1287 = _RANDOM[12'h507];
        v0_1288 = _RANDOM[12'h508];
        v0_1289 = _RANDOM[12'h509];
        v0_1290 = _RANDOM[12'h50A];
        v0_1291 = _RANDOM[12'h50B];
        v0_1292 = _RANDOM[12'h50C];
        v0_1293 = _RANDOM[12'h50D];
        v0_1294 = _RANDOM[12'h50E];
        v0_1295 = _RANDOM[12'h50F];
        v0_1296 = _RANDOM[12'h510];
        v0_1297 = _RANDOM[12'h511];
        v0_1298 = _RANDOM[12'h512];
        v0_1299 = _RANDOM[12'h513];
        v0_1300 = _RANDOM[12'h514];
        v0_1301 = _RANDOM[12'h515];
        v0_1302 = _RANDOM[12'h516];
        v0_1303 = _RANDOM[12'h517];
        v0_1304 = _RANDOM[12'h518];
        v0_1305 = _RANDOM[12'h519];
        v0_1306 = _RANDOM[12'h51A];
        v0_1307 = _RANDOM[12'h51B];
        v0_1308 = _RANDOM[12'h51C];
        v0_1309 = _RANDOM[12'h51D];
        v0_1310 = _RANDOM[12'h51E];
        v0_1311 = _RANDOM[12'h51F];
        v0_1312 = _RANDOM[12'h520];
        v0_1313 = _RANDOM[12'h521];
        v0_1314 = _RANDOM[12'h522];
        v0_1315 = _RANDOM[12'h523];
        v0_1316 = _RANDOM[12'h524];
        v0_1317 = _RANDOM[12'h525];
        v0_1318 = _RANDOM[12'h526];
        v0_1319 = _RANDOM[12'h527];
        v0_1320 = _RANDOM[12'h528];
        v0_1321 = _RANDOM[12'h529];
        v0_1322 = _RANDOM[12'h52A];
        v0_1323 = _RANDOM[12'h52B];
        v0_1324 = _RANDOM[12'h52C];
        v0_1325 = _RANDOM[12'h52D];
        v0_1326 = _RANDOM[12'h52E];
        v0_1327 = _RANDOM[12'h52F];
        v0_1328 = _RANDOM[12'h530];
        v0_1329 = _RANDOM[12'h531];
        v0_1330 = _RANDOM[12'h532];
        v0_1331 = _RANDOM[12'h533];
        v0_1332 = _RANDOM[12'h534];
        v0_1333 = _RANDOM[12'h535];
        v0_1334 = _RANDOM[12'h536];
        v0_1335 = _RANDOM[12'h537];
        v0_1336 = _RANDOM[12'h538];
        v0_1337 = _RANDOM[12'h539];
        v0_1338 = _RANDOM[12'h53A];
        v0_1339 = _RANDOM[12'h53B];
        v0_1340 = _RANDOM[12'h53C];
        v0_1341 = _RANDOM[12'h53D];
        v0_1342 = _RANDOM[12'h53E];
        v0_1343 = _RANDOM[12'h53F];
        v0_1344 = _RANDOM[12'h540];
        v0_1345 = _RANDOM[12'h541];
        v0_1346 = _RANDOM[12'h542];
        v0_1347 = _RANDOM[12'h543];
        v0_1348 = _RANDOM[12'h544];
        v0_1349 = _RANDOM[12'h545];
        v0_1350 = _RANDOM[12'h546];
        v0_1351 = _RANDOM[12'h547];
        v0_1352 = _RANDOM[12'h548];
        v0_1353 = _RANDOM[12'h549];
        v0_1354 = _RANDOM[12'h54A];
        v0_1355 = _RANDOM[12'h54B];
        v0_1356 = _RANDOM[12'h54C];
        v0_1357 = _RANDOM[12'h54D];
        v0_1358 = _RANDOM[12'h54E];
        v0_1359 = _RANDOM[12'h54F];
        v0_1360 = _RANDOM[12'h550];
        v0_1361 = _RANDOM[12'h551];
        v0_1362 = _RANDOM[12'h552];
        v0_1363 = _RANDOM[12'h553];
        v0_1364 = _RANDOM[12'h554];
        v0_1365 = _RANDOM[12'h555];
        v0_1366 = _RANDOM[12'h556];
        v0_1367 = _RANDOM[12'h557];
        v0_1368 = _RANDOM[12'h558];
        v0_1369 = _RANDOM[12'h559];
        v0_1370 = _RANDOM[12'h55A];
        v0_1371 = _RANDOM[12'h55B];
        v0_1372 = _RANDOM[12'h55C];
        v0_1373 = _RANDOM[12'h55D];
        v0_1374 = _RANDOM[12'h55E];
        v0_1375 = _RANDOM[12'h55F];
        v0_1376 = _RANDOM[12'h560];
        v0_1377 = _RANDOM[12'h561];
        v0_1378 = _RANDOM[12'h562];
        v0_1379 = _RANDOM[12'h563];
        v0_1380 = _RANDOM[12'h564];
        v0_1381 = _RANDOM[12'h565];
        v0_1382 = _RANDOM[12'h566];
        v0_1383 = _RANDOM[12'h567];
        v0_1384 = _RANDOM[12'h568];
        v0_1385 = _RANDOM[12'h569];
        v0_1386 = _RANDOM[12'h56A];
        v0_1387 = _RANDOM[12'h56B];
        v0_1388 = _RANDOM[12'h56C];
        v0_1389 = _RANDOM[12'h56D];
        v0_1390 = _RANDOM[12'h56E];
        v0_1391 = _RANDOM[12'h56F];
        v0_1392 = _RANDOM[12'h570];
        v0_1393 = _RANDOM[12'h571];
        v0_1394 = _RANDOM[12'h572];
        v0_1395 = _RANDOM[12'h573];
        v0_1396 = _RANDOM[12'h574];
        v0_1397 = _RANDOM[12'h575];
        v0_1398 = _RANDOM[12'h576];
        v0_1399 = _RANDOM[12'h577];
        v0_1400 = _RANDOM[12'h578];
        v0_1401 = _RANDOM[12'h579];
        v0_1402 = _RANDOM[12'h57A];
        v0_1403 = _RANDOM[12'h57B];
        v0_1404 = _RANDOM[12'h57C];
        v0_1405 = _RANDOM[12'h57D];
        v0_1406 = _RANDOM[12'h57E];
        v0_1407 = _RANDOM[12'h57F];
        v0_1408 = _RANDOM[12'h580];
        v0_1409 = _RANDOM[12'h581];
        v0_1410 = _RANDOM[12'h582];
        v0_1411 = _RANDOM[12'h583];
        v0_1412 = _RANDOM[12'h584];
        v0_1413 = _RANDOM[12'h585];
        v0_1414 = _RANDOM[12'h586];
        v0_1415 = _RANDOM[12'h587];
        v0_1416 = _RANDOM[12'h588];
        v0_1417 = _RANDOM[12'h589];
        v0_1418 = _RANDOM[12'h58A];
        v0_1419 = _RANDOM[12'h58B];
        v0_1420 = _RANDOM[12'h58C];
        v0_1421 = _RANDOM[12'h58D];
        v0_1422 = _RANDOM[12'h58E];
        v0_1423 = _RANDOM[12'h58F];
        v0_1424 = _RANDOM[12'h590];
        v0_1425 = _RANDOM[12'h591];
        v0_1426 = _RANDOM[12'h592];
        v0_1427 = _RANDOM[12'h593];
        v0_1428 = _RANDOM[12'h594];
        v0_1429 = _RANDOM[12'h595];
        v0_1430 = _RANDOM[12'h596];
        v0_1431 = _RANDOM[12'h597];
        v0_1432 = _RANDOM[12'h598];
        v0_1433 = _RANDOM[12'h599];
        v0_1434 = _RANDOM[12'h59A];
        v0_1435 = _RANDOM[12'h59B];
        v0_1436 = _RANDOM[12'h59C];
        v0_1437 = _RANDOM[12'h59D];
        v0_1438 = _RANDOM[12'h59E];
        v0_1439 = _RANDOM[12'h59F];
        v0_1440 = _RANDOM[12'h5A0];
        v0_1441 = _RANDOM[12'h5A1];
        v0_1442 = _RANDOM[12'h5A2];
        v0_1443 = _RANDOM[12'h5A3];
        v0_1444 = _RANDOM[12'h5A4];
        v0_1445 = _RANDOM[12'h5A5];
        v0_1446 = _RANDOM[12'h5A6];
        v0_1447 = _RANDOM[12'h5A7];
        v0_1448 = _RANDOM[12'h5A8];
        v0_1449 = _RANDOM[12'h5A9];
        v0_1450 = _RANDOM[12'h5AA];
        v0_1451 = _RANDOM[12'h5AB];
        v0_1452 = _RANDOM[12'h5AC];
        v0_1453 = _RANDOM[12'h5AD];
        v0_1454 = _RANDOM[12'h5AE];
        v0_1455 = _RANDOM[12'h5AF];
        v0_1456 = _RANDOM[12'h5B0];
        v0_1457 = _RANDOM[12'h5B1];
        v0_1458 = _RANDOM[12'h5B2];
        v0_1459 = _RANDOM[12'h5B3];
        v0_1460 = _RANDOM[12'h5B4];
        v0_1461 = _RANDOM[12'h5B5];
        v0_1462 = _RANDOM[12'h5B6];
        v0_1463 = _RANDOM[12'h5B7];
        v0_1464 = _RANDOM[12'h5B8];
        v0_1465 = _RANDOM[12'h5B9];
        v0_1466 = _RANDOM[12'h5BA];
        v0_1467 = _RANDOM[12'h5BB];
        v0_1468 = _RANDOM[12'h5BC];
        v0_1469 = _RANDOM[12'h5BD];
        v0_1470 = _RANDOM[12'h5BE];
        v0_1471 = _RANDOM[12'h5BF];
        v0_1472 = _RANDOM[12'h5C0];
        v0_1473 = _RANDOM[12'h5C1];
        v0_1474 = _RANDOM[12'h5C2];
        v0_1475 = _RANDOM[12'h5C3];
        v0_1476 = _RANDOM[12'h5C4];
        v0_1477 = _RANDOM[12'h5C5];
        v0_1478 = _RANDOM[12'h5C6];
        v0_1479 = _RANDOM[12'h5C7];
        v0_1480 = _RANDOM[12'h5C8];
        v0_1481 = _RANDOM[12'h5C9];
        v0_1482 = _RANDOM[12'h5CA];
        v0_1483 = _RANDOM[12'h5CB];
        v0_1484 = _RANDOM[12'h5CC];
        v0_1485 = _RANDOM[12'h5CD];
        v0_1486 = _RANDOM[12'h5CE];
        v0_1487 = _RANDOM[12'h5CF];
        v0_1488 = _RANDOM[12'h5D0];
        v0_1489 = _RANDOM[12'h5D1];
        v0_1490 = _RANDOM[12'h5D2];
        v0_1491 = _RANDOM[12'h5D3];
        v0_1492 = _RANDOM[12'h5D4];
        v0_1493 = _RANDOM[12'h5D5];
        v0_1494 = _RANDOM[12'h5D6];
        v0_1495 = _RANDOM[12'h5D7];
        v0_1496 = _RANDOM[12'h5D8];
        v0_1497 = _RANDOM[12'h5D9];
        v0_1498 = _RANDOM[12'h5DA];
        v0_1499 = _RANDOM[12'h5DB];
        v0_1500 = _RANDOM[12'h5DC];
        v0_1501 = _RANDOM[12'h5DD];
        v0_1502 = _RANDOM[12'h5DE];
        v0_1503 = _RANDOM[12'h5DF];
        v0_1504 = _RANDOM[12'h5E0];
        v0_1505 = _RANDOM[12'h5E1];
        v0_1506 = _RANDOM[12'h5E2];
        v0_1507 = _RANDOM[12'h5E3];
        v0_1508 = _RANDOM[12'h5E4];
        v0_1509 = _RANDOM[12'h5E5];
        v0_1510 = _RANDOM[12'h5E6];
        v0_1511 = _RANDOM[12'h5E7];
        v0_1512 = _RANDOM[12'h5E8];
        v0_1513 = _RANDOM[12'h5E9];
        v0_1514 = _RANDOM[12'h5EA];
        v0_1515 = _RANDOM[12'h5EB];
        v0_1516 = _RANDOM[12'h5EC];
        v0_1517 = _RANDOM[12'h5ED];
        v0_1518 = _RANDOM[12'h5EE];
        v0_1519 = _RANDOM[12'h5EF];
        v0_1520 = _RANDOM[12'h5F0];
        v0_1521 = _RANDOM[12'h5F1];
        v0_1522 = _RANDOM[12'h5F2];
        v0_1523 = _RANDOM[12'h5F3];
        v0_1524 = _RANDOM[12'h5F4];
        v0_1525 = _RANDOM[12'h5F5];
        v0_1526 = _RANDOM[12'h5F6];
        v0_1527 = _RANDOM[12'h5F7];
        v0_1528 = _RANDOM[12'h5F8];
        v0_1529 = _RANDOM[12'h5F9];
        v0_1530 = _RANDOM[12'h5FA];
        v0_1531 = _RANDOM[12'h5FB];
        v0_1532 = _RANDOM[12'h5FC];
        v0_1533 = _RANDOM[12'h5FD];
        v0_1534 = _RANDOM[12'h5FE];
        v0_1535 = _RANDOM[12'h5FF];
        v0_1536 = _RANDOM[12'h600];
        v0_1537 = _RANDOM[12'h601];
        v0_1538 = _RANDOM[12'h602];
        v0_1539 = _RANDOM[12'h603];
        v0_1540 = _RANDOM[12'h604];
        v0_1541 = _RANDOM[12'h605];
        v0_1542 = _RANDOM[12'h606];
        v0_1543 = _RANDOM[12'h607];
        v0_1544 = _RANDOM[12'h608];
        v0_1545 = _RANDOM[12'h609];
        v0_1546 = _RANDOM[12'h60A];
        v0_1547 = _RANDOM[12'h60B];
        v0_1548 = _RANDOM[12'h60C];
        v0_1549 = _RANDOM[12'h60D];
        v0_1550 = _RANDOM[12'h60E];
        v0_1551 = _RANDOM[12'h60F];
        v0_1552 = _RANDOM[12'h610];
        v0_1553 = _RANDOM[12'h611];
        v0_1554 = _RANDOM[12'h612];
        v0_1555 = _RANDOM[12'h613];
        v0_1556 = _RANDOM[12'h614];
        v0_1557 = _RANDOM[12'h615];
        v0_1558 = _RANDOM[12'h616];
        v0_1559 = _RANDOM[12'h617];
        v0_1560 = _RANDOM[12'h618];
        v0_1561 = _RANDOM[12'h619];
        v0_1562 = _RANDOM[12'h61A];
        v0_1563 = _RANDOM[12'h61B];
        v0_1564 = _RANDOM[12'h61C];
        v0_1565 = _RANDOM[12'h61D];
        v0_1566 = _RANDOM[12'h61E];
        v0_1567 = _RANDOM[12'h61F];
        v0_1568 = _RANDOM[12'h620];
        v0_1569 = _RANDOM[12'h621];
        v0_1570 = _RANDOM[12'h622];
        v0_1571 = _RANDOM[12'h623];
        v0_1572 = _RANDOM[12'h624];
        v0_1573 = _RANDOM[12'h625];
        v0_1574 = _RANDOM[12'h626];
        v0_1575 = _RANDOM[12'h627];
        v0_1576 = _RANDOM[12'h628];
        v0_1577 = _RANDOM[12'h629];
        v0_1578 = _RANDOM[12'h62A];
        v0_1579 = _RANDOM[12'h62B];
        v0_1580 = _RANDOM[12'h62C];
        v0_1581 = _RANDOM[12'h62D];
        v0_1582 = _RANDOM[12'h62E];
        v0_1583 = _RANDOM[12'h62F];
        v0_1584 = _RANDOM[12'h630];
        v0_1585 = _RANDOM[12'h631];
        v0_1586 = _RANDOM[12'h632];
        v0_1587 = _RANDOM[12'h633];
        v0_1588 = _RANDOM[12'h634];
        v0_1589 = _RANDOM[12'h635];
        v0_1590 = _RANDOM[12'h636];
        v0_1591 = _RANDOM[12'h637];
        v0_1592 = _RANDOM[12'h638];
        v0_1593 = _RANDOM[12'h639];
        v0_1594 = _RANDOM[12'h63A];
        v0_1595 = _RANDOM[12'h63B];
        v0_1596 = _RANDOM[12'h63C];
        v0_1597 = _RANDOM[12'h63D];
        v0_1598 = _RANDOM[12'h63E];
        v0_1599 = _RANDOM[12'h63F];
        v0_1600 = _RANDOM[12'h640];
        v0_1601 = _RANDOM[12'h641];
        v0_1602 = _RANDOM[12'h642];
        v0_1603 = _RANDOM[12'h643];
        v0_1604 = _RANDOM[12'h644];
        v0_1605 = _RANDOM[12'h645];
        v0_1606 = _RANDOM[12'h646];
        v0_1607 = _RANDOM[12'h647];
        v0_1608 = _RANDOM[12'h648];
        v0_1609 = _RANDOM[12'h649];
        v0_1610 = _RANDOM[12'h64A];
        v0_1611 = _RANDOM[12'h64B];
        v0_1612 = _RANDOM[12'h64C];
        v0_1613 = _RANDOM[12'h64D];
        v0_1614 = _RANDOM[12'h64E];
        v0_1615 = _RANDOM[12'h64F];
        v0_1616 = _RANDOM[12'h650];
        v0_1617 = _RANDOM[12'h651];
        v0_1618 = _RANDOM[12'h652];
        v0_1619 = _RANDOM[12'h653];
        v0_1620 = _RANDOM[12'h654];
        v0_1621 = _RANDOM[12'h655];
        v0_1622 = _RANDOM[12'h656];
        v0_1623 = _RANDOM[12'h657];
        v0_1624 = _RANDOM[12'h658];
        v0_1625 = _RANDOM[12'h659];
        v0_1626 = _RANDOM[12'h65A];
        v0_1627 = _RANDOM[12'h65B];
        v0_1628 = _RANDOM[12'h65C];
        v0_1629 = _RANDOM[12'h65D];
        v0_1630 = _RANDOM[12'h65E];
        v0_1631 = _RANDOM[12'h65F];
        v0_1632 = _RANDOM[12'h660];
        v0_1633 = _RANDOM[12'h661];
        v0_1634 = _RANDOM[12'h662];
        v0_1635 = _RANDOM[12'h663];
        v0_1636 = _RANDOM[12'h664];
        v0_1637 = _RANDOM[12'h665];
        v0_1638 = _RANDOM[12'h666];
        v0_1639 = _RANDOM[12'h667];
        v0_1640 = _RANDOM[12'h668];
        v0_1641 = _RANDOM[12'h669];
        v0_1642 = _RANDOM[12'h66A];
        v0_1643 = _RANDOM[12'h66B];
        v0_1644 = _RANDOM[12'h66C];
        v0_1645 = _RANDOM[12'h66D];
        v0_1646 = _RANDOM[12'h66E];
        v0_1647 = _RANDOM[12'h66F];
        v0_1648 = _RANDOM[12'h670];
        v0_1649 = _RANDOM[12'h671];
        v0_1650 = _RANDOM[12'h672];
        v0_1651 = _RANDOM[12'h673];
        v0_1652 = _RANDOM[12'h674];
        v0_1653 = _RANDOM[12'h675];
        v0_1654 = _RANDOM[12'h676];
        v0_1655 = _RANDOM[12'h677];
        v0_1656 = _RANDOM[12'h678];
        v0_1657 = _RANDOM[12'h679];
        v0_1658 = _RANDOM[12'h67A];
        v0_1659 = _RANDOM[12'h67B];
        v0_1660 = _RANDOM[12'h67C];
        v0_1661 = _RANDOM[12'h67D];
        v0_1662 = _RANDOM[12'h67E];
        v0_1663 = _RANDOM[12'h67F];
        v0_1664 = _RANDOM[12'h680];
        v0_1665 = _RANDOM[12'h681];
        v0_1666 = _RANDOM[12'h682];
        v0_1667 = _RANDOM[12'h683];
        v0_1668 = _RANDOM[12'h684];
        v0_1669 = _RANDOM[12'h685];
        v0_1670 = _RANDOM[12'h686];
        v0_1671 = _RANDOM[12'h687];
        v0_1672 = _RANDOM[12'h688];
        v0_1673 = _RANDOM[12'h689];
        v0_1674 = _RANDOM[12'h68A];
        v0_1675 = _RANDOM[12'h68B];
        v0_1676 = _RANDOM[12'h68C];
        v0_1677 = _RANDOM[12'h68D];
        v0_1678 = _RANDOM[12'h68E];
        v0_1679 = _RANDOM[12'h68F];
        v0_1680 = _RANDOM[12'h690];
        v0_1681 = _RANDOM[12'h691];
        v0_1682 = _RANDOM[12'h692];
        v0_1683 = _RANDOM[12'h693];
        v0_1684 = _RANDOM[12'h694];
        v0_1685 = _RANDOM[12'h695];
        v0_1686 = _RANDOM[12'h696];
        v0_1687 = _RANDOM[12'h697];
        v0_1688 = _RANDOM[12'h698];
        v0_1689 = _RANDOM[12'h699];
        v0_1690 = _RANDOM[12'h69A];
        v0_1691 = _RANDOM[12'h69B];
        v0_1692 = _RANDOM[12'h69C];
        v0_1693 = _RANDOM[12'h69D];
        v0_1694 = _RANDOM[12'h69E];
        v0_1695 = _RANDOM[12'h69F];
        v0_1696 = _RANDOM[12'h6A0];
        v0_1697 = _RANDOM[12'h6A1];
        v0_1698 = _RANDOM[12'h6A2];
        v0_1699 = _RANDOM[12'h6A3];
        v0_1700 = _RANDOM[12'h6A4];
        v0_1701 = _RANDOM[12'h6A5];
        v0_1702 = _RANDOM[12'h6A6];
        v0_1703 = _RANDOM[12'h6A7];
        v0_1704 = _RANDOM[12'h6A8];
        v0_1705 = _RANDOM[12'h6A9];
        v0_1706 = _RANDOM[12'h6AA];
        v0_1707 = _RANDOM[12'h6AB];
        v0_1708 = _RANDOM[12'h6AC];
        v0_1709 = _RANDOM[12'h6AD];
        v0_1710 = _RANDOM[12'h6AE];
        v0_1711 = _RANDOM[12'h6AF];
        v0_1712 = _RANDOM[12'h6B0];
        v0_1713 = _RANDOM[12'h6B1];
        v0_1714 = _RANDOM[12'h6B2];
        v0_1715 = _RANDOM[12'h6B3];
        v0_1716 = _RANDOM[12'h6B4];
        v0_1717 = _RANDOM[12'h6B5];
        v0_1718 = _RANDOM[12'h6B6];
        v0_1719 = _RANDOM[12'h6B7];
        v0_1720 = _RANDOM[12'h6B8];
        v0_1721 = _RANDOM[12'h6B9];
        v0_1722 = _RANDOM[12'h6BA];
        v0_1723 = _RANDOM[12'h6BB];
        v0_1724 = _RANDOM[12'h6BC];
        v0_1725 = _RANDOM[12'h6BD];
        v0_1726 = _RANDOM[12'h6BE];
        v0_1727 = _RANDOM[12'h6BF];
        v0_1728 = _RANDOM[12'h6C0];
        v0_1729 = _RANDOM[12'h6C1];
        v0_1730 = _RANDOM[12'h6C2];
        v0_1731 = _RANDOM[12'h6C3];
        v0_1732 = _RANDOM[12'h6C4];
        v0_1733 = _RANDOM[12'h6C5];
        v0_1734 = _RANDOM[12'h6C6];
        v0_1735 = _RANDOM[12'h6C7];
        v0_1736 = _RANDOM[12'h6C8];
        v0_1737 = _RANDOM[12'h6C9];
        v0_1738 = _RANDOM[12'h6CA];
        v0_1739 = _RANDOM[12'h6CB];
        v0_1740 = _RANDOM[12'h6CC];
        v0_1741 = _RANDOM[12'h6CD];
        v0_1742 = _RANDOM[12'h6CE];
        v0_1743 = _RANDOM[12'h6CF];
        v0_1744 = _RANDOM[12'h6D0];
        v0_1745 = _RANDOM[12'h6D1];
        v0_1746 = _RANDOM[12'h6D2];
        v0_1747 = _RANDOM[12'h6D3];
        v0_1748 = _RANDOM[12'h6D4];
        v0_1749 = _RANDOM[12'h6D5];
        v0_1750 = _RANDOM[12'h6D6];
        v0_1751 = _RANDOM[12'h6D7];
        v0_1752 = _RANDOM[12'h6D8];
        v0_1753 = _RANDOM[12'h6D9];
        v0_1754 = _RANDOM[12'h6DA];
        v0_1755 = _RANDOM[12'h6DB];
        v0_1756 = _RANDOM[12'h6DC];
        v0_1757 = _RANDOM[12'h6DD];
        v0_1758 = _RANDOM[12'h6DE];
        v0_1759 = _RANDOM[12'h6DF];
        v0_1760 = _RANDOM[12'h6E0];
        v0_1761 = _RANDOM[12'h6E1];
        v0_1762 = _RANDOM[12'h6E2];
        v0_1763 = _RANDOM[12'h6E3];
        v0_1764 = _RANDOM[12'h6E4];
        v0_1765 = _RANDOM[12'h6E5];
        v0_1766 = _RANDOM[12'h6E6];
        v0_1767 = _RANDOM[12'h6E7];
        v0_1768 = _RANDOM[12'h6E8];
        v0_1769 = _RANDOM[12'h6E9];
        v0_1770 = _RANDOM[12'h6EA];
        v0_1771 = _RANDOM[12'h6EB];
        v0_1772 = _RANDOM[12'h6EC];
        v0_1773 = _RANDOM[12'h6ED];
        v0_1774 = _RANDOM[12'h6EE];
        v0_1775 = _RANDOM[12'h6EF];
        v0_1776 = _RANDOM[12'h6F0];
        v0_1777 = _RANDOM[12'h6F1];
        v0_1778 = _RANDOM[12'h6F2];
        v0_1779 = _RANDOM[12'h6F3];
        v0_1780 = _RANDOM[12'h6F4];
        v0_1781 = _RANDOM[12'h6F5];
        v0_1782 = _RANDOM[12'h6F6];
        v0_1783 = _RANDOM[12'h6F7];
        v0_1784 = _RANDOM[12'h6F8];
        v0_1785 = _RANDOM[12'h6F9];
        v0_1786 = _RANDOM[12'h6FA];
        v0_1787 = _RANDOM[12'h6FB];
        v0_1788 = _RANDOM[12'h6FC];
        v0_1789 = _RANDOM[12'h6FD];
        v0_1790 = _RANDOM[12'h6FE];
        v0_1791 = _RANDOM[12'h6FF];
        v0_1792 = _RANDOM[12'h700];
        v0_1793 = _RANDOM[12'h701];
        v0_1794 = _RANDOM[12'h702];
        v0_1795 = _RANDOM[12'h703];
        v0_1796 = _RANDOM[12'h704];
        v0_1797 = _RANDOM[12'h705];
        v0_1798 = _RANDOM[12'h706];
        v0_1799 = _RANDOM[12'h707];
        v0_1800 = _RANDOM[12'h708];
        v0_1801 = _RANDOM[12'h709];
        v0_1802 = _RANDOM[12'h70A];
        v0_1803 = _RANDOM[12'h70B];
        v0_1804 = _RANDOM[12'h70C];
        v0_1805 = _RANDOM[12'h70D];
        v0_1806 = _RANDOM[12'h70E];
        v0_1807 = _RANDOM[12'h70F];
        v0_1808 = _RANDOM[12'h710];
        v0_1809 = _RANDOM[12'h711];
        v0_1810 = _RANDOM[12'h712];
        v0_1811 = _RANDOM[12'h713];
        v0_1812 = _RANDOM[12'h714];
        v0_1813 = _RANDOM[12'h715];
        v0_1814 = _RANDOM[12'h716];
        v0_1815 = _RANDOM[12'h717];
        v0_1816 = _RANDOM[12'h718];
        v0_1817 = _RANDOM[12'h719];
        v0_1818 = _RANDOM[12'h71A];
        v0_1819 = _RANDOM[12'h71B];
        v0_1820 = _RANDOM[12'h71C];
        v0_1821 = _RANDOM[12'h71D];
        v0_1822 = _RANDOM[12'h71E];
        v0_1823 = _RANDOM[12'h71F];
        v0_1824 = _RANDOM[12'h720];
        v0_1825 = _RANDOM[12'h721];
        v0_1826 = _RANDOM[12'h722];
        v0_1827 = _RANDOM[12'h723];
        v0_1828 = _RANDOM[12'h724];
        v0_1829 = _RANDOM[12'h725];
        v0_1830 = _RANDOM[12'h726];
        v0_1831 = _RANDOM[12'h727];
        v0_1832 = _RANDOM[12'h728];
        v0_1833 = _RANDOM[12'h729];
        v0_1834 = _RANDOM[12'h72A];
        v0_1835 = _RANDOM[12'h72B];
        v0_1836 = _RANDOM[12'h72C];
        v0_1837 = _RANDOM[12'h72D];
        v0_1838 = _RANDOM[12'h72E];
        v0_1839 = _RANDOM[12'h72F];
        v0_1840 = _RANDOM[12'h730];
        v0_1841 = _RANDOM[12'h731];
        v0_1842 = _RANDOM[12'h732];
        v0_1843 = _RANDOM[12'h733];
        v0_1844 = _RANDOM[12'h734];
        v0_1845 = _RANDOM[12'h735];
        v0_1846 = _RANDOM[12'h736];
        v0_1847 = _RANDOM[12'h737];
        v0_1848 = _RANDOM[12'h738];
        v0_1849 = _RANDOM[12'h739];
        v0_1850 = _RANDOM[12'h73A];
        v0_1851 = _RANDOM[12'h73B];
        v0_1852 = _RANDOM[12'h73C];
        v0_1853 = _RANDOM[12'h73D];
        v0_1854 = _RANDOM[12'h73E];
        v0_1855 = _RANDOM[12'h73F];
        v0_1856 = _RANDOM[12'h740];
        v0_1857 = _RANDOM[12'h741];
        v0_1858 = _RANDOM[12'h742];
        v0_1859 = _RANDOM[12'h743];
        v0_1860 = _RANDOM[12'h744];
        v0_1861 = _RANDOM[12'h745];
        v0_1862 = _RANDOM[12'h746];
        v0_1863 = _RANDOM[12'h747];
        v0_1864 = _RANDOM[12'h748];
        v0_1865 = _RANDOM[12'h749];
        v0_1866 = _RANDOM[12'h74A];
        v0_1867 = _RANDOM[12'h74B];
        v0_1868 = _RANDOM[12'h74C];
        v0_1869 = _RANDOM[12'h74D];
        v0_1870 = _RANDOM[12'h74E];
        v0_1871 = _RANDOM[12'h74F];
        v0_1872 = _RANDOM[12'h750];
        v0_1873 = _RANDOM[12'h751];
        v0_1874 = _RANDOM[12'h752];
        v0_1875 = _RANDOM[12'h753];
        v0_1876 = _RANDOM[12'h754];
        v0_1877 = _RANDOM[12'h755];
        v0_1878 = _RANDOM[12'h756];
        v0_1879 = _RANDOM[12'h757];
        v0_1880 = _RANDOM[12'h758];
        v0_1881 = _RANDOM[12'h759];
        v0_1882 = _RANDOM[12'h75A];
        v0_1883 = _RANDOM[12'h75B];
        v0_1884 = _RANDOM[12'h75C];
        v0_1885 = _RANDOM[12'h75D];
        v0_1886 = _RANDOM[12'h75E];
        v0_1887 = _RANDOM[12'h75F];
        v0_1888 = _RANDOM[12'h760];
        v0_1889 = _RANDOM[12'h761];
        v0_1890 = _RANDOM[12'h762];
        v0_1891 = _RANDOM[12'h763];
        v0_1892 = _RANDOM[12'h764];
        v0_1893 = _RANDOM[12'h765];
        v0_1894 = _RANDOM[12'h766];
        v0_1895 = _RANDOM[12'h767];
        v0_1896 = _RANDOM[12'h768];
        v0_1897 = _RANDOM[12'h769];
        v0_1898 = _RANDOM[12'h76A];
        v0_1899 = _RANDOM[12'h76B];
        v0_1900 = _RANDOM[12'h76C];
        v0_1901 = _RANDOM[12'h76D];
        v0_1902 = _RANDOM[12'h76E];
        v0_1903 = _RANDOM[12'h76F];
        v0_1904 = _RANDOM[12'h770];
        v0_1905 = _RANDOM[12'h771];
        v0_1906 = _RANDOM[12'h772];
        v0_1907 = _RANDOM[12'h773];
        v0_1908 = _RANDOM[12'h774];
        v0_1909 = _RANDOM[12'h775];
        v0_1910 = _RANDOM[12'h776];
        v0_1911 = _RANDOM[12'h777];
        v0_1912 = _RANDOM[12'h778];
        v0_1913 = _RANDOM[12'h779];
        v0_1914 = _RANDOM[12'h77A];
        v0_1915 = _RANDOM[12'h77B];
        v0_1916 = _RANDOM[12'h77C];
        v0_1917 = _RANDOM[12'h77D];
        v0_1918 = _RANDOM[12'h77E];
        v0_1919 = _RANDOM[12'h77F];
        v0_1920 = _RANDOM[12'h780];
        v0_1921 = _RANDOM[12'h781];
        v0_1922 = _RANDOM[12'h782];
        v0_1923 = _RANDOM[12'h783];
        v0_1924 = _RANDOM[12'h784];
        v0_1925 = _RANDOM[12'h785];
        v0_1926 = _RANDOM[12'h786];
        v0_1927 = _RANDOM[12'h787];
        v0_1928 = _RANDOM[12'h788];
        v0_1929 = _RANDOM[12'h789];
        v0_1930 = _RANDOM[12'h78A];
        v0_1931 = _RANDOM[12'h78B];
        v0_1932 = _RANDOM[12'h78C];
        v0_1933 = _RANDOM[12'h78D];
        v0_1934 = _RANDOM[12'h78E];
        v0_1935 = _RANDOM[12'h78F];
        v0_1936 = _RANDOM[12'h790];
        v0_1937 = _RANDOM[12'h791];
        v0_1938 = _RANDOM[12'h792];
        v0_1939 = _RANDOM[12'h793];
        v0_1940 = _RANDOM[12'h794];
        v0_1941 = _RANDOM[12'h795];
        v0_1942 = _RANDOM[12'h796];
        v0_1943 = _RANDOM[12'h797];
        v0_1944 = _RANDOM[12'h798];
        v0_1945 = _RANDOM[12'h799];
        v0_1946 = _RANDOM[12'h79A];
        v0_1947 = _RANDOM[12'h79B];
        v0_1948 = _RANDOM[12'h79C];
        v0_1949 = _RANDOM[12'h79D];
        v0_1950 = _RANDOM[12'h79E];
        v0_1951 = _RANDOM[12'h79F];
        v0_1952 = _RANDOM[12'h7A0];
        v0_1953 = _RANDOM[12'h7A1];
        v0_1954 = _RANDOM[12'h7A2];
        v0_1955 = _RANDOM[12'h7A3];
        v0_1956 = _RANDOM[12'h7A4];
        v0_1957 = _RANDOM[12'h7A5];
        v0_1958 = _RANDOM[12'h7A6];
        v0_1959 = _RANDOM[12'h7A7];
        v0_1960 = _RANDOM[12'h7A8];
        v0_1961 = _RANDOM[12'h7A9];
        v0_1962 = _RANDOM[12'h7AA];
        v0_1963 = _RANDOM[12'h7AB];
        v0_1964 = _RANDOM[12'h7AC];
        v0_1965 = _RANDOM[12'h7AD];
        v0_1966 = _RANDOM[12'h7AE];
        v0_1967 = _RANDOM[12'h7AF];
        v0_1968 = _RANDOM[12'h7B0];
        v0_1969 = _RANDOM[12'h7B1];
        v0_1970 = _RANDOM[12'h7B2];
        v0_1971 = _RANDOM[12'h7B3];
        v0_1972 = _RANDOM[12'h7B4];
        v0_1973 = _RANDOM[12'h7B5];
        v0_1974 = _RANDOM[12'h7B6];
        v0_1975 = _RANDOM[12'h7B7];
        v0_1976 = _RANDOM[12'h7B8];
        v0_1977 = _RANDOM[12'h7B9];
        v0_1978 = _RANDOM[12'h7BA];
        v0_1979 = _RANDOM[12'h7BB];
        v0_1980 = _RANDOM[12'h7BC];
        v0_1981 = _RANDOM[12'h7BD];
        v0_1982 = _RANDOM[12'h7BE];
        v0_1983 = _RANDOM[12'h7BF];
        v0_1984 = _RANDOM[12'h7C0];
        v0_1985 = _RANDOM[12'h7C1];
        v0_1986 = _RANDOM[12'h7C2];
        v0_1987 = _RANDOM[12'h7C3];
        v0_1988 = _RANDOM[12'h7C4];
        v0_1989 = _RANDOM[12'h7C5];
        v0_1990 = _RANDOM[12'h7C6];
        v0_1991 = _RANDOM[12'h7C7];
        v0_1992 = _RANDOM[12'h7C8];
        v0_1993 = _RANDOM[12'h7C9];
        v0_1994 = _RANDOM[12'h7CA];
        v0_1995 = _RANDOM[12'h7CB];
        v0_1996 = _RANDOM[12'h7CC];
        v0_1997 = _RANDOM[12'h7CD];
        v0_1998 = _RANDOM[12'h7CE];
        v0_1999 = _RANDOM[12'h7CF];
        v0_2000 = _RANDOM[12'h7D0];
        v0_2001 = _RANDOM[12'h7D1];
        v0_2002 = _RANDOM[12'h7D2];
        v0_2003 = _RANDOM[12'h7D3];
        v0_2004 = _RANDOM[12'h7D4];
        v0_2005 = _RANDOM[12'h7D5];
        v0_2006 = _RANDOM[12'h7D6];
        v0_2007 = _RANDOM[12'h7D7];
        v0_2008 = _RANDOM[12'h7D8];
        v0_2009 = _RANDOM[12'h7D9];
        v0_2010 = _RANDOM[12'h7DA];
        v0_2011 = _RANDOM[12'h7DB];
        v0_2012 = _RANDOM[12'h7DC];
        v0_2013 = _RANDOM[12'h7DD];
        v0_2014 = _RANDOM[12'h7DE];
        v0_2015 = _RANDOM[12'h7DF];
        v0_2016 = _RANDOM[12'h7E0];
        v0_2017 = _RANDOM[12'h7E1];
        v0_2018 = _RANDOM[12'h7E2];
        v0_2019 = _RANDOM[12'h7E3];
        v0_2020 = _RANDOM[12'h7E4];
        v0_2021 = _RANDOM[12'h7E5];
        v0_2022 = _RANDOM[12'h7E6];
        v0_2023 = _RANDOM[12'h7E7];
        v0_2024 = _RANDOM[12'h7E8];
        v0_2025 = _RANDOM[12'h7E9];
        v0_2026 = _RANDOM[12'h7EA];
        v0_2027 = _RANDOM[12'h7EB];
        v0_2028 = _RANDOM[12'h7EC];
        v0_2029 = _RANDOM[12'h7ED];
        v0_2030 = _RANDOM[12'h7EE];
        v0_2031 = _RANDOM[12'h7EF];
        v0_2032 = _RANDOM[12'h7F0];
        v0_2033 = _RANDOM[12'h7F1];
        v0_2034 = _RANDOM[12'h7F2];
        v0_2035 = _RANDOM[12'h7F3];
        v0_2036 = _RANDOM[12'h7F4];
        v0_2037 = _RANDOM[12'h7F5];
        v0_2038 = _RANDOM[12'h7F6];
        v0_2039 = _RANDOM[12'h7F7];
        v0_2040 = _RANDOM[12'h7F8];
        v0_2041 = _RANDOM[12'h7F9];
        v0_2042 = _RANDOM[12'h7FA];
        v0_2043 = _RANDOM[12'h7FB];
        v0_2044 = _RANDOM[12'h7FC];
        v0_2045 = _RANDOM[12'h7FD];
        v0_2046 = _RANDOM[12'h7FE];
        v0_2047 = _RANDOM[12'h7FF];
        queueCount_0 = _RANDOM[12'h800][6:0];
        queueCount_1 = _RANDOM[12'h800][13:7];
        queueCount_2 = _RANDOM[12'h800][20:14];
        queueCount_3 = _RANDOM[12'h800][27:21];
        queueCount_4 = {_RANDOM[12'h800][31:28], _RANDOM[12'h801][2:0]};
        queueCount_5 = _RANDOM[12'h801][9:3];
        queueCount_6 = _RANDOM[12'h801][16:10];
        queueCount_7 = _RANDOM[12'h801][23:17];
        queueCount_0_1 = _RANDOM[12'h801][30:24];
        queueCount_1_1 = {_RANDOM[12'h801][31], _RANDOM[12'h802][5:0]};
        queueCount_2_1 = _RANDOM[12'h802][12:6];
        queueCount_3_1 = _RANDOM[12'h802][19:13];
        queueCount_4_1 = _RANDOM[12'h802][26:20];
        queueCount_5_1 = {_RANDOM[12'h802][31:27], _RANDOM[12'h803][1:0]};
        queueCount_6_1 = _RANDOM[12'h803][8:2];
        queueCount_7_1 = _RANDOM[12'h803][15:9];
        queueCount_0_2 = _RANDOM[12'h803][22:16];
        queueCount_1_2 = _RANDOM[12'h803][29:23];
        queueCount_2_2 = {_RANDOM[12'h803][31:30], _RANDOM[12'h804][4:0]};
        queueCount_3_2 = _RANDOM[12'h804][11:5];
        queueCount_4_2 = _RANDOM[12'h804][18:12];
        queueCount_5_2 = _RANDOM[12'h804][25:19];
        queueCount_6_2 = {_RANDOM[12'h804][31:26], _RANDOM[12'h805][0]};
        queueCount_7_2 = _RANDOM[12'h805][7:1];
        queueCount_0_3 = _RANDOM[12'h805][14:8];
        queueCount_1_3 = _RANDOM[12'h805][21:15];
        queueCount_2_3 = _RANDOM[12'h805][28:22];
        queueCount_3_3 = {_RANDOM[12'h805][31:29], _RANDOM[12'h806][3:0]};
        queueCount_4_3 = _RANDOM[12'h806][10:4];
        queueCount_5_3 = _RANDOM[12'h806][17:11];
        queueCount_6_3 = _RANDOM[12'h806][24:18];
        queueCount_7_3 = _RANDOM[12'h806][31:25];
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  wire [12:0]         sourceQueue_deq_bits;
  wire [31:0]         axi4Port_aw_bits_addr_0;
  assign axi4Port_aw_bits_addr_0 = _storeUnit_memRequest_bits_address;
  assign dataQueue_enq_bits_index = _storeUnit_memRequest_bits_index;
  assign dataQueue_enq_bits_address = _storeUnit_memRequest_bits_address;
  wire [6:0]          simpleSourceQueue_deq_bits;
  wire [31:0]         simpleAccessPorts_aw_bits_addr_0;
  assign simpleAccessPorts_aw_bits_addr_0 = _otherUnit_memWriteRequest_bits_address;
  wire [3:0]          otherUnitTargetQueue_enq_bits;
  assign otherUnitTargetQueue_enq_bits = _otherUnit_status_targetLane;
  assign simpleDataQueue_enq_bits_source = _otherUnit_memWriteRequest_bits_source;
  assign simpleDataQueue_enq_bits_address = _otherUnit_memWriteRequest_bits_address;
  assign simpleDataQueue_enq_bits_size = _otherUnit_memWriteRequest_bits_size;
  wire                writeQueueVec_0_empty;
  assign writeQueueVec_0_empty = _writeQueueVec_fifo_empty;
  wire                writeQueueVec_0_full;
  assign writeQueueVec_0_full = _writeQueueVec_fifo_full;
  wire                writeQueueVec_1_empty;
  assign writeQueueVec_1_empty = _writeQueueVec_fifo_1_empty;
  wire                writeQueueVec_1_full;
  assign writeQueueVec_1_full = _writeQueueVec_fifo_1_full;
  wire                writeQueueVec_2_empty;
  assign writeQueueVec_2_empty = _writeQueueVec_fifo_2_empty;
  wire                writeQueueVec_2_full;
  assign writeQueueVec_2_full = _writeQueueVec_fifo_2_full;
  wire                writeQueueVec_3_empty;
  assign writeQueueVec_3_empty = _writeQueueVec_fifo_3_empty;
  wire                writeQueueVec_3_full;
  assign writeQueueVec_3_full = _writeQueueVec_fifo_3_full;
  assign otherUnitTargetQueue_empty = _otherUnitTargetQueue_fifo_empty;
  wire                otherUnitTargetQueue_full;
  assign otherUnitTargetQueue_full = _otherUnitTargetQueue_fifo_full;
  wire                otherUnitDataQueueVec_0_empty;
  assign otherUnitDataQueueVec_0_empty = _otherUnitDataQueueVec_fifo_empty;
  wire                otherUnitDataQueueVec_0_full;
  assign otherUnitDataQueueVec_0_full = _otherUnitDataQueueVec_fifo_full;
  wire                otherUnitDataQueueVec_1_empty;
  assign otherUnitDataQueueVec_1_empty = _otherUnitDataQueueVec_fifo_1_empty;
  wire                otherUnitDataQueueVec_1_full;
  assign otherUnitDataQueueVec_1_full = _otherUnitDataQueueVec_fifo_1_full;
  wire                otherUnitDataQueueVec_2_empty;
  assign otherUnitDataQueueVec_2_empty = _otherUnitDataQueueVec_fifo_2_empty;
  wire                otherUnitDataQueueVec_2_full;
  assign otherUnitDataQueueVec_2_full = _otherUnitDataQueueVec_fifo_2_full;
  wire                otherUnitDataQueueVec_3_empty;
  assign otherUnitDataQueueVec_3_empty = _otherUnitDataQueueVec_fifo_3_empty;
  wire                otherUnitDataQueueVec_3_full;
  assign otherUnitDataQueueVec_3_full = _otherUnitDataQueueVec_fifo_3_full;
  wire                writeIndexQueue_empty;
  assign writeIndexQueue_empty = _writeIndexQueue_fifo_empty;
  wire                writeIndexQueue_full;
  assign writeIndexQueue_full = _writeIndexQueue_fifo_full;
  wire                writeIndexQueue_1_empty;
  assign writeIndexQueue_1_empty = _writeIndexQueue_fifo_1_empty;
  wire                writeIndexQueue_1_full;
  assign writeIndexQueue_1_full = _writeIndexQueue_fifo_1_full;
  wire                writeIndexQueue_2_empty;
  assign writeIndexQueue_2_empty = _writeIndexQueue_fifo_2_empty;
  wire                writeIndexQueue_2_full;
  assign writeIndexQueue_2_full = _writeIndexQueue_fifo_2_full;
  wire                writeIndexQueue_3_empty;
  assign writeIndexQueue_3_empty = _writeIndexQueue_fifo_3_empty;
  wire                writeIndexQueue_3_full;
  assign writeIndexQueue_3_full = _writeIndexQueue_fifo_3_full;
  wire                sourceQueue_empty;
  assign sourceQueue_empty = _sourceQueue_fifo_empty;
  wire                sourceQueue_full;
  assign sourceQueue_full = _sourceQueue_fifo_full;
  wire                dataQueue_empty;
  assign dataQueue_empty = _dataQueue_fifo_empty;
  wire                dataQueue_full;
  assign dataQueue_full = _dataQueue_fifo_full;
  wire                simpleSourceQueue_empty;
  assign simpleSourceQueue_empty = _simpleSourceQueue_fifo_empty;
  wire                simpleSourceQueue_full;
  assign simpleSourceQueue_full = _simpleSourceQueue_fifo_full;
  wire                simpleDataQueue_empty;
  assign simpleDataQueue_empty = _simpleDataQueue_fifo_empty;
  wire                simpleDataQueue_full;
  assign simpleDataQueue_full = _simpleDataQueue_fifo_full;
  LoadUnit loadUnit (
    .clock                                                  (clock),
    .reset                                                  (reset),
    .lsuRequest_valid                                       (reqEnq_0),
    .lsuRequest_bits_instructionInformation_nf              (request_bits_instructionInformation_nf_0),
    .lsuRequest_bits_instructionInformation_mew             (request_bits_instructionInformation_mew_0),
    .lsuRequest_bits_instructionInformation_mop             (request_bits_instructionInformation_mop_0),
    .lsuRequest_bits_instructionInformation_lumop           (request_bits_instructionInformation_lumop_0),
    .lsuRequest_bits_instructionInformation_eew             (request_bits_instructionInformation_eew_0),
    .lsuRequest_bits_instructionInformation_vs3             (request_bits_instructionInformation_vs3_0),
    .lsuRequest_bits_instructionInformation_isStore         (request_bits_instructionInformation_isStore_0),
    .lsuRequest_bits_instructionInformation_maskedLoadStore (request_bits_instructionInformation_maskedLoadStore_0),
    .lsuRequest_bits_rs1Data                                (request_bits_rs1Data_0),
    .lsuRequest_bits_rs2Data                                (request_bits_rs2Data_0),
    .lsuRequest_bits_instructionIndex                       (request_bits_instructionIndex_0),
    .csrInterface_vl                                        (csrInterface_vl),
    .csrInterface_vStart                                    (csrInterface_vStart),
    .csrInterface_vlmul                                     (csrInterface_vlmul),
    .csrInterface_vSew                                      (csrInterface_vSew),
    .csrInterface_vxrm                                      (csrInterface_vxrm),
    .csrInterface_vta                                       (csrInterface_vta),
    .csrInterface_vma                                       (csrInterface_vma),
    .maskInput                                              (_GEN_1023[maskSelect]),
    .maskSelect_valid                                       (_loadUnit_maskSelect_valid),
    .maskSelect_bits                                        (_loadUnit_maskSelect_bits),
    .addressConflict                                        (stallLoad),
    .memRequest_ready                                       (sourceQueue_enq_ready & axi4Port_ar_ready_0),
    .memRequest_valid                                       (_loadUnit_memRequest_valid),
    .memRequest_bits_src                                    (sourceQueue_enq_bits),
    .memRequest_bits_address                                (axi4Port_ar_bits_addr_0),
    .memResponse_ready                                      (axi4Port_r_ready_0),
    .memResponse_valid                                      (axi4Port_r_valid_0),
    .memResponse_bits_data                                  (axi4Port_r_bits_data_0),
    .memResponse_bits_index                                 (sourceQueue_deq_bits),
    .status_idle                                            (_loadUnit_status_idle),
    .status_last                                            (_loadUnit_status_last),
    .status_instructionIndex                                (_loadUnit_status_instructionIndex),
    .status_changeMaskGroup                                 (/* unused */),
    .status_startAddress                                    (_loadUnit_status_startAddress),
    .status_endAddress                                      (_loadUnit_status_endAddress),
    .vrfWritePort_0_ready                                   (writeQueueVec_0_enq_ready & ~(otherTryToWrite[0])),
    .vrfWritePort_0_valid                                   (_loadUnit_vrfWritePort_0_valid),
    .vrfWritePort_0_bits_vd                                 (_loadUnit_vrfWritePort_0_bits_vd),
    .vrfWritePort_0_bits_offset                             (_loadUnit_vrfWritePort_0_bits_offset),
    .vrfWritePort_0_bits_mask                               (_loadUnit_vrfWritePort_0_bits_mask),
    .vrfWritePort_0_bits_data                               (_loadUnit_vrfWritePort_0_bits_data),
    .vrfWritePort_0_bits_instructionIndex                   (_loadUnit_vrfWritePort_0_bits_instructionIndex),
    .vrfWritePort_1_ready                                   (writeQueueVec_1_enq_ready & ~(otherTryToWrite[1])),
    .vrfWritePort_1_valid                                   (_loadUnit_vrfWritePort_1_valid),
    .vrfWritePort_1_bits_vd                                 (_loadUnit_vrfWritePort_1_bits_vd),
    .vrfWritePort_1_bits_offset                             (_loadUnit_vrfWritePort_1_bits_offset),
    .vrfWritePort_1_bits_mask                               (_loadUnit_vrfWritePort_1_bits_mask),
    .vrfWritePort_1_bits_data                               (_loadUnit_vrfWritePort_1_bits_data),
    .vrfWritePort_1_bits_instructionIndex                   (_loadUnit_vrfWritePort_1_bits_instructionIndex),
    .vrfWritePort_2_ready                                   (writeQueueVec_2_enq_ready & ~(otherTryToWrite[2])),
    .vrfWritePort_2_valid                                   (_loadUnit_vrfWritePort_2_valid),
    .vrfWritePort_2_bits_vd                                 (_loadUnit_vrfWritePort_2_bits_vd),
    .vrfWritePort_2_bits_offset                             (_loadUnit_vrfWritePort_2_bits_offset),
    .vrfWritePort_2_bits_mask                               (_loadUnit_vrfWritePort_2_bits_mask),
    .vrfWritePort_2_bits_data                               (_loadUnit_vrfWritePort_2_bits_data),
    .vrfWritePort_2_bits_instructionIndex                   (_loadUnit_vrfWritePort_2_bits_instructionIndex),
    .vrfWritePort_3_ready                                   (writeQueueVec_3_enq_ready & ~(otherTryToWrite[3])),
    .vrfWritePort_3_valid                                   (_loadUnit_vrfWritePort_3_valid),
    .vrfWritePort_3_bits_vd                                 (_loadUnit_vrfWritePort_3_bits_vd),
    .vrfWritePort_3_bits_offset                             (_loadUnit_vrfWritePort_3_bits_offset),
    .vrfWritePort_3_bits_mask                               (_loadUnit_vrfWritePort_3_bits_mask),
    .vrfWritePort_3_bits_data                               (_loadUnit_vrfWritePort_3_bits_data),
    .vrfWritePort_3_bits_instructionIndex                   (_loadUnit_vrfWritePort_3_bits_instructionIndex)
  );
  StoreUnit storeUnit (
    .clock                                                  (clock),
    .reset                                                  (reset),
    .lsuRequest_valid                                       (reqEnq_1),
    .lsuRequest_bits_instructionInformation_nf              (request_bits_instructionInformation_nf_0),
    .lsuRequest_bits_instructionInformation_mew             (request_bits_instructionInformation_mew_0),
    .lsuRequest_bits_instructionInformation_mop             (request_bits_instructionInformation_mop_0),
    .lsuRequest_bits_instructionInformation_lumop           (request_bits_instructionInformation_lumop_0),
    .lsuRequest_bits_instructionInformation_eew             (request_bits_instructionInformation_eew_0),
    .lsuRequest_bits_instructionInformation_vs3             (request_bits_instructionInformation_vs3_0),
    .lsuRequest_bits_instructionInformation_isStore         (request_bits_instructionInformation_isStore_0),
    .lsuRequest_bits_instructionInformation_maskedLoadStore (request_bits_instructionInformation_maskedLoadStore_0),
    .lsuRequest_bits_rs1Data                                (request_bits_rs1Data_0),
    .lsuRequest_bits_rs2Data                                (request_bits_rs2Data_0),
    .lsuRequest_bits_instructionIndex                       (request_bits_instructionIndex_0),
    .csrInterface_vl                                        (csrInterface_vl),
    .csrInterface_vStart                                    (csrInterface_vStart),
    .csrInterface_vlmul                                     (csrInterface_vlmul),
    .csrInterface_vSew                                      (csrInterface_vSew),
    .csrInterface_vxrm                                      (csrInterface_vxrm),
    .csrInterface_vta                                       (csrInterface_vta),
    .csrInterface_vma                                       (csrInterface_vma),
    .maskInput                                              (_GEN_1024[maskSelect_1]),
    .maskSelect_valid                                       (_storeUnit_maskSelect_valid),
    .maskSelect_bits                                        (_storeUnit_maskSelect_bits),
    .memRequest_ready                                       (axi4Port_aw_ready_0 & dataQueue_enq_ready),
    .memRequest_valid                                       (_storeUnit_memRequest_valid),
    .memRequest_bits_data                                   (dataQueue_enq_bits_data),
    .memRequest_bits_mask                                   (dataQueue_enq_bits_mask),
    .memRequest_bits_index                                  (_storeUnit_memRequest_bits_index),
    .memRequest_bits_address                                (_storeUnit_memRequest_bits_address),
    .status_idle                                            (_storeUnit_status_idle),
    .status_last                                            (_storeUnit_status_last),
    .status_instructionIndex                                (_storeUnit_status_instructionIndex),
    .status_changeMaskGroup                                 (/* unused */),
    .status_startAddress                                    (_storeUnit_status_startAddress),
    .status_endAddress                                      (_storeUnit_status_endAddress),
    .vrfReadDataPorts_0_ready                               (vrfReadDataPorts_0_ready_0 & ~(otherTryReadVrf[0])),
    .vrfReadDataPorts_0_valid                               (_storeUnit_vrfReadDataPorts_0_valid),
    .vrfReadDataPorts_0_bits_vs                             (_storeUnit_vrfReadDataPorts_0_bits_vs),
    .vrfReadDataPorts_0_bits_offset                         (_storeUnit_vrfReadDataPorts_0_bits_offset),
    .vrfReadDataPorts_0_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_0_bits_instructionIndex),
    .vrfReadDataPorts_1_ready                               (vrfReadDataPorts_1_ready_0 & ~(otherTryReadVrf[1])),
    .vrfReadDataPorts_1_valid                               (_storeUnit_vrfReadDataPorts_1_valid),
    .vrfReadDataPorts_1_bits_vs                             (_storeUnit_vrfReadDataPorts_1_bits_vs),
    .vrfReadDataPorts_1_bits_offset                         (_storeUnit_vrfReadDataPorts_1_bits_offset),
    .vrfReadDataPorts_1_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_1_bits_instructionIndex),
    .vrfReadDataPorts_2_ready                               (vrfReadDataPorts_2_ready_0 & ~(otherTryReadVrf[2])),
    .vrfReadDataPorts_2_valid                               (_storeUnit_vrfReadDataPorts_2_valid),
    .vrfReadDataPorts_2_bits_vs                             (_storeUnit_vrfReadDataPorts_2_bits_vs),
    .vrfReadDataPorts_2_bits_offset                         (_storeUnit_vrfReadDataPorts_2_bits_offset),
    .vrfReadDataPorts_2_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_2_bits_instructionIndex),
    .vrfReadDataPorts_3_ready                               (vrfReadDataPorts_3_ready_0 & ~(otherTryReadVrf[3])),
    .vrfReadDataPorts_3_valid                               (_storeUnit_vrfReadDataPorts_3_valid),
    .vrfReadDataPorts_3_bits_vs                             (_storeUnit_vrfReadDataPorts_3_bits_vs),
    .vrfReadDataPorts_3_bits_offset                         (_storeUnit_vrfReadDataPorts_3_bits_offset),
    .vrfReadDataPorts_3_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_3_bits_instructionIndex),
    .vrfReadResults_0_valid                                 (vrfReadResults_0_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_0_bits                                  (vrfReadResults_0_bits),
    .vrfReadResults_1_valid                                 (vrfReadResults_1_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_1_bits                                  (vrfReadResults_1_bits),
    .vrfReadResults_2_valid                                 (vrfReadResults_2_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_2_bits                                  (vrfReadResults_2_bits),
    .vrfReadResults_3_valid                                 (vrfReadResults_3_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_3_bits                                  (vrfReadResults_3_bits),
    .storeResponse                                          (axi4Port_b_valid_0)
  );
  SimpleAccessUnit otherUnit (
    .clock                                                  (clock),
    .reset                                                  (reset),
    .lsuRequest_valid                                       (reqEnq_2),
    .lsuRequest_bits_instructionInformation_nf              (request_bits_instructionInformation_nf_0),
    .lsuRequest_bits_instructionInformation_mew             (request_bits_instructionInformation_mew_0),
    .lsuRequest_bits_instructionInformation_mop             (request_bits_instructionInformation_mop_0),
    .lsuRequest_bits_instructionInformation_lumop           (request_bits_instructionInformation_lumop_0),
    .lsuRequest_bits_instructionInformation_eew             (request_bits_instructionInformation_eew_0),
    .lsuRequest_bits_instructionInformation_vs3             (request_bits_instructionInformation_vs3_0),
    .lsuRequest_bits_instructionInformation_isStore         (request_bits_instructionInformation_isStore_0),
    .lsuRequest_bits_instructionInformation_maskedLoadStore (request_bits_instructionInformation_maskedLoadStore_0),
    .lsuRequest_bits_rs1Data                                (request_bits_rs1Data_0),
    .lsuRequest_bits_rs2Data                                (request_bits_rs2Data_0),
    .lsuRequest_bits_instructionIndex                       (request_bits_instructionIndex_0),
    .vrfReadDataPorts_ready                                 (otherUnit_vrfReadDataPorts_ready),
    .vrfReadDataPorts_valid                                 (_otherUnit_vrfReadDataPorts_valid),
    .vrfReadDataPorts_bits_vs                               (_otherUnit_vrfReadDataPorts_bits_vs),
    .vrfReadDataPorts_bits_offset                           (_otherUnit_vrfReadDataPorts_bits_offset),
    .vrfReadDataPorts_bits_instructionIndex                 (_otherUnit_vrfReadDataPorts_bits_instructionIndex),
    .vrfReadResults_valid                                   (otherUnitTargetQueue_deq_ready),
    .vrfReadResults_bits
      ((otherUnitTargetQueue_deq_bits[0] ? otherUnitDataQueueVec_0_deq_bits : 32'h0) | (otherUnitTargetQueue_deq_bits[1] ? otherUnitDataQueueVec_1_deq_bits : 32'h0)
       | (otherUnitTargetQueue_deq_bits[2] ? otherUnitDataQueueVec_2_deq_bits : 32'h0) | (otherUnitTargetQueue_deq_bits[3] ? otherUnitDataQueueVec_3_deq_bits : 32'h0)),
    .offsetReadResult_0_valid                               (offsetReadResult_0_valid),
    .offsetReadResult_0_bits                                (offsetReadResult_0_bits),
    .offsetReadResult_1_valid                               (offsetReadResult_1_valid),
    .offsetReadResult_1_bits                                (offsetReadResult_1_bits),
    .offsetReadResult_2_valid                               (offsetReadResult_2_valid),
    .offsetReadResult_2_bits                                (offsetReadResult_2_bits),
    .offsetReadResult_3_valid                               (offsetReadResult_3_valid),
    .offsetReadResult_3_bits                                (offsetReadResult_3_bits),
    .maskInput                                              (_GEN_1025[maskSelect_2]),
    .maskSelect_valid                                       (_otherUnit_maskSelect_valid),
    .maskSelect_bits                                        (_otherUnit_maskSelect_bits),
    .memReadRequest_ready                                   (simpleSourceQueue_enq_ready & simpleAccessPorts_ar_ready_0),
    .memReadRequest_valid                                   (_otherUnit_memReadRequest_valid),
    .memReadRequest_bits_address                            (simpleAccessPorts_ar_bits_addr_0),
    .memReadRequest_bits_source                             (simpleSourceQueue_enq_bits),
    .memReadResponse_ready                                  (simpleAccessPorts_r_ready_0),
    .memReadResponse_valid                                  (simpleAccessPorts_r_valid_0),
    .memReadResponse_bits_data                              (simpleAccessPorts_r_bits_data_0),
    .memReadResponse_bits_source                            (simpleSourceQueue_deq_bits),
    .memWriteRequest_ready                                  (simpleAccessPorts_aw_ready_0 & simpleDataQueue_enq_ready),
    .memWriteRequest_valid                                  (_otherUnit_memWriteRequest_valid),
    .memWriteRequest_bits_data                              (simpleDataQueue_enq_bits_data),
    .memWriteRequest_bits_mask                              (simpleDataQueue_enq_bits_mask),
    .memWriteRequest_bits_source                            (_otherUnit_memWriteRequest_bits_source),
    .memWriteRequest_bits_address                           (_otherUnit_memWriteRequest_bits_address),
    .memWriteRequest_bits_size                              (_otherUnit_memWriteRequest_bits_size),
    .vrfWritePort_ready                                     (|(_otherUnit_status_targetLane & {otherUnit_vrfWritePort_ready_hi, otherUnit_vrfWritePort_ready_lo})),
    .vrfWritePort_valid                                     (_otherUnit_vrfWritePort_valid),
    .vrfWritePort_bits_vd                                   (_otherUnit_vrfWritePort_bits_vd),
    .vrfWritePort_bits_offset                               (_otherUnit_vrfWritePort_bits_offset),
    .vrfWritePort_bits_mask                                 (_otherUnit_vrfWritePort_bits_mask),
    .vrfWritePort_bits_data                                 (_otherUnit_vrfWritePort_bits_data),
    .vrfWritePort_bits_last                                 (_otherUnit_vrfWritePort_bits_last),
    .vrfWritePort_bits_instructionIndex                     (_otherUnit_vrfWritePort_bits_instructionIndex),
    .csrInterface_vl                                        (csrInterface_vl),
    .csrInterface_vStart                                    (csrInterface_vStart),
    .csrInterface_vlmul                                     (csrInterface_vlmul),
    .csrInterface_vSew                                      (csrInterface_vSew),
    .csrInterface_vxrm                                      (csrInterface_vxrm),
    .csrInterface_vta                                       (csrInterface_vta),
    .csrInterface_vma                                       (csrInterface_vma),
    .status_idle                                            (_otherUnit_status_idle),
    .status_last                                            (_otherUnit_status_last),
    .status_instructionIndex                                (_otherUnit_status_instructionIndex),
    .status_targetLane                                      (_otherUnit_status_targetLane),
    .status_isStore                                         (_otherUnit_status_isStore),
    .offsetRelease_0                                        (_otherUnit_offsetRelease_0),
    .offsetRelease_1                                        (_otherUnit_offsetRelease_1),
    .offsetRelease_2                                        (_otherUnit_offsetRelease_2),
    .offsetRelease_3                                        (_otherUnit_offsetRelease_3)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(58)
  ) writeQueueVec_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_0_writeValid_T & ~(_writeQueueVec_fifo_empty & writeQueueVec_0_deq_ready))),
    .pop_req_n    (~(writeQueueVec_0_deq_ready & ~_writeQueueVec_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn),
    .empty        (_writeQueueVec_fifo_empty),
    .almost_empty (writeQueueVec_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_0_almostFull),
    .full         (_writeQueueVec_fifo_full),
    .error        (_writeQueueVec_fifo_error),
    .data_out     (_writeQueueVec_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(58)
  ) writeQueueVec_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_1_writeValid_T & ~(_writeQueueVec_fifo_1_empty & writeQueueVec_1_deq_ready))),
    .pop_req_n    (~(writeQueueVec_1_deq_ready & ~_writeQueueVec_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_1),
    .empty        (_writeQueueVec_fifo_1_empty),
    .almost_empty (writeQueueVec_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_1_almostFull),
    .full         (_writeQueueVec_fifo_1_full),
    .error        (_writeQueueVec_fifo_1_error),
    .data_out     (_writeQueueVec_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(58)
  ) writeQueueVec_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_2_writeValid_T & ~(_writeQueueVec_fifo_2_empty & writeQueueVec_2_deq_ready))),
    .pop_req_n    (~(writeQueueVec_2_deq_ready & ~_writeQueueVec_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_2),
    .empty        (_writeQueueVec_fifo_2_empty),
    .almost_empty (writeQueueVec_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_2_almostFull),
    .full         (_writeQueueVec_fifo_2_full),
    .error        (_writeQueueVec_fifo_2_error),
    .data_out     (_writeQueueVec_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(58)
  ) writeQueueVec_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_3_writeValid_T & ~(_writeQueueVec_fifo_3_empty & writeQueueVec_3_deq_ready))),
    .pop_req_n    (~(writeQueueVec_3_deq_ready & ~_writeQueueVec_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_3),
    .empty        (_writeQueueVec_fifo_3_empty),
    .almost_empty (writeQueueVec_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_3_almostFull),
    .full         (_writeQueueVec_fifo_3_full),
    .error        (_writeQueueVec_fifo_3_error),
    .data_out     (_writeQueueVec_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(4)
  ) otherUnitTargetQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitTargetQueue_enq_ready & otherUnitTargetQueue_enq_valid)),
    .pop_req_n    (~(otherUnitTargetQueue_deq_ready & ~_otherUnitTargetQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitTargetQueue_enq_bits),
    .empty        (_otherUnitTargetQueue_fifo_empty),
    .almost_empty (otherUnitTargetQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitTargetQueue_almostFull),
    .full         (_otherUnitTargetQueue_fifo_full),
    .error        (_otherUnitTargetQueue_fifo_error),
    .data_out     (otherUnitTargetQueue_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_0_enq_ready & otherUnitDataQueueVec_0_enq_valid & ~(_otherUnitDataQueueVec_fifo_empty & otherUnitDataQueueVec_0_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_0_deq_ready & ~_otherUnitDataQueueVec_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_0_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_empty),
    .almost_empty (otherUnitDataQueueVec_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_0_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_full),
    .error        (_otherUnitDataQueueVec_fifo_error),
    .data_out     (_otherUnitDataQueueVec_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_1_enq_ready & otherUnitDataQueueVec_1_enq_valid & ~(_otherUnitDataQueueVec_fifo_1_empty & otherUnitDataQueueVec_1_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_1_deq_ready & ~_otherUnitDataQueueVec_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_1_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_1_empty),
    .almost_empty (otherUnitDataQueueVec_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_1_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_1_full),
    .error        (_otherUnitDataQueueVec_fifo_1_error),
    .data_out     (_otherUnitDataQueueVec_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_2_enq_ready & otherUnitDataQueueVec_2_enq_valid & ~(_otherUnitDataQueueVec_fifo_2_empty & otherUnitDataQueueVec_2_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_2_deq_ready & ~_otherUnitDataQueueVec_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_2_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_2_empty),
    .almost_empty (otherUnitDataQueueVec_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_2_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_2_full),
    .error        (_otherUnitDataQueueVec_fifo_2_error),
    .data_out     (_otherUnitDataQueueVec_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_3_enq_ready & otherUnitDataQueueVec_3_enq_valid & ~(_otherUnitDataQueueVec_fifo_3_empty & otherUnitDataQueueVec_3_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_3_deq_ready & ~_otherUnitDataQueueVec_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_3_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_3_empty),
    .almost_empty (otherUnitDataQueueVec_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_3_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_3_full),
    .error        (_otherUnitDataQueueVec_fifo_3_error),
    .data_out     (_otherUnitDataQueueVec_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_enq_ready & writeIndexQueue_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_deq_ready & ~_writeIndexQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_enq_bits),
    .empty        (_writeIndexQueue_fifo_empty),
    .almost_empty (writeIndexQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_almostFull),
    .full         (_writeIndexQueue_fifo_full),
    .error        (_writeIndexQueue_fifo_error),
    .data_out     (writeIndexQueue_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_1_enq_ready & writeIndexQueue_1_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_1_deq_ready & ~_writeIndexQueue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_1_enq_bits),
    .empty        (_writeIndexQueue_fifo_1_empty),
    .almost_empty (writeIndexQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_1_almostFull),
    .full         (_writeIndexQueue_fifo_1_full),
    .error        (_writeIndexQueue_fifo_1_error),
    .data_out     (writeIndexQueue_1_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_2_enq_ready & writeIndexQueue_2_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_2_deq_ready & ~_writeIndexQueue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_2_enq_bits),
    .empty        (_writeIndexQueue_fifo_2_empty),
    .almost_empty (writeIndexQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_2_almostFull),
    .full         (_writeIndexQueue_fifo_2_full),
    .error        (_writeIndexQueue_fifo_2_error),
    .data_out     (writeIndexQueue_2_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_3_enq_ready & writeIndexQueue_3_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_3_deq_ready & ~_writeIndexQueue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_3_enq_bits),
    .empty        (_writeIndexQueue_fifo_3_empty),
    .almost_empty (writeIndexQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_3_almostFull),
    .full         (_writeIndexQueue_fifo_3_full),
    .error        (_writeIndexQueue_fifo_3_error),
    .data_out     (writeIndexQueue_3_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(32),
    .err_mode(2),
    .rst_mode(3),
    .width(13)
  ) sourceQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sourceQueue_enq_ready & sourceQueue_enq_valid)),
    .pop_req_n    (~(sourceQueue_deq_ready & ~_sourceQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (sourceQueue_enq_bits),
    .empty        (_sourceQueue_fifo_empty),
    .almost_empty (sourceQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sourceQueue_almostFull),
    .full         (_sourceQueue_fifo_full),
    .error        (_sourceQueue_fifo_error),
    .data_out     (sourceQueue_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(2),
    .err_mode(2),
    .rst_mode(3),
    .width(189)
  ) dataQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(dataQueue_enq_ready & dataQueue_enq_valid)),
    .pop_req_n    (~(dataQueue_deq_ready & ~_dataQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (dataQueue_dataIn),
    .empty        (_dataQueue_fifo_empty),
    .almost_empty (dataQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (dataQueue_almostFull),
    .full         (_dataQueue_fifo_full),
    .error        (_dataQueue_fifo_error),
    .data_out     (_dataQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(32),
    .err_mode(2),
    .rst_mode(3),
    .width(7)
  ) simpleSourceQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(simpleSourceQueue_enq_ready & simpleSourceQueue_enq_valid)),
    .pop_req_n    (~(simpleSourceQueue_deq_ready & ~_simpleSourceQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (simpleSourceQueue_enq_bits),
    .empty        (_simpleSourceQueue_fifo_empty),
    .almost_empty (simpleSourceQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (simpleSourceQueue_almostFull),
    .full         (_simpleSourceQueue_fifo_full),
    .error        (_simpleSourceQueue_fifo_error),
    .data_out     (simpleSourceQueue_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(2),
    .err_mode(2),
    .rst_mode(3),
    .width(78)
  ) simpleDataQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(simpleDataQueue_enq_ready & simpleDataQueue_enq_valid)),
    .pop_req_n    (~(simpleDataQueue_deq_ready & ~_simpleDataQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (simpleDataQueue_dataIn),
    .empty        (_simpleDataQueue_fifo_empty),
    .almost_empty (simpleDataQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (simpleDataQueue_almostFull),
    .full         (_simpleDataQueue_fifo_full),
    .error        (_simpleDataQueue_fifo_error),
    .data_out     (_simpleDataQueue_fifo_data_out)
  );
  assign request_ready = request_ready_0;
  assign axi4Port_aw_valid = axi4Port_aw_valid_0;
  assign axi4Port_aw_bits_id = axi4Port_aw_bits_id_0;
  assign axi4Port_aw_bits_addr = axi4Port_aw_bits_addr_0;
  assign axi4Port_w_valid = axi4Port_w_valid_0;
  assign axi4Port_w_bits_data = axi4Port_w_bits_data_0;
  assign axi4Port_w_bits_strb = axi4Port_w_bits_strb_0;
  assign axi4Port_ar_valid = axi4Port_ar_valid_0;
  assign axi4Port_ar_bits_addr = axi4Port_ar_bits_addr_0;
  assign axi4Port_r_ready = axi4Port_r_ready_0;
  assign simpleAccessPorts_aw_valid = simpleAccessPorts_aw_valid_0;
  assign simpleAccessPorts_aw_bits_id = simpleAccessPorts_aw_bits_id_0;
  assign simpleAccessPorts_aw_bits_addr = simpleAccessPorts_aw_bits_addr_0;
  assign simpleAccessPorts_aw_bits_size = simpleAccessPorts_aw_bits_size_0;
  assign simpleAccessPorts_w_valid = simpleAccessPorts_w_valid_0;
  assign simpleAccessPorts_w_bits_data = simpleAccessPorts_w_bits_data_0;
  assign simpleAccessPorts_w_bits_strb = simpleAccessPorts_w_bits_strb_0;
  assign simpleAccessPorts_ar_valid = simpleAccessPorts_ar_valid_0;
  assign simpleAccessPorts_ar_bits_addr = simpleAccessPorts_ar_bits_addr_0;
  assign simpleAccessPorts_r_ready = simpleAccessPorts_r_ready_0;
  assign vrfReadDataPorts_0_valid = vrfReadDataPorts_0_valid_0;
  assign vrfReadDataPorts_0_bits_vs = vrfReadDataPorts_0_bits_vs_0;
  assign vrfReadDataPorts_0_bits_offset = vrfReadDataPorts_0_bits_offset_0;
  assign vrfReadDataPorts_0_bits_instructionIndex = vrfReadDataPorts_0_bits_instructionIndex_0;
  assign vrfReadDataPorts_1_valid = vrfReadDataPorts_1_valid_0;
  assign vrfReadDataPorts_1_bits_vs = vrfReadDataPorts_1_bits_vs_0;
  assign vrfReadDataPorts_1_bits_offset = vrfReadDataPorts_1_bits_offset_0;
  assign vrfReadDataPorts_1_bits_instructionIndex = vrfReadDataPorts_1_bits_instructionIndex_0;
  assign vrfReadDataPorts_2_valid = vrfReadDataPorts_2_valid_0;
  assign vrfReadDataPorts_2_bits_vs = vrfReadDataPorts_2_bits_vs_0;
  assign vrfReadDataPorts_2_bits_offset = vrfReadDataPorts_2_bits_offset_0;
  assign vrfReadDataPorts_2_bits_instructionIndex = vrfReadDataPorts_2_bits_instructionIndex_0;
  assign vrfReadDataPorts_3_valid = vrfReadDataPorts_3_valid_0;
  assign vrfReadDataPorts_3_bits_vs = vrfReadDataPorts_3_bits_vs_0;
  assign vrfReadDataPorts_3_bits_offset = vrfReadDataPorts_3_bits_offset_0;
  assign vrfReadDataPorts_3_bits_instructionIndex = vrfReadDataPorts_3_bits_instructionIndex_0;
  assign vrfWritePort_0_valid = vrfWritePort_0_valid_0;
  assign vrfWritePort_0_bits_vd = vrfWritePort_0_bits_vd_0;
  assign vrfWritePort_0_bits_offset = vrfWritePort_0_bits_offset_0;
  assign vrfWritePort_0_bits_mask = vrfWritePort_0_bits_mask_0;
  assign vrfWritePort_0_bits_data = vrfWritePort_0_bits_data_0;
  assign vrfWritePort_0_bits_last = vrfWritePort_0_bits_last_0;
  assign vrfWritePort_0_bits_instructionIndex = vrfWritePort_0_bits_instructionIndex_0;
  assign vrfWritePort_1_valid = vrfWritePort_1_valid_0;
  assign vrfWritePort_1_bits_vd = vrfWritePort_1_bits_vd_0;
  assign vrfWritePort_1_bits_offset = vrfWritePort_1_bits_offset_0;
  assign vrfWritePort_1_bits_mask = vrfWritePort_1_bits_mask_0;
  assign vrfWritePort_1_bits_data = vrfWritePort_1_bits_data_0;
  assign vrfWritePort_1_bits_last = vrfWritePort_1_bits_last_0;
  assign vrfWritePort_1_bits_instructionIndex = vrfWritePort_1_bits_instructionIndex_0;
  assign vrfWritePort_2_valid = vrfWritePort_2_valid_0;
  assign vrfWritePort_2_bits_vd = vrfWritePort_2_bits_vd_0;
  assign vrfWritePort_2_bits_offset = vrfWritePort_2_bits_offset_0;
  assign vrfWritePort_2_bits_mask = vrfWritePort_2_bits_mask_0;
  assign vrfWritePort_2_bits_data = vrfWritePort_2_bits_data_0;
  assign vrfWritePort_2_bits_last = vrfWritePort_2_bits_last_0;
  assign vrfWritePort_2_bits_instructionIndex = vrfWritePort_2_bits_instructionIndex_0;
  assign vrfWritePort_3_valid = vrfWritePort_3_valid_0;
  assign vrfWritePort_3_bits_vd = vrfWritePort_3_bits_vd_0;
  assign vrfWritePort_3_bits_offset = vrfWritePort_3_bits_offset_0;
  assign vrfWritePort_3_bits_mask = vrfWritePort_3_bits_mask_0;
  assign vrfWritePort_3_bits_data = vrfWritePort_3_bits_data_0;
  assign vrfWritePort_3_bits_last = vrfWritePort_3_bits_last_0;
  assign vrfWritePort_3_bits_instructionIndex = vrfWritePort_3_bits_instructionIndex_0;
  assign dataInWriteQueue_0 = {dataInWriteQueue_0_hi, dataInWriteQueue_0_lo} | dataInMSHR;
  assign dataInWriteQueue_1 = {dataInWriteQueue_1_hi, dataInWriteQueue_1_lo} | dataInMSHR;
  assign dataInWriteQueue_2 = {dataInWriteQueue_2_hi, dataInWriteQueue_2_lo} | dataInMSHR;
  assign dataInWriteQueue_3 = {dataInWriteQueue_3_hi, dataInWriteQueue_3_lo} | dataInMSHR;
  assign lastReport = (_loadUnit_status_last ? 8'h1 << _GEN_1026 : 8'h0) | (_storeUnit_status_last ? 8'h1 << _storeUnit_status_instructionIndex : 8'h0) | (_otherUnit_status_last ? 8'h1 << _GEN_1027 : 8'h0);
  assign tokenIO_offsetGroupRelease = {tokenIO_offsetGroupRelease_hi, tokenIO_offsetGroupRelease_lo};
endmodule

