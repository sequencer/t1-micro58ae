
// Include register initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for register randomization.

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_
module MaskCompress(
  input          clock,
                 reset,
                 in_valid,
                 in_bits_maskType,
  input  [1:0]   in_bits_eew,
  input  [2:0]   in_bits_uop,
  input  [31:0]  in_bits_readFromScalar,
                 in_bits_source1,
                 in_bits_mask,
  input  [511:0] in_bits_source2,
                 in_bits_pipeData,
  input  [5:0]   in_bits_groupCounter,
  input  [15:0]  in_bits_ffoInput,
                 in_bits_validInput,
  input          in_bits_lastCompress,
  output [511:0] out_data,
  output [63:0]  out_mask,
  output [5:0]   out_groupCounter,
  output [15:0]  out_ffoOutput,
  output         out_compressValid,
  input          newInstruction,
                 ffoInstruction,
  output [31:0]  writeData,
  output         stageValid
);

  wire          compressDataVec_useTail_63 = 1'h0;
  wire          compressTailMask_elementValid_63 = 1'h0;
  reg           in_1_valid;
  reg           in_1_bits_maskType;
  reg  [1:0]    in_1_bits_eew;
  reg  [2:0]    in_1_bits_uop;
  reg  [31:0]   in_1_bits_readFromScalar;
  reg  [31:0]   in_1_bits_source1;
  reg  [31:0]   in_1_bits_mask;
  reg  [511:0]  in_1_bits_source2;
  reg  [511:0]  in_1_bits_pipeData;
  reg  [5:0]    in_1_bits_groupCounter;
  reg  [15:0]   in_1_bits_ffoInput;
  reg  [15:0]   in_1_bits_validInput;
  reg           in_1_bits_lastCompress;
  wire          compress = in_1_bits_uop == 3'h1;
  wire          viota = in_1_bits_uop == 3'h0;
  wire          mv = in_1_bits_uop == 3'h2;
  wire          mvRd = in_1_bits_uop == 3'h3;
  wire          writeRD = &(in_1_bits_uop[1:0]);
  wire          ffoType = &(in_1_bits_uop[2:1]);
  wire [3:0]    _eew1H_T = 4'h1 << in_1_bits_eew;
  wire [2:0]    eew1H = _eew1H_T[2:0];
  reg  [10:0]   compressInit;
  wire [10:0]   compressVec_0 = compressInit;
  wire [63:0]   maskInput = {32'h0, in_1_bits_source1 & in_1_bits_mask};
  wire          compressMaskVec_0 = maskInput[0];
  wire          compressMaskVec_1 = maskInput[1];
  wire          compressMaskVec_2 = maskInput[2];
  wire          compressMaskVec_3 = maskInput[3];
  wire          compressMaskVec_4 = maskInput[4];
  wire          compressMaskVec_5 = maskInput[5];
  wire          compressMaskVec_6 = maskInput[6];
  wire          compressMaskVec_7 = maskInput[7];
  wire          compressMaskVec_8 = maskInput[8];
  wire          compressMaskVec_9 = maskInput[9];
  wire          compressMaskVec_10 = maskInput[10];
  wire          compressMaskVec_11 = maskInput[11];
  wire          compressMaskVec_12 = maskInput[12];
  wire          compressMaskVec_13 = maskInput[13];
  wire          compressMaskVec_14 = maskInput[14];
  wire          compressMaskVec_15 = maskInput[15];
  wire          compressMaskVec_16 = maskInput[16];
  wire          compressMaskVec_17 = maskInput[17];
  wire          compressMaskVec_18 = maskInput[18];
  wire          compressMaskVec_19 = maskInput[19];
  wire          compressMaskVec_20 = maskInput[20];
  wire          compressMaskVec_21 = maskInput[21];
  wire          compressMaskVec_22 = maskInput[22];
  wire          compressMaskVec_23 = maskInput[23];
  wire          compressMaskVec_24 = maskInput[24];
  wire          compressMaskVec_25 = maskInput[25];
  wire          compressMaskVec_26 = maskInput[26];
  wire          compressMaskVec_27 = maskInput[27];
  wire          compressMaskVec_28 = maskInput[28];
  wire          compressMaskVec_29 = maskInput[29];
  wire          compressMaskVec_30 = maskInput[30];
  wire          compressMaskVec_31 = maskInput[31];
  wire          compressMaskVec_32 = maskInput[32];
  wire          compressMaskVec_33 = maskInput[33];
  wire          compressMaskVec_34 = maskInput[34];
  wire          compressMaskVec_35 = maskInput[35];
  wire          compressMaskVec_36 = maskInput[36];
  wire          compressMaskVec_37 = maskInput[37];
  wire          compressMaskVec_38 = maskInput[38];
  wire          compressMaskVec_39 = maskInput[39];
  wire          compressMaskVec_40 = maskInput[40];
  wire          compressMaskVec_41 = maskInput[41];
  wire          compressMaskVec_42 = maskInput[42];
  wire          compressMaskVec_43 = maskInput[43];
  wire          compressMaskVec_44 = maskInput[44];
  wire          compressMaskVec_45 = maskInput[45];
  wire          compressMaskVec_46 = maskInput[46];
  wire          compressMaskVec_47 = maskInput[47];
  wire          compressMaskVec_48 = maskInput[48];
  wire          compressMaskVec_49 = maskInput[49];
  wire          compressMaskVec_50 = maskInput[50];
  wire          compressMaskVec_51 = maskInput[51];
  wire          compressMaskVec_52 = maskInput[52];
  wire          compressMaskVec_53 = maskInput[53];
  wire          compressMaskVec_54 = maskInput[54];
  wire          compressMaskVec_55 = maskInput[55];
  wire          compressMaskVec_56 = maskInput[56];
  wire          compressMaskVec_57 = maskInput[57];
  wire          compressMaskVec_58 = maskInput[58];
  wire          compressMaskVec_59 = maskInput[59];
  wire          compressMaskVec_60 = maskInput[60];
  wire          compressMaskVec_61 = maskInput[61];
  wire          compressMaskVec_62 = maskInput[62];
  wire          compressMaskVec_63 = maskInput[63];
  wire [10:0]   compressCount =
    compressInit
    + {4'h0,
       {1'h0,
        {1'h0,
         {1'h0,
          {1'h0, {1'h0, {1'h0, compressMaskVec_0} + {1'h0, compressMaskVec_1}} + {1'h0, {1'h0, compressMaskVec_2} + {1'h0, compressMaskVec_3}}}
            + {1'h0, {1'h0, {1'h0, compressMaskVec_4} + {1'h0, compressMaskVec_5}} + {1'h0, {1'h0, compressMaskVec_6} + {1'h0, compressMaskVec_7}}}}
           + {1'h0,
              {1'h0, {1'h0, {1'h0, compressMaskVec_8} + {1'h0, compressMaskVec_9}} + {1'h0, {1'h0, compressMaskVec_10} + {1'h0, compressMaskVec_11}}}
                + {1'h0, {1'h0, {1'h0, compressMaskVec_12} + {1'h0, compressMaskVec_13}} + {1'h0, {1'h0, compressMaskVec_14} + {1'h0, compressMaskVec_15}}}}}
          + {1'h0,
             {1'h0,
              {1'h0, {1'h0, {1'h0, compressMaskVec_16} + {1'h0, compressMaskVec_17}} + {1'h0, {1'h0, compressMaskVec_18} + {1'h0, compressMaskVec_19}}}
                + {1'h0, {1'h0, {1'h0, compressMaskVec_20} + {1'h0, compressMaskVec_21}} + {1'h0, {1'h0, compressMaskVec_22} + {1'h0, compressMaskVec_23}}}}
               + {1'h0,
                  {1'h0, {1'h0, {1'h0, compressMaskVec_24} + {1'h0, compressMaskVec_25}} + {1'h0, {1'h0, compressMaskVec_26} + {1'h0, compressMaskVec_27}}}
                    + {1'h0, {1'h0, {1'h0, compressMaskVec_28} + {1'h0, compressMaskVec_29}} + {1'h0, {1'h0, compressMaskVec_30} + {1'h0, compressMaskVec_31}}}}}}
         + {1'h0,
            {1'h0,
             {1'h0,
              {1'h0, {1'h0, {1'h0, compressMaskVec_32} + {1'h0, compressMaskVec_33}} + {1'h0, {1'h0, compressMaskVec_34} + {1'h0, compressMaskVec_35}}}
                + {1'h0, {1'h0, {1'h0, compressMaskVec_36} + {1'h0, compressMaskVec_37}} + {1'h0, {1'h0, compressMaskVec_38} + {1'h0, compressMaskVec_39}}}}
               + {1'h0,
                  {1'h0, {1'h0, {1'h0, compressMaskVec_40} + {1'h0, compressMaskVec_41}} + {1'h0, {1'h0, compressMaskVec_42} + {1'h0, compressMaskVec_43}}}
                    + {1'h0, {1'h0, {1'h0, compressMaskVec_44} + {1'h0, compressMaskVec_45}} + {1'h0, {1'h0, compressMaskVec_46} + {1'h0, compressMaskVec_47}}}}}
              + {1'h0,
                 {1'h0,
                  {1'h0, {1'h0, {1'h0, compressMaskVec_48} + {1'h0, compressMaskVec_49}} + {1'h0, {1'h0, compressMaskVec_50} + {1'h0, compressMaskVec_51}}}
                    + {1'h0, {1'h0, {1'h0, compressMaskVec_52} + {1'h0, compressMaskVec_53}} + {1'h0, {1'h0, compressMaskVec_54} + {1'h0, compressMaskVec_55}}}}
                   + {1'h0,
                      {1'h0, {1'h0, {1'h0, compressMaskVec_56} + {1'h0, compressMaskVec_57}} + {1'h0, {1'h0, compressMaskVec_58} + {1'h0, compressMaskVec_59}}}
                        + {1'h0, {1'h0, {1'h0, compressMaskVec_60} + {1'h0, compressMaskVec_61}} + {1'h0, {1'h0, compressMaskVec_62} + {1'h0, compressMaskVec_63}}}}}}};
  wire [10:0]   compressVec_1 = compressInit + {10'h0, compressMaskVec_0};
  wire [10:0]   compressVec_2 = compressVec_1 + {10'h0, compressMaskVec_1};
  wire [10:0]   compressVec_3 = compressVec_2 + {10'h0, compressMaskVec_2};
  wire [10:0]   compressVec_4 = compressVec_3 + {10'h0, compressMaskVec_3};
  wire [10:0]   compressVec_5 = compressVec_4 + {10'h0, compressMaskVec_4};
  wire [10:0]   compressVec_6 = compressVec_5 + {10'h0, compressMaskVec_5};
  wire [10:0]   compressVec_7 = compressVec_6 + {10'h0, compressMaskVec_6};
  wire [10:0]   compressVec_8 = compressVec_7 + {10'h0, compressMaskVec_7};
  wire [10:0]   compressVec_9 = compressVec_8 + {10'h0, compressMaskVec_8};
  wire [10:0]   compressVec_10 = compressVec_9 + {10'h0, compressMaskVec_9};
  wire [10:0]   compressVec_11 = compressVec_10 + {10'h0, compressMaskVec_10};
  wire [10:0]   compressVec_12 = compressVec_11 + {10'h0, compressMaskVec_11};
  wire [10:0]   compressVec_13 = compressVec_12 + {10'h0, compressMaskVec_12};
  wire [10:0]   compressVec_14 = compressVec_13 + {10'h0, compressMaskVec_13};
  wire [10:0]   compressVec_15 = compressVec_14 + {10'h0, compressMaskVec_14};
  wire [10:0]   compressVec_16 = compressVec_15 + {10'h0, compressMaskVec_15};
  wire [10:0]   compressVec_17 = compressVec_16 + {10'h0, compressMaskVec_16};
  wire [10:0]   compressVec_18 = compressVec_17 + {10'h0, compressMaskVec_17};
  wire [10:0]   compressVec_19 = compressVec_18 + {10'h0, compressMaskVec_18};
  wire [10:0]   compressVec_20 = compressVec_19 + {10'h0, compressMaskVec_19};
  wire [10:0]   compressVec_21 = compressVec_20 + {10'h0, compressMaskVec_20};
  wire [10:0]   compressVec_22 = compressVec_21 + {10'h0, compressMaskVec_21};
  wire [10:0]   compressVec_23 = compressVec_22 + {10'h0, compressMaskVec_22};
  wire [10:0]   compressVec_24 = compressVec_23 + {10'h0, compressMaskVec_23};
  wire [10:0]   compressVec_25 = compressVec_24 + {10'h0, compressMaskVec_24};
  wire [10:0]   compressVec_26 = compressVec_25 + {10'h0, compressMaskVec_25};
  wire [10:0]   compressVec_27 = compressVec_26 + {10'h0, compressMaskVec_26};
  wire [10:0]   compressVec_28 = compressVec_27 + {10'h0, compressMaskVec_27};
  wire [10:0]   compressVec_29 = compressVec_28 + {10'h0, compressMaskVec_28};
  wire [10:0]   compressVec_30 = compressVec_29 + {10'h0, compressMaskVec_29};
  wire [10:0]   compressVec_31 = compressVec_30 + {10'h0, compressMaskVec_30};
  wire [10:0]   compressVec_32 = compressVec_31 + {10'h0, compressMaskVec_31};
  wire [10:0]   compressVec_33 = compressVec_32 + {10'h0, compressMaskVec_32};
  wire [10:0]   compressVec_34 = compressVec_33 + {10'h0, compressMaskVec_33};
  wire [10:0]   compressVec_35 = compressVec_34 + {10'h0, compressMaskVec_34};
  wire [10:0]   compressVec_36 = compressVec_35 + {10'h0, compressMaskVec_35};
  wire [10:0]   compressVec_37 = compressVec_36 + {10'h0, compressMaskVec_36};
  wire [10:0]   compressVec_38 = compressVec_37 + {10'h0, compressMaskVec_37};
  wire [10:0]   compressVec_39 = compressVec_38 + {10'h0, compressMaskVec_38};
  wire [10:0]   compressVec_40 = compressVec_39 + {10'h0, compressMaskVec_39};
  wire [10:0]   compressVec_41 = compressVec_40 + {10'h0, compressMaskVec_40};
  wire [10:0]   compressVec_42 = compressVec_41 + {10'h0, compressMaskVec_41};
  wire [10:0]   compressVec_43 = compressVec_42 + {10'h0, compressMaskVec_42};
  wire [10:0]   compressVec_44 = compressVec_43 + {10'h0, compressMaskVec_43};
  wire [10:0]   compressVec_45 = compressVec_44 + {10'h0, compressMaskVec_44};
  wire [10:0]   compressVec_46 = compressVec_45 + {10'h0, compressMaskVec_45};
  wire [10:0]   compressVec_47 = compressVec_46 + {10'h0, compressMaskVec_46};
  wire [10:0]   compressVec_48 = compressVec_47 + {10'h0, compressMaskVec_47};
  wire [10:0]   compressVec_49 = compressVec_48 + {10'h0, compressMaskVec_48};
  wire [10:0]   compressVec_50 = compressVec_49 + {10'h0, compressMaskVec_49};
  wire [10:0]   compressVec_51 = compressVec_50 + {10'h0, compressMaskVec_50};
  wire [10:0]   compressVec_52 = compressVec_51 + {10'h0, compressMaskVec_51};
  wire [10:0]   compressVec_53 = compressVec_52 + {10'h0, compressMaskVec_52};
  wire [10:0]   compressVec_54 = compressVec_53 + {10'h0, compressMaskVec_53};
  wire [10:0]   compressVec_55 = compressVec_54 + {10'h0, compressMaskVec_54};
  wire [10:0]   compressVec_56 = compressVec_55 + {10'h0, compressMaskVec_55};
  wire [10:0]   compressVec_57 = compressVec_56 + {10'h0, compressMaskVec_56};
  wire [10:0]   compressVec_58 = compressVec_57 + {10'h0, compressMaskVec_57};
  wire [10:0]   compressVec_59 = compressVec_58 + {10'h0, compressMaskVec_58};
  wire [10:0]   compressVec_60 = compressVec_59 + {10'h0, compressMaskVec_59};
  wire [10:0]   compressVec_61 = compressVec_60 + {10'h0, compressMaskVec_60};
  wire [10:0]   compressVec_62 = compressVec_61 + {10'h0, compressMaskVec_61};
  wire [10:0]   compressVec_63 = compressVec_62 + {10'h0, compressMaskVec_62};
  reg  [31:0]   ffoIndex;
  reg           ffoValid;
  wire          countSplit_0_1 = compressCount[6];
  wire [5:0]    countSplit_0_2 = compressCount[5:0];
  wire          countSplit_1_1 = compressCount[5];
  wire [4:0]    countSplit_1_2 = compressCount[4:0];
  wire          countSplit_2_1 = compressCount[4];
  wire [3:0]    countSplit_2_2 = compressCount[3:0];
  wire          compressDeqValid = eew1H[0] & countSplit_0_1 | eew1H[1] & countSplit_1_1 | eew1H[2] & countSplit_2_1 | ~compress;
  wire [5:0]    _compressCountSelect_T_3 = eew1H[0] ? countSplit_0_2 : 6'h0;
  wire [4:0]    _GEN = _compressCountSelect_T_3[4:0] | (eew1H[1] ? countSplit_1_2 : 5'h0);
  wire [5:0]    compressCountSelect = {_compressCountSelect_T_3[5], _GEN[4], _GEN[3:0] | (eew1H[2] ? countSplit_2_2 : 4'h0)};
  reg  [10:0]   compressVecPipe_0;
  reg  [10:0]   compressVecPipe_1;
  reg  [10:0]   compressVecPipe_2;
  reg  [10:0]   compressVecPipe_3;
  reg  [10:0]   compressVecPipe_4;
  reg  [10:0]   compressVecPipe_5;
  reg  [10:0]   compressVecPipe_6;
  reg  [10:0]   compressVecPipe_7;
  reg  [10:0]   compressVecPipe_8;
  reg  [10:0]   compressVecPipe_9;
  reg  [10:0]   compressVecPipe_10;
  reg  [10:0]   compressVecPipe_11;
  reg  [10:0]   compressVecPipe_12;
  reg  [10:0]   compressVecPipe_13;
  reg  [10:0]   compressVecPipe_14;
  reg  [10:0]   compressVecPipe_15;
  reg  [10:0]   compressVecPipe_16;
  reg  [10:0]   compressVecPipe_17;
  reg  [10:0]   compressVecPipe_18;
  reg  [10:0]   compressVecPipe_19;
  reg  [10:0]   compressVecPipe_20;
  reg  [10:0]   compressVecPipe_21;
  reg  [10:0]   compressVecPipe_22;
  reg  [10:0]   compressVecPipe_23;
  reg  [10:0]   compressVecPipe_24;
  reg  [10:0]   compressVecPipe_25;
  reg  [10:0]   compressVecPipe_26;
  reg  [10:0]   compressVecPipe_27;
  reg  [10:0]   compressVecPipe_28;
  reg  [10:0]   compressVecPipe_29;
  reg  [10:0]   compressVecPipe_30;
  reg  [10:0]   compressVecPipe_31;
  reg  [10:0]   compressVecPipe_32;
  reg  [10:0]   compressVecPipe_33;
  reg  [10:0]   compressVecPipe_34;
  reg  [10:0]   compressVecPipe_35;
  reg  [10:0]   compressVecPipe_36;
  reg  [10:0]   compressVecPipe_37;
  reg  [10:0]   compressVecPipe_38;
  reg  [10:0]   compressVecPipe_39;
  reg  [10:0]   compressVecPipe_40;
  reg  [10:0]   compressVecPipe_41;
  reg  [10:0]   compressVecPipe_42;
  reg  [10:0]   compressVecPipe_43;
  reg  [10:0]   compressVecPipe_44;
  reg  [10:0]   compressVecPipe_45;
  reg  [10:0]   compressVecPipe_46;
  reg  [10:0]   compressVecPipe_47;
  reg  [10:0]   compressVecPipe_48;
  reg  [10:0]   compressVecPipe_49;
  reg  [10:0]   compressVecPipe_50;
  reg  [10:0]   compressVecPipe_51;
  reg  [10:0]   compressVecPipe_52;
  reg  [10:0]   compressVecPipe_53;
  reg  [10:0]   compressVecPipe_54;
  reg  [10:0]   compressVecPipe_55;
  reg  [10:0]   compressVecPipe_56;
  reg  [10:0]   compressVecPipe_57;
  reg  [10:0]   compressVecPipe_58;
  reg  [10:0]   compressVecPipe_59;
  reg  [10:0]   compressVecPipe_60;
  reg  [10:0]   compressVecPipe_61;
  reg  [10:0]   compressVecPipe_62;
  reg  [10:0]   compressVecPipe_63;
  reg           compressMaskVecPipe_0;
  reg           compressMaskVecPipe_1;
  reg           compressMaskVecPipe_2;
  reg           compressMaskVecPipe_3;
  reg           compressMaskVecPipe_4;
  reg           compressMaskVecPipe_5;
  reg           compressMaskVecPipe_6;
  reg           compressMaskVecPipe_7;
  reg           compressMaskVecPipe_8;
  reg           compressMaskVecPipe_9;
  reg           compressMaskVecPipe_10;
  reg           compressMaskVecPipe_11;
  reg           compressMaskVecPipe_12;
  reg           compressMaskVecPipe_13;
  reg           compressMaskVecPipe_14;
  reg           compressMaskVecPipe_15;
  reg           compressMaskVecPipe_16;
  reg           compressMaskVecPipe_17;
  reg           compressMaskVecPipe_18;
  reg           compressMaskVecPipe_19;
  reg           compressMaskVecPipe_20;
  reg           compressMaskVecPipe_21;
  reg           compressMaskVecPipe_22;
  reg           compressMaskVecPipe_23;
  reg           compressMaskVecPipe_24;
  reg           compressMaskVecPipe_25;
  reg           compressMaskVecPipe_26;
  reg           compressMaskVecPipe_27;
  reg           compressMaskVecPipe_28;
  reg           compressMaskVecPipe_29;
  reg           compressMaskVecPipe_30;
  reg           compressMaskVecPipe_31;
  reg           compressMaskVecPipe_32;
  reg           compressMaskVecPipe_33;
  reg           compressMaskVecPipe_34;
  reg           compressMaskVecPipe_35;
  reg           compressMaskVecPipe_36;
  reg           compressMaskVecPipe_37;
  reg           compressMaskVecPipe_38;
  reg           compressMaskVecPipe_39;
  reg           compressMaskVecPipe_40;
  reg           compressMaskVecPipe_41;
  reg           compressMaskVecPipe_42;
  reg           compressMaskVecPipe_43;
  reg           compressMaskVecPipe_44;
  reg           compressMaskVecPipe_45;
  reg           compressMaskVecPipe_46;
  reg           compressMaskVecPipe_47;
  reg           compressMaskVecPipe_48;
  reg           compressMaskVecPipe_49;
  reg           compressMaskVecPipe_50;
  reg           compressMaskVecPipe_51;
  reg           compressMaskVecPipe_52;
  reg           compressMaskVecPipe_53;
  reg           compressMaskVecPipe_54;
  reg           compressMaskVecPipe_55;
  reg           compressMaskVecPipe_56;
  reg           compressMaskVecPipe_57;
  reg           compressMaskVecPipe_58;
  reg           compressMaskVecPipe_59;
  reg           compressMaskVecPipe_60;
  reg           compressMaskVecPipe_61;
  reg           compressMaskVecPipe_62;
  reg           compressMaskVecPipe_63;
  reg  [31:0]   maskPipe;
  reg  [511:0]  source2Pipe;
  reg           lastCompressPipe;
  reg           stage2Valid;
  reg           newInstructionPipe;
  reg  [10:0]   compressInitPipe;
  reg           compressDeqValidPipe;
  reg  [5:0]    groupCounterPipe;
  wire [7:0]    viotaResult_res_0 = compressVecPipe_0[7:0];
  wire [7:0]    viotaResult_res_1 = compressVecPipe_1[7:0];
  wire [7:0]    viotaResult_res_2 = compressVecPipe_2[7:0];
  wire [7:0]    viotaResult_res_3 = compressVecPipe_3[7:0];
  wire [15:0]   viotaResult_lo = {viotaResult_res_1, viotaResult_res_0};
  wire [15:0]   viotaResult_hi = {viotaResult_res_3, viotaResult_res_2};
  wire [7:0]    viotaResult_res_0_1 = compressVecPipe_4[7:0];
  wire [7:0]    viotaResult_res_1_1 = compressVecPipe_5[7:0];
  wire [7:0]    viotaResult_res_2_1 = compressVecPipe_6[7:0];
  wire [7:0]    viotaResult_res_3_1 = compressVecPipe_7[7:0];
  wire [15:0]   viotaResult_lo_1 = {viotaResult_res_1_1, viotaResult_res_0_1};
  wire [15:0]   viotaResult_hi_1 = {viotaResult_res_3_1, viotaResult_res_2_1};
  wire [7:0]    viotaResult_res_0_2 = compressVecPipe_8[7:0];
  wire [7:0]    viotaResult_res_1_2 = compressVecPipe_9[7:0];
  wire [7:0]    viotaResult_res_2_2 = compressVecPipe_10[7:0];
  wire [7:0]    viotaResult_res_3_2 = compressVecPipe_11[7:0];
  wire [15:0]   viotaResult_lo_2 = {viotaResult_res_1_2, viotaResult_res_0_2};
  wire [15:0]   viotaResult_hi_2 = {viotaResult_res_3_2, viotaResult_res_2_2};
  wire [7:0]    viotaResult_res_0_3 = compressVecPipe_12[7:0];
  wire [7:0]    viotaResult_res_1_3 = compressVecPipe_13[7:0];
  wire [7:0]    viotaResult_res_2_3 = compressVecPipe_14[7:0];
  wire [7:0]    viotaResult_res_3_3 = compressVecPipe_15[7:0];
  wire [15:0]   viotaResult_lo_3 = {viotaResult_res_1_3, viotaResult_res_0_3};
  wire [15:0]   viotaResult_hi_3 = {viotaResult_res_3_3, viotaResult_res_2_3};
  wire [7:0]    viotaResult_res_0_4 = compressVecPipe_16[7:0];
  wire [7:0]    viotaResult_res_1_4 = compressVecPipe_17[7:0];
  wire [7:0]    viotaResult_res_2_4 = compressVecPipe_18[7:0];
  wire [7:0]    viotaResult_res_3_4 = compressVecPipe_19[7:0];
  wire [15:0]   viotaResult_lo_4 = {viotaResult_res_1_4, viotaResult_res_0_4};
  wire [15:0]   viotaResult_hi_4 = {viotaResult_res_3_4, viotaResult_res_2_4};
  wire [7:0]    viotaResult_res_0_5 = compressVecPipe_20[7:0];
  wire [7:0]    viotaResult_res_1_5 = compressVecPipe_21[7:0];
  wire [7:0]    viotaResult_res_2_5 = compressVecPipe_22[7:0];
  wire [7:0]    viotaResult_res_3_5 = compressVecPipe_23[7:0];
  wire [15:0]   viotaResult_lo_5 = {viotaResult_res_1_5, viotaResult_res_0_5};
  wire [15:0]   viotaResult_hi_5 = {viotaResult_res_3_5, viotaResult_res_2_5};
  wire [7:0]    viotaResult_res_0_6 = compressVecPipe_24[7:0];
  wire [7:0]    viotaResult_res_1_6 = compressVecPipe_25[7:0];
  wire [7:0]    viotaResult_res_2_6 = compressVecPipe_26[7:0];
  wire [7:0]    viotaResult_res_3_6 = compressVecPipe_27[7:0];
  wire [15:0]   viotaResult_lo_6 = {viotaResult_res_1_6, viotaResult_res_0_6};
  wire [15:0]   viotaResult_hi_6 = {viotaResult_res_3_6, viotaResult_res_2_6};
  wire [7:0]    viotaResult_res_0_7 = compressVecPipe_28[7:0];
  wire [7:0]    viotaResult_res_1_7 = compressVecPipe_29[7:0];
  wire [7:0]    viotaResult_res_2_7 = compressVecPipe_30[7:0];
  wire [7:0]    viotaResult_res_3_7 = compressVecPipe_31[7:0];
  wire [15:0]   viotaResult_lo_7 = {viotaResult_res_1_7, viotaResult_res_0_7};
  wire [15:0]   viotaResult_hi_7 = {viotaResult_res_3_7, viotaResult_res_2_7};
  wire [7:0]    viotaResult_res_0_8 = compressVecPipe_32[7:0];
  wire [7:0]    viotaResult_res_1_8 = compressVecPipe_33[7:0];
  wire [7:0]    viotaResult_res_2_8 = compressVecPipe_34[7:0];
  wire [7:0]    viotaResult_res_3_8 = compressVecPipe_35[7:0];
  wire [15:0]   viotaResult_lo_8 = {viotaResult_res_1_8, viotaResult_res_0_8};
  wire [15:0]   viotaResult_hi_8 = {viotaResult_res_3_8, viotaResult_res_2_8};
  wire [7:0]    viotaResult_res_0_9 = compressVecPipe_36[7:0];
  wire [7:0]    viotaResult_res_1_9 = compressVecPipe_37[7:0];
  wire [7:0]    viotaResult_res_2_9 = compressVecPipe_38[7:0];
  wire [7:0]    viotaResult_res_3_9 = compressVecPipe_39[7:0];
  wire [15:0]   viotaResult_lo_9 = {viotaResult_res_1_9, viotaResult_res_0_9};
  wire [15:0]   viotaResult_hi_9 = {viotaResult_res_3_9, viotaResult_res_2_9};
  wire [7:0]    viotaResult_res_0_10 = compressVecPipe_40[7:0];
  wire [7:0]    viotaResult_res_1_10 = compressVecPipe_41[7:0];
  wire [7:0]    viotaResult_res_2_10 = compressVecPipe_42[7:0];
  wire [7:0]    viotaResult_res_3_10 = compressVecPipe_43[7:0];
  wire [15:0]   viotaResult_lo_10 = {viotaResult_res_1_10, viotaResult_res_0_10};
  wire [15:0]   viotaResult_hi_10 = {viotaResult_res_3_10, viotaResult_res_2_10};
  wire [7:0]    viotaResult_res_0_11 = compressVecPipe_44[7:0];
  wire [7:0]    viotaResult_res_1_11 = compressVecPipe_45[7:0];
  wire [7:0]    viotaResult_res_2_11 = compressVecPipe_46[7:0];
  wire [7:0]    viotaResult_res_3_11 = compressVecPipe_47[7:0];
  wire [15:0]   viotaResult_lo_11 = {viotaResult_res_1_11, viotaResult_res_0_11};
  wire [15:0]   viotaResult_hi_11 = {viotaResult_res_3_11, viotaResult_res_2_11};
  wire [7:0]    viotaResult_res_0_12 = compressVecPipe_48[7:0];
  wire [7:0]    viotaResult_res_1_12 = compressVecPipe_49[7:0];
  wire [7:0]    viotaResult_res_2_12 = compressVecPipe_50[7:0];
  wire [7:0]    viotaResult_res_3_12 = compressVecPipe_51[7:0];
  wire [15:0]   viotaResult_lo_12 = {viotaResult_res_1_12, viotaResult_res_0_12};
  wire [15:0]   viotaResult_hi_12 = {viotaResult_res_3_12, viotaResult_res_2_12};
  wire [7:0]    viotaResult_res_0_13 = compressVecPipe_52[7:0];
  wire [7:0]    viotaResult_res_1_13 = compressVecPipe_53[7:0];
  wire [7:0]    viotaResult_res_2_13 = compressVecPipe_54[7:0];
  wire [7:0]    viotaResult_res_3_13 = compressVecPipe_55[7:0];
  wire [15:0]   viotaResult_lo_13 = {viotaResult_res_1_13, viotaResult_res_0_13};
  wire [15:0]   viotaResult_hi_13 = {viotaResult_res_3_13, viotaResult_res_2_13};
  wire [7:0]    viotaResult_res_0_14 = compressVecPipe_56[7:0];
  wire [7:0]    viotaResult_res_1_14 = compressVecPipe_57[7:0];
  wire [7:0]    viotaResult_res_2_14 = compressVecPipe_58[7:0];
  wire [7:0]    viotaResult_res_3_14 = compressVecPipe_59[7:0];
  wire [15:0]   viotaResult_lo_14 = {viotaResult_res_1_14, viotaResult_res_0_14};
  wire [15:0]   viotaResult_hi_14 = {viotaResult_res_3_14, viotaResult_res_2_14};
  wire [7:0]    viotaResult_res_0_15 = compressVecPipe_60[7:0];
  wire [7:0]    viotaResult_res_1_15 = compressVecPipe_61[7:0];
  wire [7:0]    viotaResult_res_2_15 = compressVecPipe_62[7:0];
  wire [7:0]    viotaResult_res_3_15 = compressVecPipe_63[7:0];
  wire [15:0]   viotaResult_lo_15 = {viotaResult_res_1_15, viotaResult_res_0_15};
  wire [15:0]   viotaResult_hi_15 = {viotaResult_res_3_15, viotaResult_res_2_15};
  wire [63:0]   viotaResult_lo_lo_lo = {viotaResult_hi_1, viotaResult_lo_1, viotaResult_hi, viotaResult_lo};
  wire [63:0]   viotaResult_lo_lo_hi = {viotaResult_hi_3, viotaResult_lo_3, viotaResult_hi_2, viotaResult_lo_2};
  wire [127:0]  viotaResult_lo_lo = {viotaResult_lo_lo_hi, viotaResult_lo_lo_lo};
  wire [63:0]   viotaResult_lo_hi_lo = {viotaResult_hi_5, viotaResult_lo_5, viotaResult_hi_4, viotaResult_lo_4};
  wire [63:0]   viotaResult_lo_hi_hi = {viotaResult_hi_7, viotaResult_lo_7, viotaResult_hi_6, viotaResult_lo_6};
  wire [127:0]  viotaResult_lo_hi = {viotaResult_lo_hi_hi, viotaResult_lo_hi_lo};
  wire [255:0]  viotaResult_lo_16 = {viotaResult_lo_hi, viotaResult_lo_lo};
  wire [63:0]   viotaResult_hi_lo_lo = {viotaResult_hi_9, viotaResult_lo_9, viotaResult_hi_8, viotaResult_lo_8};
  wire [63:0]   viotaResult_hi_lo_hi = {viotaResult_hi_11, viotaResult_lo_11, viotaResult_hi_10, viotaResult_lo_10};
  wire [127:0]  viotaResult_hi_lo = {viotaResult_hi_lo_hi, viotaResult_hi_lo_lo};
  wire [63:0]   viotaResult_hi_hi_lo = {viotaResult_hi_13, viotaResult_lo_13, viotaResult_hi_12, viotaResult_lo_12};
  wire [63:0]   viotaResult_hi_hi_hi = {viotaResult_hi_15, viotaResult_lo_15, viotaResult_hi_14, viotaResult_lo_14};
  wire [127:0]  viotaResult_hi_hi = {viotaResult_hi_hi_hi, viotaResult_hi_hi_lo};
  wire [255:0]  viotaResult_hi_16 = {viotaResult_hi_hi, viotaResult_hi_lo};
  wire [15:0]   viotaResult_res_0_16 = {5'h0, compressVecPipe_0};
  wire [15:0]   viotaResult_res_1_16 = {5'h0, compressVecPipe_1};
  wire [15:0]   viotaResult_res_0_17 = {5'h0, compressVecPipe_2};
  wire [15:0]   viotaResult_res_1_17 = {5'h0, compressVecPipe_3};
  wire [15:0]   viotaResult_res_0_18 = {5'h0, compressVecPipe_4};
  wire [15:0]   viotaResult_res_1_18 = {5'h0, compressVecPipe_5};
  wire [15:0]   viotaResult_res_0_19 = {5'h0, compressVecPipe_6};
  wire [15:0]   viotaResult_res_1_19 = {5'h0, compressVecPipe_7};
  wire [15:0]   viotaResult_res_0_20 = {5'h0, compressVecPipe_8};
  wire [15:0]   viotaResult_res_1_20 = {5'h0, compressVecPipe_9};
  wire [15:0]   viotaResult_res_0_21 = {5'h0, compressVecPipe_10};
  wire [15:0]   viotaResult_res_1_21 = {5'h0, compressVecPipe_11};
  wire [15:0]   viotaResult_res_0_22 = {5'h0, compressVecPipe_12};
  wire [15:0]   viotaResult_res_1_22 = {5'h0, compressVecPipe_13};
  wire [15:0]   viotaResult_res_0_23 = {5'h0, compressVecPipe_14};
  wire [15:0]   viotaResult_res_1_23 = {5'h0, compressVecPipe_15};
  wire [15:0]   viotaResult_res_0_24 = {5'h0, compressVecPipe_16};
  wire [15:0]   viotaResult_res_1_24 = {5'h0, compressVecPipe_17};
  wire [15:0]   viotaResult_res_0_25 = {5'h0, compressVecPipe_18};
  wire [15:0]   viotaResult_res_1_25 = {5'h0, compressVecPipe_19};
  wire [15:0]   viotaResult_res_0_26 = {5'h0, compressVecPipe_20};
  wire [15:0]   viotaResult_res_1_26 = {5'h0, compressVecPipe_21};
  wire [15:0]   viotaResult_res_0_27 = {5'h0, compressVecPipe_22};
  wire [15:0]   viotaResult_res_1_27 = {5'h0, compressVecPipe_23};
  wire [15:0]   viotaResult_res_0_28 = {5'h0, compressVecPipe_24};
  wire [15:0]   viotaResult_res_1_28 = {5'h0, compressVecPipe_25};
  wire [15:0]   viotaResult_res_0_29 = {5'h0, compressVecPipe_26};
  wire [15:0]   viotaResult_res_1_29 = {5'h0, compressVecPipe_27};
  wire [15:0]   viotaResult_res_0_30 = {5'h0, compressVecPipe_28};
  wire [15:0]   viotaResult_res_1_30 = {5'h0, compressVecPipe_29};
  wire [15:0]   viotaResult_res_0_31 = {5'h0, compressVecPipe_30};
  wire [15:0]   viotaResult_res_1_31 = {5'h0, compressVecPipe_31};
  wire [63:0]   viotaResult_lo_lo_lo_1 = {viotaResult_res_1_17, viotaResult_res_0_17, viotaResult_res_1_16, viotaResult_res_0_16};
  wire [63:0]   viotaResult_lo_lo_hi_1 = {viotaResult_res_1_19, viotaResult_res_0_19, viotaResult_res_1_18, viotaResult_res_0_18};
  wire [127:0]  viotaResult_lo_lo_1 = {viotaResult_lo_lo_hi_1, viotaResult_lo_lo_lo_1};
  wire [63:0]   viotaResult_lo_hi_lo_1 = {viotaResult_res_1_21, viotaResult_res_0_21, viotaResult_res_1_20, viotaResult_res_0_20};
  wire [63:0]   viotaResult_lo_hi_hi_1 = {viotaResult_res_1_23, viotaResult_res_0_23, viotaResult_res_1_22, viotaResult_res_0_22};
  wire [127:0]  viotaResult_lo_hi_1 = {viotaResult_lo_hi_hi_1, viotaResult_lo_hi_lo_1};
  wire [255:0]  viotaResult_lo_17 = {viotaResult_lo_hi_1, viotaResult_lo_lo_1};
  wire [63:0]   viotaResult_hi_lo_lo_1 = {viotaResult_res_1_25, viotaResult_res_0_25, viotaResult_res_1_24, viotaResult_res_0_24};
  wire [63:0]   viotaResult_hi_lo_hi_1 = {viotaResult_res_1_27, viotaResult_res_0_27, viotaResult_res_1_26, viotaResult_res_0_26};
  wire [127:0]  viotaResult_hi_lo_1 = {viotaResult_hi_lo_hi_1, viotaResult_hi_lo_lo_1};
  wire [63:0]   viotaResult_hi_hi_lo_1 = {viotaResult_res_1_29, viotaResult_res_0_29, viotaResult_res_1_28, viotaResult_res_0_28};
  wire [63:0]   viotaResult_hi_hi_hi_1 = {viotaResult_res_1_31, viotaResult_res_0_31, viotaResult_res_1_30, viotaResult_res_0_30};
  wire [127:0]  viotaResult_hi_hi_1 = {viotaResult_hi_hi_hi_1, viotaResult_hi_hi_lo_1};
  wire [255:0]  viotaResult_hi_17 = {viotaResult_hi_hi_1, viotaResult_hi_lo_1};
  wire [31:0]   viotaResult_res_0_32 = {21'h0, compressVecPipe_0};
  wire [31:0]   viotaResult_res_0_33 = {21'h0, compressVecPipe_1};
  wire [31:0]   viotaResult_res_0_34 = {21'h0, compressVecPipe_2};
  wire [31:0]   viotaResult_res_0_35 = {21'h0, compressVecPipe_3};
  wire [31:0]   viotaResult_res_0_36 = {21'h0, compressVecPipe_4};
  wire [31:0]   viotaResult_res_0_37 = {21'h0, compressVecPipe_5};
  wire [31:0]   viotaResult_res_0_38 = {21'h0, compressVecPipe_6};
  wire [31:0]   viotaResult_res_0_39 = {21'h0, compressVecPipe_7};
  wire [31:0]   viotaResult_res_0_40 = {21'h0, compressVecPipe_8};
  wire [31:0]   viotaResult_res_0_41 = {21'h0, compressVecPipe_9};
  wire [31:0]   viotaResult_res_0_42 = {21'h0, compressVecPipe_10};
  wire [31:0]   viotaResult_res_0_43 = {21'h0, compressVecPipe_11};
  wire [31:0]   viotaResult_res_0_44 = {21'h0, compressVecPipe_12};
  wire [31:0]   viotaResult_res_0_45 = {21'h0, compressVecPipe_13};
  wire [31:0]   viotaResult_res_0_46 = {21'h0, compressVecPipe_14};
  wire [31:0]   viotaResult_res_0_47 = {21'h0, compressVecPipe_15};
  wire [63:0]   viotaResult_lo_lo_lo_2 = {viotaResult_res_0_33, viotaResult_res_0_32};
  wire [63:0]   viotaResult_lo_lo_hi_2 = {viotaResult_res_0_35, viotaResult_res_0_34};
  wire [127:0]  viotaResult_lo_lo_2 = {viotaResult_lo_lo_hi_2, viotaResult_lo_lo_lo_2};
  wire [63:0]   viotaResult_lo_hi_lo_2 = {viotaResult_res_0_37, viotaResult_res_0_36};
  wire [63:0]   viotaResult_lo_hi_hi_2 = {viotaResult_res_0_39, viotaResult_res_0_38};
  wire [127:0]  viotaResult_lo_hi_2 = {viotaResult_lo_hi_hi_2, viotaResult_lo_hi_lo_2};
  wire [255:0]  viotaResult_lo_18 = {viotaResult_lo_hi_2, viotaResult_lo_lo_2};
  wire [63:0]   viotaResult_hi_lo_lo_2 = {viotaResult_res_0_41, viotaResult_res_0_40};
  wire [63:0]   viotaResult_hi_lo_hi_2 = {viotaResult_res_0_43, viotaResult_res_0_42};
  wire [127:0]  viotaResult_hi_lo_2 = {viotaResult_hi_lo_hi_2, viotaResult_hi_lo_lo_2};
  wire [63:0]   viotaResult_hi_hi_lo_2 = {viotaResult_res_0_45, viotaResult_res_0_44};
  wire [63:0]   viotaResult_hi_hi_hi_2 = {viotaResult_res_0_47, viotaResult_res_0_46};
  wire [127:0]  viotaResult_hi_hi_2 = {viotaResult_hi_hi_hi_2, viotaResult_hi_hi_lo_2};
  wire [255:0]  viotaResult_hi_18 = {viotaResult_hi_hi_2, viotaResult_hi_lo_2};
  wire [511:0]  viotaResult = (eew1H[0] ? {viotaResult_hi_16, viotaResult_lo_16} : 512'h0) | (eew1H[1] ? {viotaResult_hi_17, viotaResult_lo_17} : 512'h0) | (eew1H[2] ? {viotaResult_hi_18, viotaResult_lo_18} : 512'h0);
  wire          viotaMask_res_0 = maskPipe[0];
  wire          viotaMask_res_1 = maskPipe[1];
  wire          viotaMask_res_2 = maskPipe[2];
  wire          viotaMask_res_3 = maskPipe[3];
  wire [1:0]    viotaMask_lo = {viotaMask_res_1, viotaMask_res_0};
  wire [1:0]    viotaMask_hi = {viotaMask_res_3, viotaMask_res_2};
  wire          viotaMask_res_0_1 = maskPipe[4];
  wire          viotaMask_res_1_1 = maskPipe[5];
  wire          viotaMask_res_2_1 = maskPipe[6];
  wire          viotaMask_res_3_1 = maskPipe[7];
  wire [1:0]    viotaMask_lo_1 = {viotaMask_res_1_1, viotaMask_res_0_1};
  wire [1:0]    viotaMask_hi_1 = {viotaMask_res_3_1, viotaMask_res_2_1};
  wire          viotaMask_res_0_2 = maskPipe[8];
  wire          viotaMask_res_1_2 = maskPipe[9];
  wire          viotaMask_res_2_2 = maskPipe[10];
  wire          viotaMask_res_3_2 = maskPipe[11];
  wire [1:0]    viotaMask_lo_2 = {viotaMask_res_1_2, viotaMask_res_0_2};
  wire [1:0]    viotaMask_hi_2 = {viotaMask_res_3_2, viotaMask_res_2_2};
  wire          viotaMask_res_0_3 = maskPipe[12];
  wire          viotaMask_res_1_3 = maskPipe[13];
  wire          viotaMask_res_2_3 = maskPipe[14];
  wire          viotaMask_res_3_3 = maskPipe[15];
  wire [1:0]    viotaMask_lo_3 = {viotaMask_res_1_3, viotaMask_res_0_3};
  wire [1:0]    viotaMask_hi_3 = {viotaMask_res_3_3, viotaMask_res_2_3};
  wire          viotaMask_res_0_4 = maskPipe[16];
  wire          viotaMask_res_1_4 = maskPipe[17];
  wire          viotaMask_res_2_4 = maskPipe[18];
  wire          viotaMask_res_3_4 = maskPipe[19];
  wire [1:0]    viotaMask_lo_4 = {viotaMask_res_1_4, viotaMask_res_0_4};
  wire [1:0]    viotaMask_hi_4 = {viotaMask_res_3_4, viotaMask_res_2_4};
  wire          viotaMask_res_0_5 = maskPipe[20];
  wire          viotaMask_res_1_5 = maskPipe[21];
  wire          viotaMask_res_2_5 = maskPipe[22];
  wire          viotaMask_res_3_5 = maskPipe[23];
  wire [1:0]    viotaMask_lo_5 = {viotaMask_res_1_5, viotaMask_res_0_5};
  wire [1:0]    viotaMask_hi_5 = {viotaMask_res_3_5, viotaMask_res_2_5};
  wire          viotaMask_res_0_6 = maskPipe[24];
  wire          viotaMask_res_1_6 = maskPipe[25];
  wire          viotaMask_res_2_6 = maskPipe[26];
  wire          viotaMask_res_3_6 = maskPipe[27];
  wire [1:0]    viotaMask_lo_6 = {viotaMask_res_1_6, viotaMask_res_0_6};
  wire [1:0]    viotaMask_hi_6 = {viotaMask_res_3_6, viotaMask_res_2_6};
  wire          viotaMask_res_0_7 = maskPipe[28];
  wire          viotaMask_res_1_7 = maskPipe[29];
  wire          viotaMask_res_2_7 = maskPipe[30];
  wire          viotaMask_res_3_7 = maskPipe[31];
  wire          viotaMask_res_0_8 = maskPipe[31];
  wire          viotaMask_res_1_8 = maskPipe[31];
  wire          viotaMask_res_2_8 = maskPipe[31];
  wire          viotaMask_res_3_8 = maskPipe[31];
  wire          viotaMask_res_0_9 = maskPipe[31];
  wire          viotaMask_res_1_9 = maskPipe[31];
  wire          viotaMask_res_2_9 = maskPipe[31];
  wire          viotaMask_res_3_9 = maskPipe[31];
  wire          viotaMask_res_0_10 = maskPipe[31];
  wire          viotaMask_res_1_10 = maskPipe[31];
  wire          viotaMask_res_2_10 = maskPipe[31];
  wire          viotaMask_res_3_10 = maskPipe[31];
  wire          viotaMask_res_0_11 = maskPipe[31];
  wire          viotaMask_res_1_11 = maskPipe[31];
  wire          viotaMask_res_2_11 = maskPipe[31];
  wire          viotaMask_res_3_11 = maskPipe[31];
  wire          viotaMask_res_0_12 = maskPipe[31];
  wire          viotaMask_res_1_12 = maskPipe[31];
  wire          viotaMask_res_2_12 = maskPipe[31];
  wire          viotaMask_res_3_12 = maskPipe[31];
  wire          viotaMask_res_0_13 = maskPipe[31];
  wire          viotaMask_res_1_13 = maskPipe[31];
  wire          viotaMask_res_2_13 = maskPipe[31];
  wire          viotaMask_res_3_13 = maskPipe[31];
  wire          viotaMask_res_0_14 = maskPipe[31];
  wire          viotaMask_res_1_14 = maskPipe[31];
  wire          viotaMask_res_2_14 = maskPipe[31];
  wire          viotaMask_res_3_14 = maskPipe[31];
  wire          viotaMask_res_0_15 = maskPipe[31];
  wire          viotaMask_res_1_15 = maskPipe[31];
  wire          viotaMask_res_2_15 = maskPipe[31];
  wire          viotaMask_res_3_15 = maskPipe[31];
  wire [1:0]    viotaMask_lo_7 = {viotaMask_res_1_7, viotaMask_res_0_7};
  wire [1:0]    viotaMask_hi_7 = {viotaMask_res_3_7, viotaMask_res_2_7};
  wire [1:0]    viotaMask_lo_8 = {viotaMask_res_1_8, viotaMask_res_0_8};
  wire [1:0]    viotaMask_hi_8 = {viotaMask_res_3_8, viotaMask_res_2_8};
  wire [1:0]    viotaMask_lo_9 = {viotaMask_res_1_9, viotaMask_res_0_9};
  wire [1:0]    viotaMask_hi_9 = {viotaMask_res_3_9, viotaMask_res_2_9};
  wire [1:0]    viotaMask_lo_10 = {viotaMask_res_1_10, viotaMask_res_0_10};
  wire [1:0]    viotaMask_hi_10 = {viotaMask_res_3_10, viotaMask_res_2_10};
  wire [1:0]    viotaMask_lo_11 = {viotaMask_res_1_11, viotaMask_res_0_11};
  wire [1:0]    viotaMask_hi_11 = {viotaMask_res_3_11, viotaMask_res_2_11};
  wire [1:0]    viotaMask_lo_12 = {viotaMask_res_1_12, viotaMask_res_0_12};
  wire [1:0]    viotaMask_hi_12 = {viotaMask_res_3_12, viotaMask_res_2_12};
  wire [1:0]    viotaMask_lo_13 = {viotaMask_res_1_13, viotaMask_res_0_13};
  wire [1:0]    viotaMask_hi_13 = {viotaMask_res_3_13, viotaMask_res_2_13};
  wire [1:0]    viotaMask_lo_14 = {viotaMask_res_1_14, viotaMask_res_0_14};
  wire [1:0]    viotaMask_hi_14 = {viotaMask_res_3_14, viotaMask_res_2_14};
  wire [1:0]    viotaMask_lo_15 = {viotaMask_res_1_15, viotaMask_res_0_15};
  wire [1:0]    viotaMask_hi_15 = {viotaMask_res_3_15, viotaMask_res_2_15};
  wire [7:0]    viotaMask_lo_lo_lo = {viotaMask_hi_1, viotaMask_lo_1, viotaMask_hi, viotaMask_lo};
  wire [7:0]    viotaMask_lo_lo_hi = {viotaMask_hi_3, viotaMask_lo_3, viotaMask_hi_2, viotaMask_lo_2};
  wire [15:0]   viotaMask_lo_lo = {viotaMask_lo_lo_hi, viotaMask_lo_lo_lo};
  wire [7:0]    viotaMask_lo_hi_lo = {viotaMask_hi_5, viotaMask_lo_5, viotaMask_hi_4, viotaMask_lo_4};
  wire [7:0]    viotaMask_lo_hi_hi = {viotaMask_hi_7, viotaMask_lo_7, viotaMask_hi_6, viotaMask_lo_6};
  wire [15:0]   viotaMask_lo_hi = {viotaMask_lo_hi_hi, viotaMask_lo_hi_lo};
  wire [31:0]   viotaMask_lo_16 = {viotaMask_lo_hi, viotaMask_lo_lo};
  wire [7:0]    viotaMask_hi_lo_lo = {viotaMask_hi_9, viotaMask_lo_9, viotaMask_hi_8, viotaMask_lo_8};
  wire [7:0]    viotaMask_hi_lo_hi = {viotaMask_hi_11, viotaMask_lo_11, viotaMask_hi_10, viotaMask_lo_10};
  wire [15:0]   viotaMask_hi_lo = {viotaMask_hi_lo_hi, viotaMask_hi_lo_lo};
  wire [7:0]    viotaMask_hi_hi_lo = {viotaMask_hi_13, viotaMask_lo_13, viotaMask_hi_12, viotaMask_lo_12};
  wire [7:0]    viotaMask_hi_hi_hi = {viotaMask_hi_15, viotaMask_lo_15, viotaMask_hi_14, viotaMask_lo_14};
  wire [15:0]   viotaMask_hi_hi = {viotaMask_hi_hi_hi, viotaMask_hi_hi_lo};
  wire [31:0]   viotaMask_hi_16 = {viotaMask_hi_hi, viotaMask_hi_lo};
  wire [1:0]    viotaMask_res_0_16 = {2{viotaMask_res_0}};
  wire [1:0]    viotaMask_res_1_16 = {2{viotaMask_res_1}};
  wire [1:0]    viotaMask_res_0_17 = {2{viotaMask_res_2}};
  wire [1:0]    viotaMask_res_1_17 = {2{viotaMask_res_3}};
  wire [1:0]    viotaMask_res_0_18 = {2{viotaMask_res_0_1}};
  wire [1:0]    viotaMask_res_1_18 = {2{viotaMask_res_1_1}};
  wire [1:0]    viotaMask_res_0_19 = {2{viotaMask_res_2_1}};
  wire [1:0]    viotaMask_res_1_19 = {2{viotaMask_res_3_1}};
  wire [1:0]    viotaMask_res_0_20 = {2{viotaMask_res_0_2}};
  wire [1:0]    viotaMask_res_1_20 = {2{viotaMask_res_1_2}};
  wire [1:0]    viotaMask_res_0_21 = {2{viotaMask_res_2_2}};
  wire [1:0]    viotaMask_res_1_21 = {2{viotaMask_res_3_2}};
  wire [1:0]    viotaMask_res_0_22 = {2{viotaMask_res_0_3}};
  wire [1:0]    viotaMask_res_1_22 = {2{viotaMask_res_1_3}};
  wire [1:0]    viotaMask_res_0_23 = {2{viotaMask_res_2_3}};
  wire [1:0]    viotaMask_res_1_23 = {2{viotaMask_res_3_3}};
  wire [1:0]    viotaMask_res_0_24 = {2{viotaMask_res_0_4}};
  wire [1:0]    viotaMask_res_1_24 = {2{viotaMask_res_1_4}};
  wire [1:0]    viotaMask_res_0_25 = {2{viotaMask_res_2_4}};
  wire [1:0]    viotaMask_res_1_25 = {2{viotaMask_res_3_4}};
  wire [1:0]    viotaMask_res_0_26 = {2{viotaMask_res_0_5}};
  wire [1:0]    viotaMask_res_1_26 = {2{viotaMask_res_1_5}};
  wire [1:0]    viotaMask_res_0_27 = {2{viotaMask_res_2_5}};
  wire [1:0]    viotaMask_res_1_27 = {2{viotaMask_res_3_5}};
  wire [1:0]    viotaMask_res_0_28 = {2{viotaMask_res_0_6}};
  wire [1:0]    viotaMask_res_1_28 = {2{viotaMask_res_1_6}};
  wire [1:0]    viotaMask_res_0_29 = {2{viotaMask_res_2_6}};
  wire [1:0]    viotaMask_res_1_29 = {2{viotaMask_res_3_6}};
  wire [1:0]    viotaMask_res_0_30 = {2{viotaMask_res_0_7}};
  wire [1:0]    viotaMask_res_1_30 = {2{viotaMask_res_1_7}};
  wire [1:0]    viotaMask_res_0_31 = {2{viotaMask_res_2_7}};
  wire [1:0]    viotaMask_res_1_31 = {2{maskPipe[31]}};
  wire [7:0]    viotaMask_lo_lo_lo_1 = {viotaMask_res_1_17, viotaMask_res_0_17, viotaMask_res_1_16, viotaMask_res_0_16};
  wire [7:0]    viotaMask_lo_lo_hi_1 = {viotaMask_res_1_19, viotaMask_res_0_19, viotaMask_res_1_18, viotaMask_res_0_18};
  wire [15:0]   viotaMask_lo_lo_1 = {viotaMask_lo_lo_hi_1, viotaMask_lo_lo_lo_1};
  wire [7:0]    viotaMask_lo_hi_lo_1 = {viotaMask_res_1_21, viotaMask_res_0_21, viotaMask_res_1_20, viotaMask_res_0_20};
  wire [7:0]    viotaMask_lo_hi_hi_1 = {viotaMask_res_1_23, viotaMask_res_0_23, viotaMask_res_1_22, viotaMask_res_0_22};
  wire [15:0]   viotaMask_lo_hi_1 = {viotaMask_lo_hi_hi_1, viotaMask_lo_hi_lo_1};
  wire [31:0]   viotaMask_lo_17 = {viotaMask_lo_hi_1, viotaMask_lo_lo_1};
  wire [7:0]    viotaMask_hi_lo_lo_1 = {viotaMask_res_1_25, viotaMask_res_0_25, viotaMask_res_1_24, viotaMask_res_0_24};
  wire [7:0]    viotaMask_hi_lo_hi_1 = {viotaMask_res_1_27, viotaMask_res_0_27, viotaMask_res_1_26, viotaMask_res_0_26};
  wire [15:0]   viotaMask_hi_lo_1 = {viotaMask_hi_lo_hi_1, viotaMask_hi_lo_lo_1};
  wire [7:0]    viotaMask_hi_hi_lo_1 = {viotaMask_res_1_29, viotaMask_res_0_29, viotaMask_res_1_28, viotaMask_res_0_28};
  wire [7:0]    viotaMask_hi_hi_hi_1 = {viotaMask_res_1_31, viotaMask_res_0_31, viotaMask_res_1_30, viotaMask_res_0_30};
  wire [15:0]   viotaMask_hi_hi_1 = {viotaMask_hi_hi_hi_1, viotaMask_hi_hi_lo_1};
  wire [31:0]   viotaMask_hi_17 = {viotaMask_hi_hi_1, viotaMask_hi_lo_1};
  wire [3:0]    viotaMask_res_0_32 = {4{viotaMask_res_0}};
  wire [3:0]    viotaMask_res_0_33 = {4{viotaMask_res_1}};
  wire [3:0]    viotaMask_res_0_34 = {4{viotaMask_res_2}};
  wire [3:0]    viotaMask_res_0_35 = {4{viotaMask_res_3}};
  wire [3:0]    viotaMask_res_0_36 = {4{viotaMask_res_0_1}};
  wire [3:0]    viotaMask_res_0_37 = {4{viotaMask_res_1_1}};
  wire [3:0]    viotaMask_res_0_38 = {4{viotaMask_res_2_1}};
  wire [3:0]    viotaMask_res_0_39 = {4{viotaMask_res_3_1}};
  wire [3:0]    viotaMask_res_0_40 = {4{viotaMask_res_0_2}};
  wire [3:0]    viotaMask_res_0_41 = {4{viotaMask_res_1_2}};
  wire [3:0]    viotaMask_res_0_42 = {4{viotaMask_res_2_2}};
  wire [3:0]    viotaMask_res_0_43 = {4{viotaMask_res_3_2}};
  wire [3:0]    viotaMask_res_0_44 = {4{viotaMask_res_0_3}};
  wire [3:0]    viotaMask_res_0_45 = {4{viotaMask_res_1_3}};
  wire [3:0]    viotaMask_res_0_46 = {4{viotaMask_res_2_3}};
  wire [3:0]    viotaMask_res_0_47 = {4{viotaMask_res_3_3}};
  wire [7:0]    viotaMask_lo_lo_lo_2 = {viotaMask_res_0_33, viotaMask_res_0_32};
  wire [7:0]    viotaMask_lo_lo_hi_2 = {viotaMask_res_0_35, viotaMask_res_0_34};
  wire [15:0]   viotaMask_lo_lo_2 = {viotaMask_lo_lo_hi_2, viotaMask_lo_lo_lo_2};
  wire [7:0]    viotaMask_lo_hi_lo_2 = {viotaMask_res_0_37, viotaMask_res_0_36};
  wire [7:0]    viotaMask_lo_hi_hi_2 = {viotaMask_res_0_39, viotaMask_res_0_38};
  wire [15:0]   viotaMask_lo_hi_2 = {viotaMask_lo_hi_hi_2, viotaMask_lo_hi_lo_2};
  wire [31:0]   viotaMask_lo_18 = {viotaMask_lo_hi_2, viotaMask_lo_lo_2};
  wire [7:0]    viotaMask_hi_lo_lo_2 = {viotaMask_res_0_41, viotaMask_res_0_40};
  wire [7:0]    viotaMask_hi_lo_hi_2 = {viotaMask_res_0_43, viotaMask_res_0_42};
  wire [15:0]   viotaMask_hi_lo_2 = {viotaMask_hi_lo_hi_2, viotaMask_hi_lo_lo_2};
  wire [7:0]    viotaMask_hi_hi_lo_2 = {viotaMask_res_0_45, viotaMask_res_0_44};
  wire [7:0]    viotaMask_hi_hi_hi_2 = {viotaMask_res_0_47, viotaMask_res_0_46};
  wire [15:0]   viotaMask_hi_hi_2 = {viotaMask_hi_hi_hi_2, viotaMask_hi_hi_lo_2};
  wire [31:0]   viotaMask_hi_18 = {viotaMask_hi_hi_2, viotaMask_hi_lo_2};
  wire [63:0]   viotaMask = (eew1H[0] ? {viotaMask_hi_16, viotaMask_lo_16} : 64'h0) | (eew1H[1] ? {viotaMask_hi_17, viotaMask_lo_17} : 64'h0) | (eew1H[2] ? {viotaMask_hi_18, viotaMask_lo_18} : 64'h0);
  wire [5:0]    tailCount = compressInitPipe[5:0];
  wire [5:0]    tailCountForMask = compressInit[5:0];
  reg  [511:0]  compressDataReg;
  reg           compressTailValid;
  reg  [5:0]    compressWriteGroupCount;
  wire          _GEN_0 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h0;
  wire          compressDataVec_hitReq_0;
  assign compressDataVec_hitReq_0 = _GEN_0;
  wire          compressDataVec_hitReq_0_128;
  assign compressDataVec_hitReq_0_128 = _GEN_0;
  wire          compressDataVec_hitReq_0_192;
  assign compressDataVec_hitReq_0_192 = _GEN_0;
  wire          _GEN_1 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h0;
  wire          compressDataVec_hitReq_1;
  assign compressDataVec_hitReq_1 = _GEN_1;
  wire          compressDataVec_hitReq_1_128;
  assign compressDataVec_hitReq_1_128 = _GEN_1;
  wire          compressDataVec_hitReq_1_192;
  assign compressDataVec_hitReq_1_192 = _GEN_1;
  wire          _GEN_2 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h0;
  wire          compressDataVec_hitReq_2;
  assign compressDataVec_hitReq_2 = _GEN_2;
  wire          compressDataVec_hitReq_2_128;
  assign compressDataVec_hitReq_2_128 = _GEN_2;
  wire          compressDataVec_hitReq_2_192;
  assign compressDataVec_hitReq_2_192 = _GEN_2;
  wire          _GEN_3 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h0;
  wire          compressDataVec_hitReq_3;
  assign compressDataVec_hitReq_3 = _GEN_3;
  wire          compressDataVec_hitReq_3_128;
  assign compressDataVec_hitReq_3_128 = _GEN_3;
  wire          compressDataVec_hitReq_3_192;
  assign compressDataVec_hitReq_3_192 = _GEN_3;
  wire          _GEN_4 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h0;
  wire          compressDataVec_hitReq_4;
  assign compressDataVec_hitReq_4 = _GEN_4;
  wire          compressDataVec_hitReq_4_128;
  assign compressDataVec_hitReq_4_128 = _GEN_4;
  wire          compressDataVec_hitReq_4_192;
  assign compressDataVec_hitReq_4_192 = _GEN_4;
  wire          _GEN_5 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h0;
  wire          compressDataVec_hitReq_5;
  assign compressDataVec_hitReq_5 = _GEN_5;
  wire          compressDataVec_hitReq_5_128;
  assign compressDataVec_hitReq_5_128 = _GEN_5;
  wire          compressDataVec_hitReq_5_192;
  assign compressDataVec_hitReq_5_192 = _GEN_5;
  wire          _GEN_6 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h0;
  wire          compressDataVec_hitReq_6;
  assign compressDataVec_hitReq_6 = _GEN_6;
  wire          compressDataVec_hitReq_6_128;
  assign compressDataVec_hitReq_6_128 = _GEN_6;
  wire          compressDataVec_hitReq_6_192;
  assign compressDataVec_hitReq_6_192 = _GEN_6;
  wire          _GEN_7 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h0;
  wire          compressDataVec_hitReq_7;
  assign compressDataVec_hitReq_7 = _GEN_7;
  wire          compressDataVec_hitReq_7_128;
  assign compressDataVec_hitReq_7_128 = _GEN_7;
  wire          compressDataVec_hitReq_7_192;
  assign compressDataVec_hitReq_7_192 = _GEN_7;
  wire          _GEN_8 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h0;
  wire          compressDataVec_hitReq_8;
  assign compressDataVec_hitReq_8 = _GEN_8;
  wire          compressDataVec_hitReq_8_128;
  assign compressDataVec_hitReq_8_128 = _GEN_8;
  wire          compressDataVec_hitReq_8_192;
  assign compressDataVec_hitReq_8_192 = _GEN_8;
  wire          _GEN_9 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h0;
  wire          compressDataVec_hitReq_9;
  assign compressDataVec_hitReq_9 = _GEN_9;
  wire          compressDataVec_hitReq_9_128;
  assign compressDataVec_hitReq_9_128 = _GEN_9;
  wire          compressDataVec_hitReq_9_192;
  assign compressDataVec_hitReq_9_192 = _GEN_9;
  wire          _GEN_10 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h0;
  wire          compressDataVec_hitReq_10;
  assign compressDataVec_hitReq_10 = _GEN_10;
  wire          compressDataVec_hitReq_10_128;
  assign compressDataVec_hitReq_10_128 = _GEN_10;
  wire          compressDataVec_hitReq_10_192;
  assign compressDataVec_hitReq_10_192 = _GEN_10;
  wire          _GEN_11 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h0;
  wire          compressDataVec_hitReq_11;
  assign compressDataVec_hitReq_11 = _GEN_11;
  wire          compressDataVec_hitReq_11_128;
  assign compressDataVec_hitReq_11_128 = _GEN_11;
  wire          compressDataVec_hitReq_11_192;
  assign compressDataVec_hitReq_11_192 = _GEN_11;
  wire          _GEN_12 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h0;
  wire          compressDataVec_hitReq_12;
  assign compressDataVec_hitReq_12 = _GEN_12;
  wire          compressDataVec_hitReq_12_128;
  assign compressDataVec_hitReq_12_128 = _GEN_12;
  wire          compressDataVec_hitReq_12_192;
  assign compressDataVec_hitReq_12_192 = _GEN_12;
  wire          _GEN_13 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h0;
  wire          compressDataVec_hitReq_13;
  assign compressDataVec_hitReq_13 = _GEN_13;
  wire          compressDataVec_hitReq_13_128;
  assign compressDataVec_hitReq_13_128 = _GEN_13;
  wire          compressDataVec_hitReq_13_192;
  assign compressDataVec_hitReq_13_192 = _GEN_13;
  wire          _GEN_14 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h0;
  wire          compressDataVec_hitReq_14;
  assign compressDataVec_hitReq_14 = _GEN_14;
  wire          compressDataVec_hitReq_14_128;
  assign compressDataVec_hitReq_14_128 = _GEN_14;
  wire          compressDataVec_hitReq_14_192;
  assign compressDataVec_hitReq_14_192 = _GEN_14;
  wire          _GEN_15 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h0;
  wire          compressDataVec_hitReq_15;
  assign compressDataVec_hitReq_15 = _GEN_15;
  wire          compressDataVec_hitReq_15_128;
  assign compressDataVec_hitReq_15_128 = _GEN_15;
  wire          compressDataVec_hitReq_15_192;
  assign compressDataVec_hitReq_15_192 = _GEN_15;
  wire          _GEN_16 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h0;
  wire          compressDataVec_hitReq_16;
  assign compressDataVec_hitReq_16 = _GEN_16;
  wire          compressDataVec_hitReq_16_128;
  assign compressDataVec_hitReq_16_128 = _GEN_16;
  wire          _GEN_17 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h0;
  wire          compressDataVec_hitReq_17;
  assign compressDataVec_hitReq_17 = _GEN_17;
  wire          compressDataVec_hitReq_17_128;
  assign compressDataVec_hitReq_17_128 = _GEN_17;
  wire          _GEN_18 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h0;
  wire          compressDataVec_hitReq_18;
  assign compressDataVec_hitReq_18 = _GEN_18;
  wire          compressDataVec_hitReq_18_128;
  assign compressDataVec_hitReq_18_128 = _GEN_18;
  wire          _GEN_19 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h0;
  wire          compressDataVec_hitReq_19;
  assign compressDataVec_hitReq_19 = _GEN_19;
  wire          compressDataVec_hitReq_19_128;
  assign compressDataVec_hitReq_19_128 = _GEN_19;
  wire          _GEN_20 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h0;
  wire          compressDataVec_hitReq_20;
  assign compressDataVec_hitReq_20 = _GEN_20;
  wire          compressDataVec_hitReq_20_128;
  assign compressDataVec_hitReq_20_128 = _GEN_20;
  wire          _GEN_21 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h0;
  wire          compressDataVec_hitReq_21;
  assign compressDataVec_hitReq_21 = _GEN_21;
  wire          compressDataVec_hitReq_21_128;
  assign compressDataVec_hitReq_21_128 = _GEN_21;
  wire          _GEN_22 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h0;
  wire          compressDataVec_hitReq_22;
  assign compressDataVec_hitReq_22 = _GEN_22;
  wire          compressDataVec_hitReq_22_128;
  assign compressDataVec_hitReq_22_128 = _GEN_22;
  wire          _GEN_23 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h0;
  wire          compressDataVec_hitReq_23;
  assign compressDataVec_hitReq_23 = _GEN_23;
  wire          compressDataVec_hitReq_23_128;
  assign compressDataVec_hitReq_23_128 = _GEN_23;
  wire          _GEN_24 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h0;
  wire          compressDataVec_hitReq_24;
  assign compressDataVec_hitReq_24 = _GEN_24;
  wire          compressDataVec_hitReq_24_128;
  assign compressDataVec_hitReq_24_128 = _GEN_24;
  wire          _GEN_25 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h0;
  wire          compressDataVec_hitReq_25;
  assign compressDataVec_hitReq_25 = _GEN_25;
  wire          compressDataVec_hitReq_25_128;
  assign compressDataVec_hitReq_25_128 = _GEN_25;
  wire          _GEN_26 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h0;
  wire          compressDataVec_hitReq_26;
  assign compressDataVec_hitReq_26 = _GEN_26;
  wire          compressDataVec_hitReq_26_128;
  assign compressDataVec_hitReq_26_128 = _GEN_26;
  wire          _GEN_27 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h0;
  wire          compressDataVec_hitReq_27;
  assign compressDataVec_hitReq_27 = _GEN_27;
  wire          compressDataVec_hitReq_27_128;
  assign compressDataVec_hitReq_27_128 = _GEN_27;
  wire          _GEN_28 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h0;
  wire          compressDataVec_hitReq_28;
  assign compressDataVec_hitReq_28 = _GEN_28;
  wire          compressDataVec_hitReq_28_128;
  assign compressDataVec_hitReq_28_128 = _GEN_28;
  wire          _GEN_29 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h0;
  wire          compressDataVec_hitReq_29;
  assign compressDataVec_hitReq_29 = _GEN_29;
  wire          compressDataVec_hitReq_29_128;
  assign compressDataVec_hitReq_29_128 = _GEN_29;
  wire          _GEN_30 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h0;
  wire          compressDataVec_hitReq_30;
  assign compressDataVec_hitReq_30 = _GEN_30;
  wire          compressDataVec_hitReq_30_128;
  assign compressDataVec_hitReq_30_128 = _GEN_30;
  wire          _GEN_31 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h0;
  wire          compressDataVec_hitReq_31;
  assign compressDataVec_hitReq_31 = _GEN_31;
  wire          compressDataVec_hitReq_31_128;
  assign compressDataVec_hitReq_31_128 = _GEN_31;
  wire          compressDataVec_hitReq_32 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h0;
  wire          compressDataVec_hitReq_33 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h0;
  wire          compressDataVec_hitReq_34 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h0;
  wire          compressDataVec_hitReq_35 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h0;
  wire          compressDataVec_hitReq_36 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h0;
  wire          compressDataVec_hitReq_37 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h0;
  wire          compressDataVec_hitReq_38 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h0;
  wire          compressDataVec_hitReq_39 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h0;
  wire          compressDataVec_hitReq_40 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h0;
  wire          compressDataVec_hitReq_41 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h0;
  wire          compressDataVec_hitReq_42 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h0;
  wire          compressDataVec_hitReq_43 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h0;
  wire          compressDataVec_hitReq_44 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h0;
  wire          compressDataVec_hitReq_45 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h0;
  wire          compressDataVec_hitReq_46 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h0;
  wire          compressDataVec_hitReq_47 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h0;
  wire          compressDataVec_hitReq_48 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h0;
  wire          compressDataVec_hitReq_49 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h0;
  wire          compressDataVec_hitReq_50 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h0;
  wire          compressDataVec_hitReq_51 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h0;
  wire          compressDataVec_hitReq_52 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h0;
  wire          compressDataVec_hitReq_53 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h0;
  wire          compressDataVec_hitReq_54 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h0;
  wire          compressDataVec_hitReq_55 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h0;
  wire          compressDataVec_hitReq_56 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h0;
  wire          compressDataVec_hitReq_57 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h0;
  wire          compressDataVec_hitReq_58 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h0;
  wire          compressDataVec_hitReq_59 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h0;
  wire          compressDataVec_hitReq_60 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h0;
  wire          compressDataVec_hitReq_61 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h0;
  wire          compressDataVec_hitReq_62 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h0;
  wire          compressDataVec_hitReq_63 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h0;
  wire [7:0]    compressDataVec_selectReqData =
    (compressDataVec_hitReq_0 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7 ? source2Pipe[63:56] : 8'h0)
    | (compressDataVec_hitReq_8 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11 ? source2Pipe[95:88] : 8'h0)
    | (compressDataVec_hitReq_12 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14 ? source2Pipe[119:112] : 8'h0)
    | (compressDataVec_hitReq_15 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17 ? source2Pipe[143:136] : 8'h0)
    | (compressDataVec_hitReq_18 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20 ? source2Pipe[167:160] : 8'h0)
    | (compressDataVec_hitReq_21 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23 ? source2Pipe[191:184] : 8'h0)
    | (compressDataVec_hitReq_24 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26 ? source2Pipe[215:208] : 8'h0)
    | (compressDataVec_hitReq_27 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29 ? source2Pipe[239:232] : 8'h0)
    | (compressDataVec_hitReq_30 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32 ? source2Pipe[263:256] : 8'h0)
    | (compressDataVec_hitReq_33 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35 ? source2Pipe[287:280] : 8'h0)
    | (compressDataVec_hitReq_36 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38 ? source2Pipe[311:304] : 8'h0)
    | (compressDataVec_hitReq_39 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41 ? source2Pipe[335:328] : 8'h0)
    | (compressDataVec_hitReq_42 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44 ? source2Pipe[359:352] : 8'h0)
    | (compressDataVec_hitReq_45 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47 ? source2Pipe[383:376] : 8'h0)
    | (compressDataVec_hitReq_48 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50 ? source2Pipe[407:400] : 8'h0)
    | (compressDataVec_hitReq_51 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53 ? source2Pipe[431:424] : 8'h0)
    | (compressDataVec_hitReq_54 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56 ? source2Pipe[455:448] : 8'h0)
    | (compressDataVec_hitReq_57 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59 ? source2Pipe[479:472] : 8'h0)
    | (compressDataVec_hitReq_60 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62 ? source2Pipe[503:496] : 8'h0)
    | (compressDataVec_hitReq_63 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail;
  assign compressDataVec_useTail = |tailCount;
  wire          _GEN_32 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h1;
  wire          compressDataVec_hitReq_0_1;
  assign compressDataVec_hitReq_0_1 = _GEN_32;
  wire          compressDataVec_hitReq_0_129;
  assign compressDataVec_hitReq_0_129 = _GEN_32;
  wire          compressDataVec_hitReq_0_193;
  assign compressDataVec_hitReq_0_193 = _GEN_32;
  wire          _GEN_33 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h1;
  wire          compressDataVec_hitReq_1_1;
  assign compressDataVec_hitReq_1_1 = _GEN_33;
  wire          compressDataVec_hitReq_1_129;
  assign compressDataVec_hitReq_1_129 = _GEN_33;
  wire          compressDataVec_hitReq_1_193;
  assign compressDataVec_hitReq_1_193 = _GEN_33;
  wire          _GEN_34 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h1;
  wire          compressDataVec_hitReq_2_1;
  assign compressDataVec_hitReq_2_1 = _GEN_34;
  wire          compressDataVec_hitReq_2_129;
  assign compressDataVec_hitReq_2_129 = _GEN_34;
  wire          compressDataVec_hitReq_2_193;
  assign compressDataVec_hitReq_2_193 = _GEN_34;
  wire          _GEN_35 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h1;
  wire          compressDataVec_hitReq_3_1;
  assign compressDataVec_hitReq_3_1 = _GEN_35;
  wire          compressDataVec_hitReq_3_129;
  assign compressDataVec_hitReq_3_129 = _GEN_35;
  wire          compressDataVec_hitReq_3_193;
  assign compressDataVec_hitReq_3_193 = _GEN_35;
  wire          _GEN_36 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h1;
  wire          compressDataVec_hitReq_4_1;
  assign compressDataVec_hitReq_4_1 = _GEN_36;
  wire          compressDataVec_hitReq_4_129;
  assign compressDataVec_hitReq_4_129 = _GEN_36;
  wire          compressDataVec_hitReq_4_193;
  assign compressDataVec_hitReq_4_193 = _GEN_36;
  wire          _GEN_37 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h1;
  wire          compressDataVec_hitReq_5_1;
  assign compressDataVec_hitReq_5_1 = _GEN_37;
  wire          compressDataVec_hitReq_5_129;
  assign compressDataVec_hitReq_5_129 = _GEN_37;
  wire          compressDataVec_hitReq_5_193;
  assign compressDataVec_hitReq_5_193 = _GEN_37;
  wire          _GEN_38 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h1;
  wire          compressDataVec_hitReq_6_1;
  assign compressDataVec_hitReq_6_1 = _GEN_38;
  wire          compressDataVec_hitReq_6_129;
  assign compressDataVec_hitReq_6_129 = _GEN_38;
  wire          compressDataVec_hitReq_6_193;
  assign compressDataVec_hitReq_6_193 = _GEN_38;
  wire          _GEN_39 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h1;
  wire          compressDataVec_hitReq_7_1;
  assign compressDataVec_hitReq_7_1 = _GEN_39;
  wire          compressDataVec_hitReq_7_129;
  assign compressDataVec_hitReq_7_129 = _GEN_39;
  wire          compressDataVec_hitReq_7_193;
  assign compressDataVec_hitReq_7_193 = _GEN_39;
  wire          _GEN_40 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h1;
  wire          compressDataVec_hitReq_8_1;
  assign compressDataVec_hitReq_8_1 = _GEN_40;
  wire          compressDataVec_hitReq_8_129;
  assign compressDataVec_hitReq_8_129 = _GEN_40;
  wire          compressDataVec_hitReq_8_193;
  assign compressDataVec_hitReq_8_193 = _GEN_40;
  wire          _GEN_41 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h1;
  wire          compressDataVec_hitReq_9_1;
  assign compressDataVec_hitReq_9_1 = _GEN_41;
  wire          compressDataVec_hitReq_9_129;
  assign compressDataVec_hitReq_9_129 = _GEN_41;
  wire          compressDataVec_hitReq_9_193;
  assign compressDataVec_hitReq_9_193 = _GEN_41;
  wire          _GEN_42 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h1;
  wire          compressDataVec_hitReq_10_1;
  assign compressDataVec_hitReq_10_1 = _GEN_42;
  wire          compressDataVec_hitReq_10_129;
  assign compressDataVec_hitReq_10_129 = _GEN_42;
  wire          compressDataVec_hitReq_10_193;
  assign compressDataVec_hitReq_10_193 = _GEN_42;
  wire          _GEN_43 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h1;
  wire          compressDataVec_hitReq_11_1;
  assign compressDataVec_hitReq_11_1 = _GEN_43;
  wire          compressDataVec_hitReq_11_129;
  assign compressDataVec_hitReq_11_129 = _GEN_43;
  wire          compressDataVec_hitReq_11_193;
  assign compressDataVec_hitReq_11_193 = _GEN_43;
  wire          _GEN_44 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h1;
  wire          compressDataVec_hitReq_12_1;
  assign compressDataVec_hitReq_12_1 = _GEN_44;
  wire          compressDataVec_hitReq_12_129;
  assign compressDataVec_hitReq_12_129 = _GEN_44;
  wire          compressDataVec_hitReq_12_193;
  assign compressDataVec_hitReq_12_193 = _GEN_44;
  wire          _GEN_45 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h1;
  wire          compressDataVec_hitReq_13_1;
  assign compressDataVec_hitReq_13_1 = _GEN_45;
  wire          compressDataVec_hitReq_13_129;
  assign compressDataVec_hitReq_13_129 = _GEN_45;
  wire          compressDataVec_hitReq_13_193;
  assign compressDataVec_hitReq_13_193 = _GEN_45;
  wire          _GEN_46 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h1;
  wire          compressDataVec_hitReq_14_1;
  assign compressDataVec_hitReq_14_1 = _GEN_46;
  wire          compressDataVec_hitReq_14_129;
  assign compressDataVec_hitReq_14_129 = _GEN_46;
  wire          compressDataVec_hitReq_14_193;
  assign compressDataVec_hitReq_14_193 = _GEN_46;
  wire          _GEN_47 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h1;
  wire          compressDataVec_hitReq_15_1;
  assign compressDataVec_hitReq_15_1 = _GEN_47;
  wire          compressDataVec_hitReq_15_129;
  assign compressDataVec_hitReq_15_129 = _GEN_47;
  wire          compressDataVec_hitReq_15_193;
  assign compressDataVec_hitReq_15_193 = _GEN_47;
  wire          _GEN_48 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h1;
  wire          compressDataVec_hitReq_16_1;
  assign compressDataVec_hitReq_16_1 = _GEN_48;
  wire          compressDataVec_hitReq_16_129;
  assign compressDataVec_hitReq_16_129 = _GEN_48;
  wire          _GEN_49 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h1;
  wire          compressDataVec_hitReq_17_1;
  assign compressDataVec_hitReq_17_1 = _GEN_49;
  wire          compressDataVec_hitReq_17_129;
  assign compressDataVec_hitReq_17_129 = _GEN_49;
  wire          _GEN_50 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h1;
  wire          compressDataVec_hitReq_18_1;
  assign compressDataVec_hitReq_18_1 = _GEN_50;
  wire          compressDataVec_hitReq_18_129;
  assign compressDataVec_hitReq_18_129 = _GEN_50;
  wire          _GEN_51 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h1;
  wire          compressDataVec_hitReq_19_1;
  assign compressDataVec_hitReq_19_1 = _GEN_51;
  wire          compressDataVec_hitReq_19_129;
  assign compressDataVec_hitReq_19_129 = _GEN_51;
  wire          _GEN_52 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h1;
  wire          compressDataVec_hitReq_20_1;
  assign compressDataVec_hitReq_20_1 = _GEN_52;
  wire          compressDataVec_hitReq_20_129;
  assign compressDataVec_hitReq_20_129 = _GEN_52;
  wire          _GEN_53 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h1;
  wire          compressDataVec_hitReq_21_1;
  assign compressDataVec_hitReq_21_1 = _GEN_53;
  wire          compressDataVec_hitReq_21_129;
  assign compressDataVec_hitReq_21_129 = _GEN_53;
  wire          _GEN_54 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h1;
  wire          compressDataVec_hitReq_22_1;
  assign compressDataVec_hitReq_22_1 = _GEN_54;
  wire          compressDataVec_hitReq_22_129;
  assign compressDataVec_hitReq_22_129 = _GEN_54;
  wire          _GEN_55 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h1;
  wire          compressDataVec_hitReq_23_1;
  assign compressDataVec_hitReq_23_1 = _GEN_55;
  wire          compressDataVec_hitReq_23_129;
  assign compressDataVec_hitReq_23_129 = _GEN_55;
  wire          _GEN_56 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h1;
  wire          compressDataVec_hitReq_24_1;
  assign compressDataVec_hitReq_24_1 = _GEN_56;
  wire          compressDataVec_hitReq_24_129;
  assign compressDataVec_hitReq_24_129 = _GEN_56;
  wire          _GEN_57 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h1;
  wire          compressDataVec_hitReq_25_1;
  assign compressDataVec_hitReq_25_1 = _GEN_57;
  wire          compressDataVec_hitReq_25_129;
  assign compressDataVec_hitReq_25_129 = _GEN_57;
  wire          _GEN_58 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h1;
  wire          compressDataVec_hitReq_26_1;
  assign compressDataVec_hitReq_26_1 = _GEN_58;
  wire          compressDataVec_hitReq_26_129;
  assign compressDataVec_hitReq_26_129 = _GEN_58;
  wire          _GEN_59 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h1;
  wire          compressDataVec_hitReq_27_1;
  assign compressDataVec_hitReq_27_1 = _GEN_59;
  wire          compressDataVec_hitReq_27_129;
  assign compressDataVec_hitReq_27_129 = _GEN_59;
  wire          _GEN_60 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h1;
  wire          compressDataVec_hitReq_28_1;
  assign compressDataVec_hitReq_28_1 = _GEN_60;
  wire          compressDataVec_hitReq_28_129;
  assign compressDataVec_hitReq_28_129 = _GEN_60;
  wire          _GEN_61 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h1;
  wire          compressDataVec_hitReq_29_1;
  assign compressDataVec_hitReq_29_1 = _GEN_61;
  wire          compressDataVec_hitReq_29_129;
  assign compressDataVec_hitReq_29_129 = _GEN_61;
  wire          _GEN_62 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h1;
  wire          compressDataVec_hitReq_30_1;
  assign compressDataVec_hitReq_30_1 = _GEN_62;
  wire          compressDataVec_hitReq_30_129;
  assign compressDataVec_hitReq_30_129 = _GEN_62;
  wire          _GEN_63 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h1;
  wire          compressDataVec_hitReq_31_1;
  assign compressDataVec_hitReq_31_1 = _GEN_63;
  wire          compressDataVec_hitReq_31_129;
  assign compressDataVec_hitReq_31_129 = _GEN_63;
  wire          compressDataVec_hitReq_32_1 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h1;
  wire          compressDataVec_hitReq_33_1 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h1;
  wire          compressDataVec_hitReq_34_1 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h1;
  wire          compressDataVec_hitReq_35_1 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h1;
  wire          compressDataVec_hitReq_36_1 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h1;
  wire          compressDataVec_hitReq_37_1 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h1;
  wire          compressDataVec_hitReq_38_1 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h1;
  wire          compressDataVec_hitReq_39_1 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h1;
  wire          compressDataVec_hitReq_40_1 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h1;
  wire          compressDataVec_hitReq_41_1 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h1;
  wire          compressDataVec_hitReq_42_1 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h1;
  wire          compressDataVec_hitReq_43_1 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h1;
  wire          compressDataVec_hitReq_44_1 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h1;
  wire          compressDataVec_hitReq_45_1 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h1;
  wire          compressDataVec_hitReq_46_1 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h1;
  wire          compressDataVec_hitReq_47_1 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h1;
  wire          compressDataVec_hitReq_48_1 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h1;
  wire          compressDataVec_hitReq_49_1 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h1;
  wire          compressDataVec_hitReq_50_1 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h1;
  wire          compressDataVec_hitReq_51_1 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h1;
  wire          compressDataVec_hitReq_52_1 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h1;
  wire          compressDataVec_hitReq_53_1 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h1;
  wire          compressDataVec_hitReq_54_1 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h1;
  wire          compressDataVec_hitReq_55_1 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h1;
  wire          compressDataVec_hitReq_56_1 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h1;
  wire          compressDataVec_hitReq_57_1 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h1;
  wire          compressDataVec_hitReq_58_1 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h1;
  wire          compressDataVec_hitReq_59_1 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h1;
  wire          compressDataVec_hitReq_60_1 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h1;
  wire          compressDataVec_hitReq_61_1 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h1;
  wire          compressDataVec_hitReq_62_1 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h1;
  wire          compressDataVec_hitReq_63_1 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h1;
  wire [7:0]    compressDataVec_selectReqData_1 =
    (compressDataVec_hitReq_0_1 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_1 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_1 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_1 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_1 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_1 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_1 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_1 ? source2Pipe[63:56] : 8'h0)
    | (compressDataVec_hitReq_8_1 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_1 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_1 ? source2Pipe[87:80] : 8'h0)
    | (compressDataVec_hitReq_11_1 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_1 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_1 ? source2Pipe[111:104] : 8'h0)
    | (compressDataVec_hitReq_14_1 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_1 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_1 ? source2Pipe[135:128] : 8'h0)
    | (compressDataVec_hitReq_17_1 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_1 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_1 ? source2Pipe[159:152] : 8'h0)
    | (compressDataVec_hitReq_20_1 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_1 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_1 ? source2Pipe[183:176] : 8'h0)
    | (compressDataVec_hitReq_23_1 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_1 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_1 ? source2Pipe[207:200] : 8'h0)
    | (compressDataVec_hitReq_26_1 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_1 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_1 ? source2Pipe[231:224] : 8'h0)
    | (compressDataVec_hitReq_29_1 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_1 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_1 ? source2Pipe[255:248] : 8'h0)
    | (compressDataVec_hitReq_32_1 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_1 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_1 ? source2Pipe[279:272] : 8'h0)
    | (compressDataVec_hitReq_35_1 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_1 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_1 ? source2Pipe[303:296] : 8'h0)
    | (compressDataVec_hitReq_38_1 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_1 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_1 ? source2Pipe[327:320] : 8'h0)
    | (compressDataVec_hitReq_41_1 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_1 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_1 ? source2Pipe[351:344] : 8'h0)
    | (compressDataVec_hitReq_44_1 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_1 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_1 ? source2Pipe[375:368] : 8'h0)
    | (compressDataVec_hitReq_47_1 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_1 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_1 ? source2Pipe[399:392] : 8'h0)
    | (compressDataVec_hitReq_50_1 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_1 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_1 ? source2Pipe[423:416] : 8'h0)
    | (compressDataVec_hitReq_53_1 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_1 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_1 ? source2Pipe[447:440] : 8'h0)
    | (compressDataVec_hitReq_56_1 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_1 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_1 ? source2Pipe[471:464] : 8'h0)
    | (compressDataVec_hitReq_59_1 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_1 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_1 ? source2Pipe[495:488] : 8'h0)
    | (compressDataVec_hitReq_62_1 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_1 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_1;
  assign compressDataVec_useTail_1 = |(tailCount[5:1]);
  wire          _GEN_64 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h2;
  wire          compressDataVec_hitReq_0_2;
  assign compressDataVec_hitReq_0_2 = _GEN_64;
  wire          compressDataVec_hitReq_0_130;
  assign compressDataVec_hitReq_0_130 = _GEN_64;
  wire          compressDataVec_hitReq_0_194;
  assign compressDataVec_hitReq_0_194 = _GEN_64;
  wire          _GEN_65 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h2;
  wire          compressDataVec_hitReq_1_2;
  assign compressDataVec_hitReq_1_2 = _GEN_65;
  wire          compressDataVec_hitReq_1_130;
  assign compressDataVec_hitReq_1_130 = _GEN_65;
  wire          compressDataVec_hitReq_1_194;
  assign compressDataVec_hitReq_1_194 = _GEN_65;
  wire          _GEN_66 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h2;
  wire          compressDataVec_hitReq_2_2;
  assign compressDataVec_hitReq_2_2 = _GEN_66;
  wire          compressDataVec_hitReq_2_130;
  assign compressDataVec_hitReq_2_130 = _GEN_66;
  wire          compressDataVec_hitReq_2_194;
  assign compressDataVec_hitReq_2_194 = _GEN_66;
  wire          _GEN_67 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h2;
  wire          compressDataVec_hitReq_3_2;
  assign compressDataVec_hitReq_3_2 = _GEN_67;
  wire          compressDataVec_hitReq_3_130;
  assign compressDataVec_hitReq_3_130 = _GEN_67;
  wire          compressDataVec_hitReq_3_194;
  assign compressDataVec_hitReq_3_194 = _GEN_67;
  wire          _GEN_68 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h2;
  wire          compressDataVec_hitReq_4_2;
  assign compressDataVec_hitReq_4_2 = _GEN_68;
  wire          compressDataVec_hitReq_4_130;
  assign compressDataVec_hitReq_4_130 = _GEN_68;
  wire          compressDataVec_hitReq_4_194;
  assign compressDataVec_hitReq_4_194 = _GEN_68;
  wire          _GEN_69 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h2;
  wire          compressDataVec_hitReq_5_2;
  assign compressDataVec_hitReq_5_2 = _GEN_69;
  wire          compressDataVec_hitReq_5_130;
  assign compressDataVec_hitReq_5_130 = _GEN_69;
  wire          compressDataVec_hitReq_5_194;
  assign compressDataVec_hitReq_5_194 = _GEN_69;
  wire          _GEN_70 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h2;
  wire          compressDataVec_hitReq_6_2;
  assign compressDataVec_hitReq_6_2 = _GEN_70;
  wire          compressDataVec_hitReq_6_130;
  assign compressDataVec_hitReq_6_130 = _GEN_70;
  wire          compressDataVec_hitReq_6_194;
  assign compressDataVec_hitReq_6_194 = _GEN_70;
  wire          _GEN_71 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h2;
  wire          compressDataVec_hitReq_7_2;
  assign compressDataVec_hitReq_7_2 = _GEN_71;
  wire          compressDataVec_hitReq_7_130;
  assign compressDataVec_hitReq_7_130 = _GEN_71;
  wire          compressDataVec_hitReq_7_194;
  assign compressDataVec_hitReq_7_194 = _GEN_71;
  wire          _GEN_72 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h2;
  wire          compressDataVec_hitReq_8_2;
  assign compressDataVec_hitReq_8_2 = _GEN_72;
  wire          compressDataVec_hitReq_8_130;
  assign compressDataVec_hitReq_8_130 = _GEN_72;
  wire          compressDataVec_hitReq_8_194;
  assign compressDataVec_hitReq_8_194 = _GEN_72;
  wire          _GEN_73 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h2;
  wire          compressDataVec_hitReq_9_2;
  assign compressDataVec_hitReq_9_2 = _GEN_73;
  wire          compressDataVec_hitReq_9_130;
  assign compressDataVec_hitReq_9_130 = _GEN_73;
  wire          compressDataVec_hitReq_9_194;
  assign compressDataVec_hitReq_9_194 = _GEN_73;
  wire          _GEN_74 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h2;
  wire          compressDataVec_hitReq_10_2;
  assign compressDataVec_hitReq_10_2 = _GEN_74;
  wire          compressDataVec_hitReq_10_130;
  assign compressDataVec_hitReq_10_130 = _GEN_74;
  wire          compressDataVec_hitReq_10_194;
  assign compressDataVec_hitReq_10_194 = _GEN_74;
  wire          _GEN_75 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h2;
  wire          compressDataVec_hitReq_11_2;
  assign compressDataVec_hitReq_11_2 = _GEN_75;
  wire          compressDataVec_hitReq_11_130;
  assign compressDataVec_hitReq_11_130 = _GEN_75;
  wire          compressDataVec_hitReq_11_194;
  assign compressDataVec_hitReq_11_194 = _GEN_75;
  wire          _GEN_76 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h2;
  wire          compressDataVec_hitReq_12_2;
  assign compressDataVec_hitReq_12_2 = _GEN_76;
  wire          compressDataVec_hitReq_12_130;
  assign compressDataVec_hitReq_12_130 = _GEN_76;
  wire          compressDataVec_hitReq_12_194;
  assign compressDataVec_hitReq_12_194 = _GEN_76;
  wire          _GEN_77 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h2;
  wire          compressDataVec_hitReq_13_2;
  assign compressDataVec_hitReq_13_2 = _GEN_77;
  wire          compressDataVec_hitReq_13_130;
  assign compressDataVec_hitReq_13_130 = _GEN_77;
  wire          compressDataVec_hitReq_13_194;
  assign compressDataVec_hitReq_13_194 = _GEN_77;
  wire          _GEN_78 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h2;
  wire          compressDataVec_hitReq_14_2;
  assign compressDataVec_hitReq_14_2 = _GEN_78;
  wire          compressDataVec_hitReq_14_130;
  assign compressDataVec_hitReq_14_130 = _GEN_78;
  wire          compressDataVec_hitReq_14_194;
  assign compressDataVec_hitReq_14_194 = _GEN_78;
  wire          _GEN_79 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h2;
  wire          compressDataVec_hitReq_15_2;
  assign compressDataVec_hitReq_15_2 = _GEN_79;
  wire          compressDataVec_hitReq_15_130;
  assign compressDataVec_hitReq_15_130 = _GEN_79;
  wire          compressDataVec_hitReq_15_194;
  assign compressDataVec_hitReq_15_194 = _GEN_79;
  wire          _GEN_80 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h2;
  wire          compressDataVec_hitReq_16_2;
  assign compressDataVec_hitReq_16_2 = _GEN_80;
  wire          compressDataVec_hitReq_16_130;
  assign compressDataVec_hitReq_16_130 = _GEN_80;
  wire          _GEN_81 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h2;
  wire          compressDataVec_hitReq_17_2;
  assign compressDataVec_hitReq_17_2 = _GEN_81;
  wire          compressDataVec_hitReq_17_130;
  assign compressDataVec_hitReq_17_130 = _GEN_81;
  wire          _GEN_82 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h2;
  wire          compressDataVec_hitReq_18_2;
  assign compressDataVec_hitReq_18_2 = _GEN_82;
  wire          compressDataVec_hitReq_18_130;
  assign compressDataVec_hitReq_18_130 = _GEN_82;
  wire          _GEN_83 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h2;
  wire          compressDataVec_hitReq_19_2;
  assign compressDataVec_hitReq_19_2 = _GEN_83;
  wire          compressDataVec_hitReq_19_130;
  assign compressDataVec_hitReq_19_130 = _GEN_83;
  wire          _GEN_84 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h2;
  wire          compressDataVec_hitReq_20_2;
  assign compressDataVec_hitReq_20_2 = _GEN_84;
  wire          compressDataVec_hitReq_20_130;
  assign compressDataVec_hitReq_20_130 = _GEN_84;
  wire          _GEN_85 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h2;
  wire          compressDataVec_hitReq_21_2;
  assign compressDataVec_hitReq_21_2 = _GEN_85;
  wire          compressDataVec_hitReq_21_130;
  assign compressDataVec_hitReq_21_130 = _GEN_85;
  wire          _GEN_86 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h2;
  wire          compressDataVec_hitReq_22_2;
  assign compressDataVec_hitReq_22_2 = _GEN_86;
  wire          compressDataVec_hitReq_22_130;
  assign compressDataVec_hitReq_22_130 = _GEN_86;
  wire          _GEN_87 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h2;
  wire          compressDataVec_hitReq_23_2;
  assign compressDataVec_hitReq_23_2 = _GEN_87;
  wire          compressDataVec_hitReq_23_130;
  assign compressDataVec_hitReq_23_130 = _GEN_87;
  wire          _GEN_88 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h2;
  wire          compressDataVec_hitReq_24_2;
  assign compressDataVec_hitReq_24_2 = _GEN_88;
  wire          compressDataVec_hitReq_24_130;
  assign compressDataVec_hitReq_24_130 = _GEN_88;
  wire          _GEN_89 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h2;
  wire          compressDataVec_hitReq_25_2;
  assign compressDataVec_hitReq_25_2 = _GEN_89;
  wire          compressDataVec_hitReq_25_130;
  assign compressDataVec_hitReq_25_130 = _GEN_89;
  wire          _GEN_90 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h2;
  wire          compressDataVec_hitReq_26_2;
  assign compressDataVec_hitReq_26_2 = _GEN_90;
  wire          compressDataVec_hitReq_26_130;
  assign compressDataVec_hitReq_26_130 = _GEN_90;
  wire          _GEN_91 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h2;
  wire          compressDataVec_hitReq_27_2;
  assign compressDataVec_hitReq_27_2 = _GEN_91;
  wire          compressDataVec_hitReq_27_130;
  assign compressDataVec_hitReq_27_130 = _GEN_91;
  wire          _GEN_92 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h2;
  wire          compressDataVec_hitReq_28_2;
  assign compressDataVec_hitReq_28_2 = _GEN_92;
  wire          compressDataVec_hitReq_28_130;
  assign compressDataVec_hitReq_28_130 = _GEN_92;
  wire          _GEN_93 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h2;
  wire          compressDataVec_hitReq_29_2;
  assign compressDataVec_hitReq_29_2 = _GEN_93;
  wire          compressDataVec_hitReq_29_130;
  assign compressDataVec_hitReq_29_130 = _GEN_93;
  wire          _GEN_94 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h2;
  wire          compressDataVec_hitReq_30_2;
  assign compressDataVec_hitReq_30_2 = _GEN_94;
  wire          compressDataVec_hitReq_30_130;
  assign compressDataVec_hitReq_30_130 = _GEN_94;
  wire          _GEN_95 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h2;
  wire          compressDataVec_hitReq_31_2;
  assign compressDataVec_hitReq_31_2 = _GEN_95;
  wire          compressDataVec_hitReq_31_130;
  assign compressDataVec_hitReq_31_130 = _GEN_95;
  wire          compressDataVec_hitReq_32_2 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h2;
  wire          compressDataVec_hitReq_33_2 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h2;
  wire          compressDataVec_hitReq_34_2 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h2;
  wire          compressDataVec_hitReq_35_2 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h2;
  wire          compressDataVec_hitReq_36_2 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h2;
  wire          compressDataVec_hitReq_37_2 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h2;
  wire          compressDataVec_hitReq_38_2 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h2;
  wire          compressDataVec_hitReq_39_2 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h2;
  wire          compressDataVec_hitReq_40_2 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h2;
  wire          compressDataVec_hitReq_41_2 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h2;
  wire          compressDataVec_hitReq_42_2 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h2;
  wire          compressDataVec_hitReq_43_2 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h2;
  wire          compressDataVec_hitReq_44_2 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h2;
  wire          compressDataVec_hitReq_45_2 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h2;
  wire          compressDataVec_hitReq_46_2 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h2;
  wire          compressDataVec_hitReq_47_2 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h2;
  wire          compressDataVec_hitReq_48_2 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h2;
  wire          compressDataVec_hitReq_49_2 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h2;
  wire          compressDataVec_hitReq_50_2 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h2;
  wire          compressDataVec_hitReq_51_2 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h2;
  wire          compressDataVec_hitReq_52_2 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h2;
  wire          compressDataVec_hitReq_53_2 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h2;
  wire          compressDataVec_hitReq_54_2 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h2;
  wire          compressDataVec_hitReq_55_2 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h2;
  wire          compressDataVec_hitReq_56_2 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h2;
  wire          compressDataVec_hitReq_57_2 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h2;
  wire          compressDataVec_hitReq_58_2 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h2;
  wire          compressDataVec_hitReq_59_2 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h2;
  wire          compressDataVec_hitReq_60_2 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h2;
  wire          compressDataVec_hitReq_61_2 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h2;
  wire          compressDataVec_hitReq_62_2 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h2;
  wire          compressDataVec_hitReq_63_2 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h2;
  wire [7:0]    compressDataVec_selectReqData_2 =
    (compressDataVec_hitReq_0_2 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_2 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_2 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_2 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_2 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_2 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_2 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_2 ? source2Pipe[63:56] : 8'h0)
    | (compressDataVec_hitReq_8_2 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_2 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_2 ? source2Pipe[87:80] : 8'h0)
    | (compressDataVec_hitReq_11_2 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_2 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_2 ? source2Pipe[111:104] : 8'h0)
    | (compressDataVec_hitReq_14_2 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_2 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_2 ? source2Pipe[135:128] : 8'h0)
    | (compressDataVec_hitReq_17_2 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_2 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_2 ? source2Pipe[159:152] : 8'h0)
    | (compressDataVec_hitReq_20_2 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_2 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_2 ? source2Pipe[183:176] : 8'h0)
    | (compressDataVec_hitReq_23_2 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_2 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_2 ? source2Pipe[207:200] : 8'h0)
    | (compressDataVec_hitReq_26_2 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_2 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_2 ? source2Pipe[231:224] : 8'h0)
    | (compressDataVec_hitReq_29_2 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_2 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_2 ? source2Pipe[255:248] : 8'h0)
    | (compressDataVec_hitReq_32_2 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_2 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_2 ? source2Pipe[279:272] : 8'h0)
    | (compressDataVec_hitReq_35_2 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_2 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_2 ? source2Pipe[303:296] : 8'h0)
    | (compressDataVec_hitReq_38_2 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_2 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_2 ? source2Pipe[327:320] : 8'h0)
    | (compressDataVec_hitReq_41_2 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_2 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_2 ? source2Pipe[351:344] : 8'h0)
    | (compressDataVec_hitReq_44_2 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_2 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_2 ? source2Pipe[375:368] : 8'h0)
    | (compressDataVec_hitReq_47_2 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_2 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_2 ? source2Pipe[399:392] : 8'h0)
    | (compressDataVec_hitReq_50_2 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_2 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_2 ? source2Pipe[423:416] : 8'h0)
    | (compressDataVec_hitReq_53_2 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_2 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_2 ? source2Pipe[447:440] : 8'h0)
    | (compressDataVec_hitReq_56_2 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_2 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_2 ? source2Pipe[471:464] : 8'h0)
    | (compressDataVec_hitReq_59_2 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_2 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_2 ? source2Pipe[495:488] : 8'h0)
    | (compressDataVec_hitReq_62_2 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_2 ? source2Pipe[511:504] : 8'h0);
  wire          _GEN_96 = tailCount > 6'h2;
  wire          compressDataVec_useTail_2;
  assign compressDataVec_useTail_2 = _GEN_96;
  wire          compressDataVec_useTail_66;
  assign compressDataVec_useTail_66 = _GEN_96;
  wire          compressDataVec_useTail_98;
  assign compressDataVec_useTail_98 = _GEN_96;
  wire          _GEN_97 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h3;
  wire          compressDataVec_hitReq_0_3;
  assign compressDataVec_hitReq_0_3 = _GEN_97;
  wire          compressDataVec_hitReq_0_131;
  assign compressDataVec_hitReq_0_131 = _GEN_97;
  wire          compressDataVec_hitReq_0_195;
  assign compressDataVec_hitReq_0_195 = _GEN_97;
  wire          _GEN_98 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h3;
  wire          compressDataVec_hitReq_1_3;
  assign compressDataVec_hitReq_1_3 = _GEN_98;
  wire          compressDataVec_hitReq_1_131;
  assign compressDataVec_hitReq_1_131 = _GEN_98;
  wire          compressDataVec_hitReq_1_195;
  assign compressDataVec_hitReq_1_195 = _GEN_98;
  wire          _GEN_99 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h3;
  wire          compressDataVec_hitReq_2_3;
  assign compressDataVec_hitReq_2_3 = _GEN_99;
  wire          compressDataVec_hitReq_2_131;
  assign compressDataVec_hitReq_2_131 = _GEN_99;
  wire          compressDataVec_hitReq_2_195;
  assign compressDataVec_hitReq_2_195 = _GEN_99;
  wire          _GEN_100 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h3;
  wire          compressDataVec_hitReq_3_3;
  assign compressDataVec_hitReq_3_3 = _GEN_100;
  wire          compressDataVec_hitReq_3_131;
  assign compressDataVec_hitReq_3_131 = _GEN_100;
  wire          compressDataVec_hitReq_3_195;
  assign compressDataVec_hitReq_3_195 = _GEN_100;
  wire          _GEN_101 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h3;
  wire          compressDataVec_hitReq_4_3;
  assign compressDataVec_hitReq_4_3 = _GEN_101;
  wire          compressDataVec_hitReq_4_131;
  assign compressDataVec_hitReq_4_131 = _GEN_101;
  wire          compressDataVec_hitReq_4_195;
  assign compressDataVec_hitReq_4_195 = _GEN_101;
  wire          _GEN_102 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h3;
  wire          compressDataVec_hitReq_5_3;
  assign compressDataVec_hitReq_5_3 = _GEN_102;
  wire          compressDataVec_hitReq_5_131;
  assign compressDataVec_hitReq_5_131 = _GEN_102;
  wire          compressDataVec_hitReq_5_195;
  assign compressDataVec_hitReq_5_195 = _GEN_102;
  wire          _GEN_103 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h3;
  wire          compressDataVec_hitReq_6_3;
  assign compressDataVec_hitReq_6_3 = _GEN_103;
  wire          compressDataVec_hitReq_6_131;
  assign compressDataVec_hitReq_6_131 = _GEN_103;
  wire          compressDataVec_hitReq_6_195;
  assign compressDataVec_hitReq_6_195 = _GEN_103;
  wire          _GEN_104 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h3;
  wire          compressDataVec_hitReq_7_3;
  assign compressDataVec_hitReq_7_3 = _GEN_104;
  wire          compressDataVec_hitReq_7_131;
  assign compressDataVec_hitReq_7_131 = _GEN_104;
  wire          compressDataVec_hitReq_7_195;
  assign compressDataVec_hitReq_7_195 = _GEN_104;
  wire          _GEN_105 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h3;
  wire          compressDataVec_hitReq_8_3;
  assign compressDataVec_hitReq_8_3 = _GEN_105;
  wire          compressDataVec_hitReq_8_131;
  assign compressDataVec_hitReq_8_131 = _GEN_105;
  wire          compressDataVec_hitReq_8_195;
  assign compressDataVec_hitReq_8_195 = _GEN_105;
  wire          _GEN_106 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h3;
  wire          compressDataVec_hitReq_9_3;
  assign compressDataVec_hitReq_9_3 = _GEN_106;
  wire          compressDataVec_hitReq_9_131;
  assign compressDataVec_hitReq_9_131 = _GEN_106;
  wire          compressDataVec_hitReq_9_195;
  assign compressDataVec_hitReq_9_195 = _GEN_106;
  wire          _GEN_107 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h3;
  wire          compressDataVec_hitReq_10_3;
  assign compressDataVec_hitReq_10_3 = _GEN_107;
  wire          compressDataVec_hitReq_10_131;
  assign compressDataVec_hitReq_10_131 = _GEN_107;
  wire          compressDataVec_hitReq_10_195;
  assign compressDataVec_hitReq_10_195 = _GEN_107;
  wire          _GEN_108 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h3;
  wire          compressDataVec_hitReq_11_3;
  assign compressDataVec_hitReq_11_3 = _GEN_108;
  wire          compressDataVec_hitReq_11_131;
  assign compressDataVec_hitReq_11_131 = _GEN_108;
  wire          compressDataVec_hitReq_11_195;
  assign compressDataVec_hitReq_11_195 = _GEN_108;
  wire          _GEN_109 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h3;
  wire          compressDataVec_hitReq_12_3;
  assign compressDataVec_hitReq_12_3 = _GEN_109;
  wire          compressDataVec_hitReq_12_131;
  assign compressDataVec_hitReq_12_131 = _GEN_109;
  wire          compressDataVec_hitReq_12_195;
  assign compressDataVec_hitReq_12_195 = _GEN_109;
  wire          _GEN_110 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h3;
  wire          compressDataVec_hitReq_13_3;
  assign compressDataVec_hitReq_13_3 = _GEN_110;
  wire          compressDataVec_hitReq_13_131;
  assign compressDataVec_hitReq_13_131 = _GEN_110;
  wire          compressDataVec_hitReq_13_195;
  assign compressDataVec_hitReq_13_195 = _GEN_110;
  wire          _GEN_111 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h3;
  wire          compressDataVec_hitReq_14_3;
  assign compressDataVec_hitReq_14_3 = _GEN_111;
  wire          compressDataVec_hitReq_14_131;
  assign compressDataVec_hitReq_14_131 = _GEN_111;
  wire          compressDataVec_hitReq_14_195;
  assign compressDataVec_hitReq_14_195 = _GEN_111;
  wire          _GEN_112 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h3;
  wire          compressDataVec_hitReq_15_3;
  assign compressDataVec_hitReq_15_3 = _GEN_112;
  wire          compressDataVec_hitReq_15_131;
  assign compressDataVec_hitReq_15_131 = _GEN_112;
  wire          compressDataVec_hitReq_15_195;
  assign compressDataVec_hitReq_15_195 = _GEN_112;
  wire          _GEN_113 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h3;
  wire          compressDataVec_hitReq_16_3;
  assign compressDataVec_hitReq_16_3 = _GEN_113;
  wire          compressDataVec_hitReq_16_131;
  assign compressDataVec_hitReq_16_131 = _GEN_113;
  wire          _GEN_114 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h3;
  wire          compressDataVec_hitReq_17_3;
  assign compressDataVec_hitReq_17_3 = _GEN_114;
  wire          compressDataVec_hitReq_17_131;
  assign compressDataVec_hitReq_17_131 = _GEN_114;
  wire          _GEN_115 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h3;
  wire          compressDataVec_hitReq_18_3;
  assign compressDataVec_hitReq_18_3 = _GEN_115;
  wire          compressDataVec_hitReq_18_131;
  assign compressDataVec_hitReq_18_131 = _GEN_115;
  wire          _GEN_116 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h3;
  wire          compressDataVec_hitReq_19_3;
  assign compressDataVec_hitReq_19_3 = _GEN_116;
  wire          compressDataVec_hitReq_19_131;
  assign compressDataVec_hitReq_19_131 = _GEN_116;
  wire          _GEN_117 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h3;
  wire          compressDataVec_hitReq_20_3;
  assign compressDataVec_hitReq_20_3 = _GEN_117;
  wire          compressDataVec_hitReq_20_131;
  assign compressDataVec_hitReq_20_131 = _GEN_117;
  wire          _GEN_118 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h3;
  wire          compressDataVec_hitReq_21_3;
  assign compressDataVec_hitReq_21_3 = _GEN_118;
  wire          compressDataVec_hitReq_21_131;
  assign compressDataVec_hitReq_21_131 = _GEN_118;
  wire          _GEN_119 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h3;
  wire          compressDataVec_hitReq_22_3;
  assign compressDataVec_hitReq_22_3 = _GEN_119;
  wire          compressDataVec_hitReq_22_131;
  assign compressDataVec_hitReq_22_131 = _GEN_119;
  wire          _GEN_120 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h3;
  wire          compressDataVec_hitReq_23_3;
  assign compressDataVec_hitReq_23_3 = _GEN_120;
  wire          compressDataVec_hitReq_23_131;
  assign compressDataVec_hitReq_23_131 = _GEN_120;
  wire          _GEN_121 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h3;
  wire          compressDataVec_hitReq_24_3;
  assign compressDataVec_hitReq_24_3 = _GEN_121;
  wire          compressDataVec_hitReq_24_131;
  assign compressDataVec_hitReq_24_131 = _GEN_121;
  wire          _GEN_122 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h3;
  wire          compressDataVec_hitReq_25_3;
  assign compressDataVec_hitReq_25_3 = _GEN_122;
  wire          compressDataVec_hitReq_25_131;
  assign compressDataVec_hitReq_25_131 = _GEN_122;
  wire          _GEN_123 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h3;
  wire          compressDataVec_hitReq_26_3;
  assign compressDataVec_hitReq_26_3 = _GEN_123;
  wire          compressDataVec_hitReq_26_131;
  assign compressDataVec_hitReq_26_131 = _GEN_123;
  wire          _GEN_124 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h3;
  wire          compressDataVec_hitReq_27_3;
  assign compressDataVec_hitReq_27_3 = _GEN_124;
  wire          compressDataVec_hitReq_27_131;
  assign compressDataVec_hitReq_27_131 = _GEN_124;
  wire          _GEN_125 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h3;
  wire          compressDataVec_hitReq_28_3;
  assign compressDataVec_hitReq_28_3 = _GEN_125;
  wire          compressDataVec_hitReq_28_131;
  assign compressDataVec_hitReq_28_131 = _GEN_125;
  wire          _GEN_126 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h3;
  wire          compressDataVec_hitReq_29_3;
  assign compressDataVec_hitReq_29_3 = _GEN_126;
  wire          compressDataVec_hitReq_29_131;
  assign compressDataVec_hitReq_29_131 = _GEN_126;
  wire          _GEN_127 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h3;
  wire          compressDataVec_hitReq_30_3;
  assign compressDataVec_hitReq_30_3 = _GEN_127;
  wire          compressDataVec_hitReq_30_131;
  assign compressDataVec_hitReq_30_131 = _GEN_127;
  wire          _GEN_128 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h3;
  wire          compressDataVec_hitReq_31_3;
  assign compressDataVec_hitReq_31_3 = _GEN_128;
  wire          compressDataVec_hitReq_31_131;
  assign compressDataVec_hitReq_31_131 = _GEN_128;
  wire          compressDataVec_hitReq_32_3 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h3;
  wire          compressDataVec_hitReq_33_3 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h3;
  wire          compressDataVec_hitReq_34_3 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h3;
  wire          compressDataVec_hitReq_35_3 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h3;
  wire          compressDataVec_hitReq_36_3 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h3;
  wire          compressDataVec_hitReq_37_3 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h3;
  wire          compressDataVec_hitReq_38_3 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h3;
  wire          compressDataVec_hitReq_39_3 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h3;
  wire          compressDataVec_hitReq_40_3 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h3;
  wire          compressDataVec_hitReq_41_3 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h3;
  wire          compressDataVec_hitReq_42_3 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h3;
  wire          compressDataVec_hitReq_43_3 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h3;
  wire          compressDataVec_hitReq_44_3 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h3;
  wire          compressDataVec_hitReq_45_3 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h3;
  wire          compressDataVec_hitReq_46_3 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h3;
  wire          compressDataVec_hitReq_47_3 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h3;
  wire          compressDataVec_hitReq_48_3 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h3;
  wire          compressDataVec_hitReq_49_3 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h3;
  wire          compressDataVec_hitReq_50_3 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h3;
  wire          compressDataVec_hitReq_51_3 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h3;
  wire          compressDataVec_hitReq_52_3 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h3;
  wire          compressDataVec_hitReq_53_3 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h3;
  wire          compressDataVec_hitReq_54_3 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h3;
  wire          compressDataVec_hitReq_55_3 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h3;
  wire          compressDataVec_hitReq_56_3 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h3;
  wire          compressDataVec_hitReq_57_3 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h3;
  wire          compressDataVec_hitReq_58_3 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h3;
  wire          compressDataVec_hitReq_59_3 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h3;
  wire          compressDataVec_hitReq_60_3 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h3;
  wire          compressDataVec_hitReq_61_3 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h3;
  wire          compressDataVec_hitReq_62_3 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h3;
  wire          compressDataVec_hitReq_63_3 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h3;
  wire [7:0]    compressDataVec_selectReqData_3 =
    (compressDataVec_hitReq_0_3 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_3 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_3 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_3 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_3 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_3 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_3 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_3 ? source2Pipe[63:56] : 8'h0)
    | (compressDataVec_hitReq_8_3 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_3 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_3 ? source2Pipe[87:80] : 8'h0)
    | (compressDataVec_hitReq_11_3 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_3 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_3 ? source2Pipe[111:104] : 8'h0)
    | (compressDataVec_hitReq_14_3 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_3 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_3 ? source2Pipe[135:128] : 8'h0)
    | (compressDataVec_hitReq_17_3 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_3 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_3 ? source2Pipe[159:152] : 8'h0)
    | (compressDataVec_hitReq_20_3 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_3 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_3 ? source2Pipe[183:176] : 8'h0)
    | (compressDataVec_hitReq_23_3 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_3 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_3 ? source2Pipe[207:200] : 8'h0)
    | (compressDataVec_hitReq_26_3 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_3 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_3 ? source2Pipe[231:224] : 8'h0)
    | (compressDataVec_hitReq_29_3 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_3 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_3 ? source2Pipe[255:248] : 8'h0)
    | (compressDataVec_hitReq_32_3 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_3 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_3 ? source2Pipe[279:272] : 8'h0)
    | (compressDataVec_hitReq_35_3 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_3 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_3 ? source2Pipe[303:296] : 8'h0)
    | (compressDataVec_hitReq_38_3 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_3 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_3 ? source2Pipe[327:320] : 8'h0)
    | (compressDataVec_hitReq_41_3 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_3 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_3 ? source2Pipe[351:344] : 8'h0)
    | (compressDataVec_hitReq_44_3 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_3 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_3 ? source2Pipe[375:368] : 8'h0)
    | (compressDataVec_hitReq_47_3 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_3 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_3 ? source2Pipe[399:392] : 8'h0)
    | (compressDataVec_hitReq_50_3 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_3 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_3 ? source2Pipe[423:416] : 8'h0)
    | (compressDataVec_hitReq_53_3 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_3 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_3 ? source2Pipe[447:440] : 8'h0)
    | (compressDataVec_hitReq_56_3 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_3 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_3 ? source2Pipe[471:464] : 8'h0)
    | (compressDataVec_hitReq_59_3 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_3 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_3 ? source2Pipe[495:488] : 8'h0)
    | (compressDataVec_hitReq_62_3 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_3 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_3;
  assign compressDataVec_useTail_3 = |(tailCount[5:2]);
  wire          _GEN_129 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h4;
  wire          compressDataVec_hitReq_0_4;
  assign compressDataVec_hitReq_0_4 = _GEN_129;
  wire          compressDataVec_hitReq_0_132;
  assign compressDataVec_hitReq_0_132 = _GEN_129;
  wire          compressDataVec_hitReq_0_196;
  assign compressDataVec_hitReq_0_196 = _GEN_129;
  wire          _GEN_130 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h4;
  wire          compressDataVec_hitReq_1_4;
  assign compressDataVec_hitReq_1_4 = _GEN_130;
  wire          compressDataVec_hitReq_1_132;
  assign compressDataVec_hitReq_1_132 = _GEN_130;
  wire          compressDataVec_hitReq_1_196;
  assign compressDataVec_hitReq_1_196 = _GEN_130;
  wire          _GEN_131 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h4;
  wire          compressDataVec_hitReq_2_4;
  assign compressDataVec_hitReq_2_4 = _GEN_131;
  wire          compressDataVec_hitReq_2_132;
  assign compressDataVec_hitReq_2_132 = _GEN_131;
  wire          compressDataVec_hitReq_2_196;
  assign compressDataVec_hitReq_2_196 = _GEN_131;
  wire          _GEN_132 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h4;
  wire          compressDataVec_hitReq_3_4;
  assign compressDataVec_hitReq_3_4 = _GEN_132;
  wire          compressDataVec_hitReq_3_132;
  assign compressDataVec_hitReq_3_132 = _GEN_132;
  wire          compressDataVec_hitReq_3_196;
  assign compressDataVec_hitReq_3_196 = _GEN_132;
  wire          _GEN_133 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h4;
  wire          compressDataVec_hitReq_4_4;
  assign compressDataVec_hitReq_4_4 = _GEN_133;
  wire          compressDataVec_hitReq_4_132;
  assign compressDataVec_hitReq_4_132 = _GEN_133;
  wire          compressDataVec_hitReq_4_196;
  assign compressDataVec_hitReq_4_196 = _GEN_133;
  wire          _GEN_134 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h4;
  wire          compressDataVec_hitReq_5_4;
  assign compressDataVec_hitReq_5_4 = _GEN_134;
  wire          compressDataVec_hitReq_5_132;
  assign compressDataVec_hitReq_5_132 = _GEN_134;
  wire          compressDataVec_hitReq_5_196;
  assign compressDataVec_hitReq_5_196 = _GEN_134;
  wire          _GEN_135 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h4;
  wire          compressDataVec_hitReq_6_4;
  assign compressDataVec_hitReq_6_4 = _GEN_135;
  wire          compressDataVec_hitReq_6_132;
  assign compressDataVec_hitReq_6_132 = _GEN_135;
  wire          compressDataVec_hitReq_6_196;
  assign compressDataVec_hitReq_6_196 = _GEN_135;
  wire          _GEN_136 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h4;
  wire          compressDataVec_hitReq_7_4;
  assign compressDataVec_hitReq_7_4 = _GEN_136;
  wire          compressDataVec_hitReq_7_132;
  assign compressDataVec_hitReq_7_132 = _GEN_136;
  wire          compressDataVec_hitReq_7_196;
  assign compressDataVec_hitReq_7_196 = _GEN_136;
  wire          _GEN_137 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h4;
  wire          compressDataVec_hitReq_8_4;
  assign compressDataVec_hitReq_8_4 = _GEN_137;
  wire          compressDataVec_hitReq_8_132;
  assign compressDataVec_hitReq_8_132 = _GEN_137;
  wire          compressDataVec_hitReq_8_196;
  assign compressDataVec_hitReq_8_196 = _GEN_137;
  wire          _GEN_138 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h4;
  wire          compressDataVec_hitReq_9_4;
  assign compressDataVec_hitReq_9_4 = _GEN_138;
  wire          compressDataVec_hitReq_9_132;
  assign compressDataVec_hitReq_9_132 = _GEN_138;
  wire          compressDataVec_hitReq_9_196;
  assign compressDataVec_hitReq_9_196 = _GEN_138;
  wire          _GEN_139 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h4;
  wire          compressDataVec_hitReq_10_4;
  assign compressDataVec_hitReq_10_4 = _GEN_139;
  wire          compressDataVec_hitReq_10_132;
  assign compressDataVec_hitReq_10_132 = _GEN_139;
  wire          compressDataVec_hitReq_10_196;
  assign compressDataVec_hitReq_10_196 = _GEN_139;
  wire          _GEN_140 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h4;
  wire          compressDataVec_hitReq_11_4;
  assign compressDataVec_hitReq_11_4 = _GEN_140;
  wire          compressDataVec_hitReq_11_132;
  assign compressDataVec_hitReq_11_132 = _GEN_140;
  wire          compressDataVec_hitReq_11_196;
  assign compressDataVec_hitReq_11_196 = _GEN_140;
  wire          _GEN_141 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h4;
  wire          compressDataVec_hitReq_12_4;
  assign compressDataVec_hitReq_12_4 = _GEN_141;
  wire          compressDataVec_hitReq_12_132;
  assign compressDataVec_hitReq_12_132 = _GEN_141;
  wire          compressDataVec_hitReq_12_196;
  assign compressDataVec_hitReq_12_196 = _GEN_141;
  wire          _GEN_142 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h4;
  wire          compressDataVec_hitReq_13_4;
  assign compressDataVec_hitReq_13_4 = _GEN_142;
  wire          compressDataVec_hitReq_13_132;
  assign compressDataVec_hitReq_13_132 = _GEN_142;
  wire          compressDataVec_hitReq_13_196;
  assign compressDataVec_hitReq_13_196 = _GEN_142;
  wire          _GEN_143 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h4;
  wire          compressDataVec_hitReq_14_4;
  assign compressDataVec_hitReq_14_4 = _GEN_143;
  wire          compressDataVec_hitReq_14_132;
  assign compressDataVec_hitReq_14_132 = _GEN_143;
  wire          compressDataVec_hitReq_14_196;
  assign compressDataVec_hitReq_14_196 = _GEN_143;
  wire          _GEN_144 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h4;
  wire          compressDataVec_hitReq_15_4;
  assign compressDataVec_hitReq_15_4 = _GEN_144;
  wire          compressDataVec_hitReq_15_132;
  assign compressDataVec_hitReq_15_132 = _GEN_144;
  wire          compressDataVec_hitReq_15_196;
  assign compressDataVec_hitReq_15_196 = _GEN_144;
  wire          _GEN_145 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h4;
  wire          compressDataVec_hitReq_16_4;
  assign compressDataVec_hitReq_16_4 = _GEN_145;
  wire          compressDataVec_hitReq_16_132;
  assign compressDataVec_hitReq_16_132 = _GEN_145;
  wire          _GEN_146 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h4;
  wire          compressDataVec_hitReq_17_4;
  assign compressDataVec_hitReq_17_4 = _GEN_146;
  wire          compressDataVec_hitReq_17_132;
  assign compressDataVec_hitReq_17_132 = _GEN_146;
  wire          _GEN_147 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h4;
  wire          compressDataVec_hitReq_18_4;
  assign compressDataVec_hitReq_18_4 = _GEN_147;
  wire          compressDataVec_hitReq_18_132;
  assign compressDataVec_hitReq_18_132 = _GEN_147;
  wire          _GEN_148 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h4;
  wire          compressDataVec_hitReq_19_4;
  assign compressDataVec_hitReq_19_4 = _GEN_148;
  wire          compressDataVec_hitReq_19_132;
  assign compressDataVec_hitReq_19_132 = _GEN_148;
  wire          _GEN_149 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h4;
  wire          compressDataVec_hitReq_20_4;
  assign compressDataVec_hitReq_20_4 = _GEN_149;
  wire          compressDataVec_hitReq_20_132;
  assign compressDataVec_hitReq_20_132 = _GEN_149;
  wire          _GEN_150 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h4;
  wire          compressDataVec_hitReq_21_4;
  assign compressDataVec_hitReq_21_4 = _GEN_150;
  wire          compressDataVec_hitReq_21_132;
  assign compressDataVec_hitReq_21_132 = _GEN_150;
  wire          _GEN_151 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h4;
  wire          compressDataVec_hitReq_22_4;
  assign compressDataVec_hitReq_22_4 = _GEN_151;
  wire          compressDataVec_hitReq_22_132;
  assign compressDataVec_hitReq_22_132 = _GEN_151;
  wire          _GEN_152 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h4;
  wire          compressDataVec_hitReq_23_4;
  assign compressDataVec_hitReq_23_4 = _GEN_152;
  wire          compressDataVec_hitReq_23_132;
  assign compressDataVec_hitReq_23_132 = _GEN_152;
  wire          _GEN_153 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h4;
  wire          compressDataVec_hitReq_24_4;
  assign compressDataVec_hitReq_24_4 = _GEN_153;
  wire          compressDataVec_hitReq_24_132;
  assign compressDataVec_hitReq_24_132 = _GEN_153;
  wire          _GEN_154 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h4;
  wire          compressDataVec_hitReq_25_4;
  assign compressDataVec_hitReq_25_4 = _GEN_154;
  wire          compressDataVec_hitReq_25_132;
  assign compressDataVec_hitReq_25_132 = _GEN_154;
  wire          _GEN_155 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h4;
  wire          compressDataVec_hitReq_26_4;
  assign compressDataVec_hitReq_26_4 = _GEN_155;
  wire          compressDataVec_hitReq_26_132;
  assign compressDataVec_hitReq_26_132 = _GEN_155;
  wire          _GEN_156 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h4;
  wire          compressDataVec_hitReq_27_4;
  assign compressDataVec_hitReq_27_4 = _GEN_156;
  wire          compressDataVec_hitReq_27_132;
  assign compressDataVec_hitReq_27_132 = _GEN_156;
  wire          _GEN_157 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h4;
  wire          compressDataVec_hitReq_28_4;
  assign compressDataVec_hitReq_28_4 = _GEN_157;
  wire          compressDataVec_hitReq_28_132;
  assign compressDataVec_hitReq_28_132 = _GEN_157;
  wire          _GEN_158 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h4;
  wire          compressDataVec_hitReq_29_4;
  assign compressDataVec_hitReq_29_4 = _GEN_158;
  wire          compressDataVec_hitReq_29_132;
  assign compressDataVec_hitReq_29_132 = _GEN_158;
  wire          _GEN_159 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h4;
  wire          compressDataVec_hitReq_30_4;
  assign compressDataVec_hitReq_30_4 = _GEN_159;
  wire          compressDataVec_hitReq_30_132;
  assign compressDataVec_hitReq_30_132 = _GEN_159;
  wire          _GEN_160 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h4;
  wire          compressDataVec_hitReq_31_4;
  assign compressDataVec_hitReq_31_4 = _GEN_160;
  wire          compressDataVec_hitReq_31_132;
  assign compressDataVec_hitReq_31_132 = _GEN_160;
  wire          compressDataVec_hitReq_32_4 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h4;
  wire          compressDataVec_hitReq_33_4 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h4;
  wire          compressDataVec_hitReq_34_4 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h4;
  wire          compressDataVec_hitReq_35_4 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h4;
  wire          compressDataVec_hitReq_36_4 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h4;
  wire          compressDataVec_hitReq_37_4 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h4;
  wire          compressDataVec_hitReq_38_4 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h4;
  wire          compressDataVec_hitReq_39_4 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h4;
  wire          compressDataVec_hitReq_40_4 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h4;
  wire          compressDataVec_hitReq_41_4 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h4;
  wire          compressDataVec_hitReq_42_4 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h4;
  wire          compressDataVec_hitReq_43_4 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h4;
  wire          compressDataVec_hitReq_44_4 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h4;
  wire          compressDataVec_hitReq_45_4 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h4;
  wire          compressDataVec_hitReq_46_4 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h4;
  wire          compressDataVec_hitReq_47_4 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h4;
  wire          compressDataVec_hitReq_48_4 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h4;
  wire          compressDataVec_hitReq_49_4 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h4;
  wire          compressDataVec_hitReq_50_4 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h4;
  wire          compressDataVec_hitReq_51_4 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h4;
  wire          compressDataVec_hitReq_52_4 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h4;
  wire          compressDataVec_hitReq_53_4 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h4;
  wire          compressDataVec_hitReq_54_4 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h4;
  wire          compressDataVec_hitReq_55_4 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h4;
  wire          compressDataVec_hitReq_56_4 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h4;
  wire          compressDataVec_hitReq_57_4 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h4;
  wire          compressDataVec_hitReq_58_4 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h4;
  wire          compressDataVec_hitReq_59_4 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h4;
  wire          compressDataVec_hitReq_60_4 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h4;
  wire          compressDataVec_hitReq_61_4 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h4;
  wire          compressDataVec_hitReq_62_4 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h4;
  wire          compressDataVec_hitReq_63_4 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h4;
  wire [7:0]    compressDataVec_selectReqData_4 =
    (compressDataVec_hitReq_0_4 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_4 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_4 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_4 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_4 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_4 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_4 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_4 ? source2Pipe[63:56] : 8'h0)
    | (compressDataVec_hitReq_8_4 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_4 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_4 ? source2Pipe[87:80] : 8'h0)
    | (compressDataVec_hitReq_11_4 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_4 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_4 ? source2Pipe[111:104] : 8'h0)
    | (compressDataVec_hitReq_14_4 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_4 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_4 ? source2Pipe[135:128] : 8'h0)
    | (compressDataVec_hitReq_17_4 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_4 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_4 ? source2Pipe[159:152] : 8'h0)
    | (compressDataVec_hitReq_20_4 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_4 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_4 ? source2Pipe[183:176] : 8'h0)
    | (compressDataVec_hitReq_23_4 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_4 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_4 ? source2Pipe[207:200] : 8'h0)
    | (compressDataVec_hitReq_26_4 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_4 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_4 ? source2Pipe[231:224] : 8'h0)
    | (compressDataVec_hitReq_29_4 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_4 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_4 ? source2Pipe[255:248] : 8'h0)
    | (compressDataVec_hitReq_32_4 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_4 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_4 ? source2Pipe[279:272] : 8'h0)
    | (compressDataVec_hitReq_35_4 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_4 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_4 ? source2Pipe[303:296] : 8'h0)
    | (compressDataVec_hitReq_38_4 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_4 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_4 ? source2Pipe[327:320] : 8'h0)
    | (compressDataVec_hitReq_41_4 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_4 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_4 ? source2Pipe[351:344] : 8'h0)
    | (compressDataVec_hitReq_44_4 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_4 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_4 ? source2Pipe[375:368] : 8'h0)
    | (compressDataVec_hitReq_47_4 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_4 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_4 ? source2Pipe[399:392] : 8'h0)
    | (compressDataVec_hitReq_50_4 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_4 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_4 ? source2Pipe[423:416] : 8'h0)
    | (compressDataVec_hitReq_53_4 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_4 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_4 ? source2Pipe[447:440] : 8'h0)
    | (compressDataVec_hitReq_56_4 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_4 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_4 ? source2Pipe[471:464] : 8'h0)
    | (compressDataVec_hitReq_59_4 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_4 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_4 ? source2Pipe[495:488] : 8'h0)
    | (compressDataVec_hitReq_62_4 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_4 ? source2Pipe[511:504] : 8'h0);
  wire          _GEN_161 = tailCount > 6'h4;
  wire          compressDataVec_useTail_4;
  assign compressDataVec_useTail_4 = _GEN_161;
  wire          compressDataVec_useTail_68;
  assign compressDataVec_useTail_68 = _GEN_161;
  wire          compressDataVec_useTail_100;
  assign compressDataVec_useTail_100 = _GEN_161;
  wire          _GEN_162 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h5;
  wire          compressDataVec_hitReq_0_5;
  assign compressDataVec_hitReq_0_5 = _GEN_162;
  wire          compressDataVec_hitReq_0_133;
  assign compressDataVec_hitReq_0_133 = _GEN_162;
  wire          compressDataVec_hitReq_0_197;
  assign compressDataVec_hitReq_0_197 = _GEN_162;
  wire          _GEN_163 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h5;
  wire          compressDataVec_hitReq_1_5;
  assign compressDataVec_hitReq_1_5 = _GEN_163;
  wire          compressDataVec_hitReq_1_133;
  assign compressDataVec_hitReq_1_133 = _GEN_163;
  wire          compressDataVec_hitReq_1_197;
  assign compressDataVec_hitReq_1_197 = _GEN_163;
  wire          _GEN_164 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h5;
  wire          compressDataVec_hitReq_2_5;
  assign compressDataVec_hitReq_2_5 = _GEN_164;
  wire          compressDataVec_hitReq_2_133;
  assign compressDataVec_hitReq_2_133 = _GEN_164;
  wire          compressDataVec_hitReq_2_197;
  assign compressDataVec_hitReq_2_197 = _GEN_164;
  wire          _GEN_165 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h5;
  wire          compressDataVec_hitReq_3_5;
  assign compressDataVec_hitReq_3_5 = _GEN_165;
  wire          compressDataVec_hitReq_3_133;
  assign compressDataVec_hitReq_3_133 = _GEN_165;
  wire          compressDataVec_hitReq_3_197;
  assign compressDataVec_hitReq_3_197 = _GEN_165;
  wire          _GEN_166 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h5;
  wire          compressDataVec_hitReq_4_5;
  assign compressDataVec_hitReq_4_5 = _GEN_166;
  wire          compressDataVec_hitReq_4_133;
  assign compressDataVec_hitReq_4_133 = _GEN_166;
  wire          compressDataVec_hitReq_4_197;
  assign compressDataVec_hitReq_4_197 = _GEN_166;
  wire          _GEN_167 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h5;
  wire          compressDataVec_hitReq_5_5;
  assign compressDataVec_hitReq_5_5 = _GEN_167;
  wire          compressDataVec_hitReq_5_133;
  assign compressDataVec_hitReq_5_133 = _GEN_167;
  wire          compressDataVec_hitReq_5_197;
  assign compressDataVec_hitReq_5_197 = _GEN_167;
  wire          _GEN_168 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h5;
  wire          compressDataVec_hitReq_6_5;
  assign compressDataVec_hitReq_6_5 = _GEN_168;
  wire          compressDataVec_hitReq_6_133;
  assign compressDataVec_hitReq_6_133 = _GEN_168;
  wire          compressDataVec_hitReq_6_197;
  assign compressDataVec_hitReq_6_197 = _GEN_168;
  wire          _GEN_169 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h5;
  wire          compressDataVec_hitReq_7_5;
  assign compressDataVec_hitReq_7_5 = _GEN_169;
  wire          compressDataVec_hitReq_7_133;
  assign compressDataVec_hitReq_7_133 = _GEN_169;
  wire          compressDataVec_hitReq_7_197;
  assign compressDataVec_hitReq_7_197 = _GEN_169;
  wire          _GEN_170 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h5;
  wire          compressDataVec_hitReq_8_5;
  assign compressDataVec_hitReq_8_5 = _GEN_170;
  wire          compressDataVec_hitReq_8_133;
  assign compressDataVec_hitReq_8_133 = _GEN_170;
  wire          compressDataVec_hitReq_8_197;
  assign compressDataVec_hitReq_8_197 = _GEN_170;
  wire          _GEN_171 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h5;
  wire          compressDataVec_hitReq_9_5;
  assign compressDataVec_hitReq_9_5 = _GEN_171;
  wire          compressDataVec_hitReq_9_133;
  assign compressDataVec_hitReq_9_133 = _GEN_171;
  wire          compressDataVec_hitReq_9_197;
  assign compressDataVec_hitReq_9_197 = _GEN_171;
  wire          _GEN_172 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h5;
  wire          compressDataVec_hitReq_10_5;
  assign compressDataVec_hitReq_10_5 = _GEN_172;
  wire          compressDataVec_hitReq_10_133;
  assign compressDataVec_hitReq_10_133 = _GEN_172;
  wire          compressDataVec_hitReq_10_197;
  assign compressDataVec_hitReq_10_197 = _GEN_172;
  wire          _GEN_173 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h5;
  wire          compressDataVec_hitReq_11_5;
  assign compressDataVec_hitReq_11_5 = _GEN_173;
  wire          compressDataVec_hitReq_11_133;
  assign compressDataVec_hitReq_11_133 = _GEN_173;
  wire          compressDataVec_hitReq_11_197;
  assign compressDataVec_hitReq_11_197 = _GEN_173;
  wire          _GEN_174 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h5;
  wire          compressDataVec_hitReq_12_5;
  assign compressDataVec_hitReq_12_5 = _GEN_174;
  wire          compressDataVec_hitReq_12_133;
  assign compressDataVec_hitReq_12_133 = _GEN_174;
  wire          compressDataVec_hitReq_12_197;
  assign compressDataVec_hitReq_12_197 = _GEN_174;
  wire          _GEN_175 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h5;
  wire          compressDataVec_hitReq_13_5;
  assign compressDataVec_hitReq_13_5 = _GEN_175;
  wire          compressDataVec_hitReq_13_133;
  assign compressDataVec_hitReq_13_133 = _GEN_175;
  wire          compressDataVec_hitReq_13_197;
  assign compressDataVec_hitReq_13_197 = _GEN_175;
  wire          _GEN_176 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h5;
  wire          compressDataVec_hitReq_14_5;
  assign compressDataVec_hitReq_14_5 = _GEN_176;
  wire          compressDataVec_hitReq_14_133;
  assign compressDataVec_hitReq_14_133 = _GEN_176;
  wire          compressDataVec_hitReq_14_197;
  assign compressDataVec_hitReq_14_197 = _GEN_176;
  wire          _GEN_177 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h5;
  wire          compressDataVec_hitReq_15_5;
  assign compressDataVec_hitReq_15_5 = _GEN_177;
  wire          compressDataVec_hitReq_15_133;
  assign compressDataVec_hitReq_15_133 = _GEN_177;
  wire          compressDataVec_hitReq_15_197;
  assign compressDataVec_hitReq_15_197 = _GEN_177;
  wire          _GEN_178 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h5;
  wire          compressDataVec_hitReq_16_5;
  assign compressDataVec_hitReq_16_5 = _GEN_178;
  wire          compressDataVec_hitReq_16_133;
  assign compressDataVec_hitReq_16_133 = _GEN_178;
  wire          _GEN_179 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h5;
  wire          compressDataVec_hitReq_17_5;
  assign compressDataVec_hitReq_17_5 = _GEN_179;
  wire          compressDataVec_hitReq_17_133;
  assign compressDataVec_hitReq_17_133 = _GEN_179;
  wire          _GEN_180 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h5;
  wire          compressDataVec_hitReq_18_5;
  assign compressDataVec_hitReq_18_5 = _GEN_180;
  wire          compressDataVec_hitReq_18_133;
  assign compressDataVec_hitReq_18_133 = _GEN_180;
  wire          _GEN_181 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h5;
  wire          compressDataVec_hitReq_19_5;
  assign compressDataVec_hitReq_19_5 = _GEN_181;
  wire          compressDataVec_hitReq_19_133;
  assign compressDataVec_hitReq_19_133 = _GEN_181;
  wire          _GEN_182 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h5;
  wire          compressDataVec_hitReq_20_5;
  assign compressDataVec_hitReq_20_5 = _GEN_182;
  wire          compressDataVec_hitReq_20_133;
  assign compressDataVec_hitReq_20_133 = _GEN_182;
  wire          _GEN_183 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h5;
  wire          compressDataVec_hitReq_21_5;
  assign compressDataVec_hitReq_21_5 = _GEN_183;
  wire          compressDataVec_hitReq_21_133;
  assign compressDataVec_hitReq_21_133 = _GEN_183;
  wire          _GEN_184 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h5;
  wire          compressDataVec_hitReq_22_5;
  assign compressDataVec_hitReq_22_5 = _GEN_184;
  wire          compressDataVec_hitReq_22_133;
  assign compressDataVec_hitReq_22_133 = _GEN_184;
  wire          _GEN_185 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h5;
  wire          compressDataVec_hitReq_23_5;
  assign compressDataVec_hitReq_23_5 = _GEN_185;
  wire          compressDataVec_hitReq_23_133;
  assign compressDataVec_hitReq_23_133 = _GEN_185;
  wire          _GEN_186 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h5;
  wire          compressDataVec_hitReq_24_5;
  assign compressDataVec_hitReq_24_5 = _GEN_186;
  wire          compressDataVec_hitReq_24_133;
  assign compressDataVec_hitReq_24_133 = _GEN_186;
  wire          _GEN_187 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h5;
  wire          compressDataVec_hitReq_25_5;
  assign compressDataVec_hitReq_25_5 = _GEN_187;
  wire          compressDataVec_hitReq_25_133;
  assign compressDataVec_hitReq_25_133 = _GEN_187;
  wire          _GEN_188 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h5;
  wire          compressDataVec_hitReq_26_5;
  assign compressDataVec_hitReq_26_5 = _GEN_188;
  wire          compressDataVec_hitReq_26_133;
  assign compressDataVec_hitReq_26_133 = _GEN_188;
  wire          _GEN_189 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h5;
  wire          compressDataVec_hitReq_27_5;
  assign compressDataVec_hitReq_27_5 = _GEN_189;
  wire          compressDataVec_hitReq_27_133;
  assign compressDataVec_hitReq_27_133 = _GEN_189;
  wire          _GEN_190 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h5;
  wire          compressDataVec_hitReq_28_5;
  assign compressDataVec_hitReq_28_5 = _GEN_190;
  wire          compressDataVec_hitReq_28_133;
  assign compressDataVec_hitReq_28_133 = _GEN_190;
  wire          _GEN_191 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h5;
  wire          compressDataVec_hitReq_29_5;
  assign compressDataVec_hitReq_29_5 = _GEN_191;
  wire          compressDataVec_hitReq_29_133;
  assign compressDataVec_hitReq_29_133 = _GEN_191;
  wire          _GEN_192 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h5;
  wire          compressDataVec_hitReq_30_5;
  assign compressDataVec_hitReq_30_5 = _GEN_192;
  wire          compressDataVec_hitReq_30_133;
  assign compressDataVec_hitReq_30_133 = _GEN_192;
  wire          _GEN_193 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h5;
  wire          compressDataVec_hitReq_31_5;
  assign compressDataVec_hitReq_31_5 = _GEN_193;
  wire          compressDataVec_hitReq_31_133;
  assign compressDataVec_hitReq_31_133 = _GEN_193;
  wire          compressDataVec_hitReq_32_5 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h5;
  wire          compressDataVec_hitReq_33_5 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h5;
  wire          compressDataVec_hitReq_34_5 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h5;
  wire          compressDataVec_hitReq_35_5 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h5;
  wire          compressDataVec_hitReq_36_5 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h5;
  wire          compressDataVec_hitReq_37_5 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h5;
  wire          compressDataVec_hitReq_38_5 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h5;
  wire          compressDataVec_hitReq_39_5 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h5;
  wire          compressDataVec_hitReq_40_5 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h5;
  wire          compressDataVec_hitReq_41_5 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h5;
  wire          compressDataVec_hitReq_42_5 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h5;
  wire          compressDataVec_hitReq_43_5 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h5;
  wire          compressDataVec_hitReq_44_5 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h5;
  wire          compressDataVec_hitReq_45_5 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h5;
  wire          compressDataVec_hitReq_46_5 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h5;
  wire          compressDataVec_hitReq_47_5 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h5;
  wire          compressDataVec_hitReq_48_5 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h5;
  wire          compressDataVec_hitReq_49_5 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h5;
  wire          compressDataVec_hitReq_50_5 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h5;
  wire          compressDataVec_hitReq_51_5 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h5;
  wire          compressDataVec_hitReq_52_5 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h5;
  wire          compressDataVec_hitReq_53_5 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h5;
  wire          compressDataVec_hitReq_54_5 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h5;
  wire          compressDataVec_hitReq_55_5 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h5;
  wire          compressDataVec_hitReq_56_5 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h5;
  wire          compressDataVec_hitReq_57_5 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h5;
  wire          compressDataVec_hitReq_58_5 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h5;
  wire          compressDataVec_hitReq_59_5 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h5;
  wire          compressDataVec_hitReq_60_5 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h5;
  wire          compressDataVec_hitReq_61_5 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h5;
  wire          compressDataVec_hitReq_62_5 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h5;
  wire          compressDataVec_hitReq_63_5 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h5;
  wire [7:0]    compressDataVec_selectReqData_5 =
    (compressDataVec_hitReq_0_5 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_5 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_5 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_5 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_5 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_5 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_5 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_5 ? source2Pipe[63:56] : 8'h0)
    | (compressDataVec_hitReq_8_5 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_5 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_5 ? source2Pipe[87:80] : 8'h0)
    | (compressDataVec_hitReq_11_5 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_5 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_5 ? source2Pipe[111:104] : 8'h0)
    | (compressDataVec_hitReq_14_5 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_5 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_5 ? source2Pipe[135:128] : 8'h0)
    | (compressDataVec_hitReq_17_5 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_5 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_5 ? source2Pipe[159:152] : 8'h0)
    | (compressDataVec_hitReq_20_5 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_5 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_5 ? source2Pipe[183:176] : 8'h0)
    | (compressDataVec_hitReq_23_5 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_5 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_5 ? source2Pipe[207:200] : 8'h0)
    | (compressDataVec_hitReq_26_5 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_5 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_5 ? source2Pipe[231:224] : 8'h0)
    | (compressDataVec_hitReq_29_5 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_5 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_5 ? source2Pipe[255:248] : 8'h0)
    | (compressDataVec_hitReq_32_5 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_5 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_5 ? source2Pipe[279:272] : 8'h0)
    | (compressDataVec_hitReq_35_5 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_5 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_5 ? source2Pipe[303:296] : 8'h0)
    | (compressDataVec_hitReq_38_5 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_5 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_5 ? source2Pipe[327:320] : 8'h0)
    | (compressDataVec_hitReq_41_5 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_5 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_5 ? source2Pipe[351:344] : 8'h0)
    | (compressDataVec_hitReq_44_5 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_5 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_5 ? source2Pipe[375:368] : 8'h0)
    | (compressDataVec_hitReq_47_5 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_5 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_5 ? source2Pipe[399:392] : 8'h0)
    | (compressDataVec_hitReq_50_5 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_5 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_5 ? source2Pipe[423:416] : 8'h0)
    | (compressDataVec_hitReq_53_5 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_5 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_5 ? source2Pipe[447:440] : 8'h0)
    | (compressDataVec_hitReq_56_5 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_5 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_5 ? source2Pipe[471:464] : 8'h0)
    | (compressDataVec_hitReq_59_5 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_5 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_5 ? source2Pipe[495:488] : 8'h0)
    | (compressDataVec_hitReq_62_5 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_5 ? source2Pipe[511:504] : 8'h0);
  wire          _GEN_194 = tailCount > 6'h5;
  wire          compressDataVec_useTail_5;
  assign compressDataVec_useTail_5 = _GEN_194;
  wire          compressDataVec_useTail_69;
  assign compressDataVec_useTail_69 = _GEN_194;
  wire          compressDataVec_useTail_101;
  assign compressDataVec_useTail_101 = _GEN_194;
  wire          _GEN_195 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h6;
  wire          compressDataVec_hitReq_0_6;
  assign compressDataVec_hitReq_0_6 = _GEN_195;
  wire          compressDataVec_hitReq_0_134;
  assign compressDataVec_hitReq_0_134 = _GEN_195;
  wire          compressDataVec_hitReq_0_198;
  assign compressDataVec_hitReq_0_198 = _GEN_195;
  wire          _GEN_196 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h6;
  wire          compressDataVec_hitReq_1_6;
  assign compressDataVec_hitReq_1_6 = _GEN_196;
  wire          compressDataVec_hitReq_1_134;
  assign compressDataVec_hitReq_1_134 = _GEN_196;
  wire          compressDataVec_hitReq_1_198;
  assign compressDataVec_hitReq_1_198 = _GEN_196;
  wire          _GEN_197 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h6;
  wire          compressDataVec_hitReq_2_6;
  assign compressDataVec_hitReq_2_6 = _GEN_197;
  wire          compressDataVec_hitReq_2_134;
  assign compressDataVec_hitReq_2_134 = _GEN_197;
  wire          compressDataVec_hitReq_2_198;
  assign compressDataVec_hitReq_2_198 = _GEN_197;
  wire          _GEN_198 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h6;
  wire          compressDataVec_hitReq_3_6;
  assign compressDataVec_hitReq_3_6 = _GEN_198;
  wire          compressDataVec_hitReq_3_134;
  assign compressDataVec_hitReq_3_134 = _GEN_198;
  wire          compressDataVec_hitReq_3_198;
  assign compressDataVec_hitReq_3_198 = _GEN_198;
  wire          _GEN_199 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h6;
  wire          compressDataVec_hitReq_4_6;
  assign compressDataVec_hitReq_4_6 = _GEN_199;
  wire          compressDataVec_hitReq_4_134;
  assign compressDataVec_hitReq_4_134 = _GEN_199;
  wire          compressDataVec_hitReq_4_198;
  assign compressDataVec_hitReq_4_198 = _GEN_199;
  wire          _GEN_200 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h6;
  wire          compressDataVec_hitReq_5_6;
  assign compressDataVec_hitReq_5_6 = _GEN_200;
  wire          compressDataVec_hitReq_5_134;
  assign compressDataVec_hitReq_5_134 = _GEN_200;
  wire          compressDataVec_hitReq_5_198;
  assign compressDataVec_hitReq_5_198 = _GEN_200;
  wire          _GEN_201 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h6;
  wire          compressDataVec_hitReq_6_6;
  assign compressDataVec_hitReq_6_6 = _GEN_201;
  wire          compressDataVec_hitReq_6_134;
  assign compressDataVec_hitReq_6_134 = _GEN_201;
  wire          compressDataVec_hitReq_6_198;
  assign compressDataVec_hitReq_6_198 = _GEN_201;
  wire          _GEN_202 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h6;
  wire          compressDataVec_hitReq_7_6;
  assign compressDataVec_hitReq_7_6 = _GEN_202;
  wire          compressDataVec_hitReq_7_134;
  assign compressDataVec_hitReq_7_134 = _GEN_202;
  wire          compressDataVec_hitReq_7_198;
  assign compressDataVec_hitReq_7_198 = _GEN_202;
  wire          _GEN_203 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h6;
  wire          compressDataVec_hitReq_8_6;
  assign compressDataVec_hitReq_8_6 = _GEN_203;
  wire          compressDataVec_hitReq_8_134;
  assign compressDataVec_hitReq_8_134 = _GEN_203;
  wire          compressDataVec_hitReq_8_198;
  assign compressDataVec_hitReq_8_198 = _GEN_203;
  wire          _GEN_204 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h6;
  wire          compressDataVec_hitReq_9_6;
  assign compressDataVec_hitReq_9_6 = _GEN_204;
  wire          compressDataVec_hitReq_9_134;
  assign compressDataVec_hitReq_9_134 = _GEN_204;
  wire          compressDataVec_hitReq_9_198;
  assign compressDataVec_hitReq_9_198 = _GEN_204;
  wire          _GEN_205 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h6;
  wire          compressDataVec_hitReq_10_6;
  assign compressDataVec_hitReq_10_6 = _GEN_205;
  wire          compressDataVec_hitReq_10_134;
  assign compressDataVec_hitReq_10_134 = _GEN_205;
  wire          compressDataVec_hitReq_10_198;
  assign compressDataVec_hitReq_10_198 = _GEN_205;
  wire          _GEN_206 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h6;
  wire          compressDataVec_hitReq_11_6;
  assign compressDataVec_hitReq_11_6 = _GEN_206;
  wire          compressDataVec_hitReq_11_134;
  assign compressDataVec_hitReq_11_134 = _GEN_206;
  wire          compressDataVec_hitReq_11_198;
  assign compressDataVec_hitReq_11_198 = _GEN_206;
  wire          _GEN_207 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h6;
  wire          compressDataVec_hitReq_12_6;
  assign compressDataVec_hitReq_12_6 = _GEN_207;
  wire          compressDataVec_hitReq_12_134;
  assign compressDataVec_hitReq_12_134 = _GEN_207;
  wire          compressDataVec_hitReq_12_198;
  assign compressDataVec_hitReq_12_198 = _GEN_207;
  wire          _GEN_208 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h6;
  wire          compressDataVec_hitReq_13_6;
  assign compressDataVec_hitReq_13_6 = _GEN_208;
  wire          compressDataVec_hitReq_13_134;
  assign compressDataVec_hitReq_13_134 = _GEN_208;
  wire          compressDataVec_hitReq_13_198;
  assign compressDataVec_hitReq_13_198 = _GEN_208;
  wire          _GEN_209 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h6;
  wire          compressDataVec_hitReq_14_6;
  assign compressDataVec_hitReq_14_6 = _GEN_209;
  wire          compressDataVec_hitReq_14_134;
  assign compressDataVec_hitReq_14_134 = _GEN_209;
  wire          compressDataVec_hitReq_14_198;
  assign compressDataVec_hitReq_14_198 = _GEN_209;
  wire          _GEN_210 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h6;
  wire          compressDataVec_hitReq_15_6;
  assign compressDataVec_hitReq_15_6 = _GEN_210;
  wire          compressDataVec_hitReq_15_134;
  assign compressDataVec_hitReq_15_134 = _GEN_210;
  wire          compressDataVec_hitReq_15_198;
  assign compressDataVec_hitReq_15_198 = _GEN_210;
  wire          _GEN_211 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h6;
  wire          compressDataVec_hitReq_16_6;
  assign compressDataVec_hitReq_16_6 = _GEN_211;
  wire          compressDataVec_hitReq_16_134;
  assign compressDataVec_hitReq_16_134 = _GEN_211;
  wire          _GEN_212 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h6;
  wire          compressDataVec_hitReq_17_6;
  assign compressDataVec_hitReq_17_6 = _GEN_212;
  wire          compressDataVec_hitReq_17_134;
  assign compressDataVec_hitReq_17_134 = _GEN_212;
  wire          _GEN_213 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h6;
  wire          compressDataVec_hitReq_18_6;
  assign compressDataVec_hitReq_18_6 = _GEN_213;
  wire          compressDataVec_hitReq_18_134;
  assign compressDataVec_hitReq_18_134 = _GEN_213;
  wire          _GEN_214 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h6;
  wire          compressDataVec_hitReq_19_6;
  assign compressDataVec_hitReq_19_6 = _GEN_214;
  wire          compressDataVec_hitReq_19_134;
  assign compressDataVec_hitReq_19_134 = _GEN_214;
  wire          _GEN_215 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h6;
  wire          compressDataVec_hitReq_20_6;
  assign compressDataVec_hitReq_20_6 = _GEN_215;
  wire          compressDataVec_hitReq_20_134;
  assign compressDataVec_hitReq_20_134 = _GEN_215;
  wire          _GEN_216 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h6;
  wire          compressDataVec_hitReq_21_6;
  assign compressDataVec_hitReq_21_6 = _GEN_216;
  wire          compressDataVec_hitReq_21_134;
  assign compressDataVec_hitReq_21_134 = _GEN_216;
  wire          _GEN_217 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h6;
  wire          compressDataVec_hitReq_22_6;
  assign compressDataVec_hitReq_22_6 = _GEN_217;
  wire          compressDataVec_hitReq_22_134;
  assign compressDataVec_hitReq_22_134 = _GEN_217;
  wire          _GEN_218 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h6;
  wire          compressDataVec_hitReq_23_6;
  assign compressDataVec_hitReq_23_6 = _GEN_218;
  wire          compressDataVec_hitReq_23_134;
  assign compressDataVec_hitReq_23_134 = _GEN_218;
  wire          _GEN_219 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h6;
  wire          compressDataVec_hitReq_24_6;
  assign compressDataVec_hitReq_24_6 = _GEN_219;
  wire          compressDataVec_hitReq_24_134;
  assign compressDataVec_hitReq_24_134 = _GEN_219;
  wire          _GEN_220 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h6;
  wire          compressDataVec_hitReq_25_6;
  assign compressDataVec_hitReq_25_6 = _GEN_220;
  wire          compressDataVec_hitReq_25_134;
  assign compressDataVec_hitReq_25_134 = _GEN_220;
  wire          _GEN_221 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h6;
  wire          compressDataVec_hitReq_26_6;
  assign compressDataVec_hitReq_26_6 = _GEN_221;
  wire          compressDataVec_hitReq_26_134;
  assign compressDataVec_hitReq_26_134 = _GEN_221;
  wire          _GEN_222 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h6;
  wire          compressDataVec_hitReq_27_6;
  assign compressDataVec_hitReq_27_6 = _GEN_222;
  wire          compressDataVec_hitReq_27_134;
  assign compressDataVec_hitReq_27_134 = _GEN_222;
  wire          _GEN_223 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h6;
  wire          compressDataVec_hitReq_28_6;
  assign compressDataVec_hitReq_28_6 = _GEN_223;
  wire          compressDataVec_hitReq_28_134;
  assign compressDataVec_hitReq_28_134 = _GEN_223;
  wire          _GEN_224 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h6;
  wire          compressDataVec_hitReq_29_6;
  assign compressDataVec_hitReq_29_6 = _GEN_224;
  wire          compressDataVec_hitReq_29_134;
  assign compressDataVec_hitReq_29_134 = _GEN_224;
  wire          _GEN_225 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h6;
  wire          compressDataVec_hitReq_30_6;
  assign compressDataVec_hitReq_30_6 = _GEN_225;
  wire          compressDataVec_hitReq_30_134;
  assign compressDataVec_hitReq_30_134 = _GEN_225;
  wire          _GEN_226 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h6;
  wire          compressDataVec_hitReq_31_6;
  assign compressDataVec_hitReq_31_6 = _GEN_226;
  wire          compressDataVec_hitReq_31_134;
  assign compressDataVec_hitReq_31_134 = _GEN_226;
  wire          compressDataVec_hitReq_32_6 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h6;
  wire          compressDataVec_hitReq_33_6 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h6;
  wire          compressDataVec_hitReq_34_6 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h6;
  wire          compressDataVec_hitReq_35_6 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h6;
  wire          compressDataVec_hitReq_36_6 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h6;
  wire          compressDataVec_hitReq_37_6 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h6;
  wire          compressDataVec_hitReq_38_6 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h6;
  wire          compressDataVec_hitReq_39_6 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h6;
  wire          compressDataVec_hitReq_40_6 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h6;
  wire          compressDataVec_hitReq_41_6 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h6;
  wire          compressDataVec_hitReq_42_6 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h6;
  wire          compressDataVec_hitReq_43_6 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h6;
  wire          compressDataVec_hitReq_44_6 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h6;
  wire          compressDataVec_hitReq_45_6 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h6;
  wire          compressDataVec_hitReq_46_6 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h6;
  wire          compressDataVec_hitReq_47_6 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h6;
  wire          compressDataVec_hitReq_48_6 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h6;
  wire          compressDataVec_hitReq_49_6 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h6;
  wire          compressDataVec_hitReq_50_6 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h6;
  wire          compressDataVec_hitReq_51_6 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h6;
  wire          compressDataVec_hitReq_52_6 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h6;
  wire          compressDataVec_hitReq_53_6 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h6;
  wire          compressDataVec_hitReq_54_6 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h6;
  wire          compressDataVec_hitReq_55_6 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h6;
  wire          compressDataVec_hitReq_56_6 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h6;
  wire          compressDataVec_hitReq_57_6 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h6;
  wire          compressDataVec_hitReq_58_6 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h6;
  wire          compressDataVec_hitReq_59_6 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h6;
  wire          compressDataVec_hitReq_60_6 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h6;
  wire          compressDataVec_hitReq_61_6 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h6;
  wire          compressDataVec_hitReq_62_6 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h6;
  wire          compressDataVec_hitReq_63_6 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h6;
  wire [7:0]    compressDataVec_selectReqData_6 =
    (compressDataVec_hitReq_0_6 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_6 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_6 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_6 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_6 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_6 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_6 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_6 ? source2Pipe[63:56] : 8'h0)
    | (compressDataVec_hitReq_8_6 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_6 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_6 ? source2Pipe[87:80] : 8'h0)
    | (compressDataVec_hitReq_11_6 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_6 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_6 ? source2Pipe[111:104] : 8'h0)
    | (compressDataVec_hitReq_14_6 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_6 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_6 ? source2Pipe[135:128] : 8'h0)
    | (compressDataVec_hitReq_17_6 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_6 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_6 ? source2Pipe[159:152] : 8'h0)
    | (compressDataVec_hitReq_20_6 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_6 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_6 ? source2Pipe[183:176] : 8'h0)
    | (compressDataVec_hitReq_23_6 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_6 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_6 ? source2Pipe[207:200] : 8'h0)
    | (compressDataVec_hitReq_26_6 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_6 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_6 ? source2Pipe[231:224] : 8'h0)
    | (compressDataVec_hitReq_29_6 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_6 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_6 ? source2Pipe[255:248] : 8'h0)
    | (compressDataVec_hitReq_32_6 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_6 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_6 ? source2Pipe[279:272] : 8'h0)
    | (compressDataVec_hitReq_35_6 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_6 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_6 ? source2Pipe[303:296] : 8'h0)
    | (compressDataVec_hitReq_38_6 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_6 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_6 ? source2Pipe[327:320] : 8'h0)
    | (compressDataVec_hitReq_41_6 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_6 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_6 ? source2Pipe[351:344] : 8'h0)
    | (compressDataVec_hitReq_44_6 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_6 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_6 ? source2Pipe[375:368] : 8'h0)
    | (compressDataVec_hitReq_47_6 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_6 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_6 ? source2Pipe[399:392] : 8'h0)
    | (compressDataVec_hitReq_50_6 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_6 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_6 ? source2Pipe[423:416] : 8'h0)
    | (compressDataVec_hitReq_53_6 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_6 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_6 ? source2Pipe[447:440] : 8'h0)
    | (compressDataVec_hitReq_56_6 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_6 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_6 ? source2Pipe[471:464] : 8'h0)
    | (compressDataVec_hitReq_59_6 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_6 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_6 ? source2Pipe[495:488] : 8'h0)
    | (compressDataVec_hitReq_62_6 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_6 ? source2Pipe[511:504] : 8'h0);
  wire          _GEN_227 = tailCount > 6'h6;
  wire          compressDataVec_useTail_6;
  assign compressDataVec_useTail_6 = _GEN_227;
  wire          compressDataVec_useTail_70;
  assign compressDataVec_useTail_70 = _GEN_227;
  wire          compressDataVec_useTail_102;
  assign compressDataVec_useTail_102 = _GEN_227;
  wire          _GEN_228 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h7;
  wire          compressDataVec_hitReq_0_7;
  assign compressDataVec_hitReq_0_7 = _GEN_228;
  wire          compressDataVec_hitReq_0_135;
  assign compressDataVec_hitReq_0_135 = _GEN_228;
  wire          compressDataVec_hitReq_0_199;
  assign compressDataVec_hitReq_0_199 = _GEN_228;
  wire          _GEN_229 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h7;
  wire          compressDataVec_hitReq_1_7;
  assign compressDataVec_hitReq_1_7 = _GEN_229;
  wire          compressDataVec_hitReq_1_135;
  assign compressDataVec_hitReq_1_135 = _GEN_229;
  wire          compressDataVec_hitReq_1_199;
  assign compressDataVec_hitReq_1_199 = _GEN_229;
  wire          _GEN_230 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h7;
  wire          compressDataVec_hitReq_2_7;
  assign compressDataVec_hitReq_2_7 = _GEN_230;
  wire          compressDataVec_hitReq_2_135;
  assign compressDataVec_hitReq_2_135 = _GEN_230;
  wire          compressDataVec_hitReq_2_199;
  assign compressDataVec_hitReq_2_199 = _GEN_230;
  wire          _GEN_231 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h7;
  wire          compressDataVec_hitReq_3_7;
  assign compressDataVec_hitReq_3_7 = _GEN_231;
  wire          compressDataVec_hitReq_3_135;
  assign compressDataVec_hitReq_3_135 = _GEN_231;
  wire          compressDataVec_hitReq_3_199;
  assign compressDataVec_hitReq_3_199 = _GEN_231;
  wire          _GEN_232 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h7;
  wire          compressDataVec_hitReq_4_7;
  assign compressDataVec_hitReq_4_7 = _GEN_232;
  wire          compressDataVec_hitReq_4_135;
  assign compressDataVec_hitReq_4_135 = _GEN_232;
  wire          compressDataVec_hitReq_4_199;
  assign compressDataVec_hitReq_4_199 = _GEN_232;
  wire          _GEN_233 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h7;
  wire          compressDataVec_hitReq_5_7;
  assign compressDataVec_hitReq_5_7 = _GEN_233;
  wire          compressDataVec_hitReq_5_135;
  assign compressDataVec_hitReq_5_135 = _GEN_233;
  wire          compressDataVec_hitReq_5_199;
  assign compressDataVec_hitReq_5_199 = _GEN_233;
  wire          _GEN_234 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h7;
  wire          compressDataVec_hitReq_6_7;
  assign compressDataVec_hitReq_6_7 = _GEN_234;
  wire          compressDataVec_hitReq_6_135;
  assign compressDataVec_hitReq_6_135 = _GEN_234;
  wire          compressDataVec_hitReq_6_199;
  assign compressDataVec_hitReq_6_199 = _GEN_234;
  wire          _GEN_235 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h7;
  wire          compressDataVec_hitReq_7_7;
  assign compressDataVec_hitReq_7_7 = _GEN_235;
  wire          compressDataVec_hitReq_7_135;
  assign compressDataVec_hitReq_7_135 = _GEN_235;
  wire          compressDataVec_hitReq_7_199;
  assign compressDataVec_hitReq_7_199 = _GEN_235;
  wire          _GEN_236 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h7;
  wire          compressDataVec_hitReq_8_7;
  assign compressDataVec_hitReq_8_7 = _GEN_236;
  wire          compressDataVec_hitReq_8_135;
  assign compressDataVec_hitReq_8_135 = _GEN_236;
  wire          compressDataVec_hitReq_8_199;
  assign compressDataVec_hitReq_8_199 = _GEN_236;
  wire          _GEN_237 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h7;
  wire          compressDataVec_hitReq_9_7;
  assign compressDataVec_hitReq_9_7 = _GEN_237;
  wire          compressDataVec_hitReq_9_135;
  assign compressDataVec_hitReq_9_135 = _GEN_237;
  wire          compressDataVec_hitReq_9_199;
  assign compressDataVec_hitReq_9_199 = _GEN_237;
  wire          _GEN_238 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h7;
  wire          compressDataVec_hitReq_10_7;
  assign compressDataVec_hitReq_10_7 = _GEN_238;
  wire          compressDataVec_hitReq_10_135;
  assign compressDataVec_hitReq_10_135 = _GEN_238;
  wire          compressDataVec_hitReq_10_199;
  assign compressDataVec_hitReq_10_199 = _GEN_238;
  wire          _GEN_239 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h7;
  wire          compressDataVec_hitReq_11_7;
  assign compressDataVec_hitReq_11_7 = _GEN_239;
  wire          compressDataVec_hitReq_11_135;
  assign compressDataVec_hitReq_11_135 = _GEN_239;
  wire          compressDataVec_hitReq_11_199;
  assign compressDataVec_hitReq_11_199 = _GEN_239;
  wire          _GEN_240 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h7;
  wire          compressDataVec_hitReq_12_7;
  assign compressDataVec_hitReq_12_7 = _GEN_240;
  wire          compressDataVec_hitReq_12_135;
  assign compressDataVec_hitReq_12_135 = _GEN_240;
  wire          compressDataVec_hitReq_12_199;
  assign compressDataVec_hitReq_12_199 = _GEN_240;
  wire          _GEN_241 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h7;
  wire          compressDataVec_hitReq_13_7;
  assign compressDataVec_hitReq_13_7 = _GEN_241;
  wire          compressDataVec_hitReq_13_135;
  assign compressDataVec_hitReq_13_135 = _GEN_241;
  wire          compressDataVec_hitReq_13_199;
  assign compressDataVec_hitReq_13_199 = _GEN_241;
  wire          _GEN_242 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h7;
  wire          compressDataVec_hitReq_14_7;
  assign compressDataVec_hitReq_14_7 = _GEN_242;
  wire          compressDataVec_hitReq_14_135;
  assign compressDataVec_hitReq_14_135 = _GEN_242;
  wire          compressDataVec_hitReq_14_199;
  assign compressDataVec_hitReq_14_199 = _GEN_242;
  wire          _GEN_243 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h7;
  wire          compressDataVec_hitReq_15_7;
  assign compressDataVec_hitReq_15_7 = _GEN_243;
  wire          compressDataVec_hitReq_15_135;
  assign compressDataVec_hitReq_15_135 = _GEN_243;
  wire          compressDataVec_hitReq_15_199;
  assign compressDataVec_hitReq_15_199 = _GEN_243;
  wire          _GEN_244 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h7;
  wire          compressDataVec_hitReq_16_7;
  assign compressDataVec_hitReq_16_7 = _GEN_244;
  wire          compressDataVec_hitReq_16_135;
  assign compressDataVec_hitReq_16_135 = _GEN_244;
  wire          _GEN_245 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h7;
  wire          compressDataVec_hitReq_17_7;
  assign compressDataVec_hitReq_17_7 = _GEN_245;
  wire          compressDataVec_hitReq_17_135;
  assign compressDataVec_hitReq_17_135 = _GEN_245;
  wire          _GEN_246 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h7;
  wire          compressDataVec_hitReq_18_7;
  assign compressDataVec_hitReq_18_7 = _GEN_246;
  wire          compressDataVec_hitReq_18_135;
  assign compressDataVec_hitReq_18_135 = _GEN_246;
  wire          _GEN_247 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h7;
  wire          compressDataVec_hitReq_19_7;
  assign compressDataVec_hitReq_19_7 = _GEN_247;
  wire          compressDataVec_hitReq_19_135;
  assign compressDataVec_hitReq_19_135 = _GEN_247;
  wire          _GEN_248 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h7;
  wire          compressDataVec_hitReq_20_7;
  assign compressDataVec_hitReq_20_7 = _GEN_248;
  wire          compressDataVec_hitReq_20_135;
  assign compressDataVec_hitReq_20_135 = _GEN_248;
  wire          _GEN_249 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h7;
  wire          compressDataVec_hitReq_21_7;
  assign compressDataVec_hitReq_21_7 = _GEN_249;
  wire          compressDataVec_hitReq_21_135;
  assign compressDataVec_hitReq_21_135 = _GEN_249;
  wire          _GEN_250 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h7;
  wire          compressDataVec_hitReq_22_7;
  assign compressDataVec_hitReq_22_7 = _GEN_250;
  wire          compressDataVec_hitReq_22_135;
  assign compressDataVec_hitReq_22_135 = _GEN_250;
  wire          _GEN_251 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h7;
  wire          compressDataVec_hitReq_23_7;
  assign compressDataVec_hitReq_23_7 = _GEN_251;
  wire          compressDataVec_hitReq_23_135;
  assign compressDataVec_hitReq_23_135 = _GEN_251;
  wire          _GEN_252 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h7;
  wire          compressDataVec_hitReq_24_7;
  assign compressDataVec_hitReq_24_7 = _GEN_252;
  wire          compressDataVec_hitReq_24_135;
  assign compressDataVec_hitReq_24_135 = _GEN_252;
  wire          _GEN_253 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h7;
  wire          compressDataVec_hitReq_25_7;
  assign compressDataVec_hitReq_25_7 = _GEN_253;
  wire          compressDataVec_hitReq_25_135;
  assign compressDataVec_hitReq_25_135 = _GEN_253;
  wire          _GEN_254 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h7;
  wire          compressDataVec_hitReq_26_7;
  assign compressDataVec_hitReq_26_7 = _GEN_254;
  wire          compressDataVec_hitReq_26_135;
  assign compressDataVec_hitReq_26_135 = _GEN_254;
  wire          _GEN_255 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h7;
  wire          compressDataVec_hitReq_27_7;
  assign compressDataVec_hitReq_27_7 = _GEN_255;
  wire          compressDataVec_hitReq_27_135;
  assign compressDataVec_hitReq_27_135 = _GEN_255;
  wire          _GEN_256 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h7;
  wire          compressDataVec_hitReq_28_7;
  assign compressDataVec_hitReq_28_7 = _GEN_256;
  wire          compressDataVec_hitReq_28_135;
  assign compressDataVec_hitReq_28_135 = _GEN_256;
  wire          _GEN_257 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h7;
  wire          compressDataVec_hitReq_29_7;
  assign compressDataVec_hitReq_29_7 = _GEN_257;
  wire          compressDataVec_hitReq_29_135;
  assign compressDataVec_hitReq_29_135 = _GEN_257;
  wire          _GEN_258 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h7;
  wire          compressDataVec_hitReq_30_7;
  assign compressDataVec_hitReq_30_7 = _GEN_258;
  wire          compressDataVec_hitReq_30_135;
  assign compressDataVec_hitReq_30_135 = _GEN_258;
  wire          _GEN_259 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h7;
  wire          compressDataVec_hitReq_31_7;
  assign compressDataVec_hitReq_31_7 = _GEN_259;
  wire          compressDataVec_hitReq_31_135;
  assign compressDataVec_hitReq_31_135 = _GEN_259;
  wire          compressDataVec_hitReq_32_7 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h7;
  wire          compressDataVec_hitReq_33_7 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h7;
  wire          compressDataVec_hitReq_34_7 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h7;
  wire          compressDataVec_hitReq_35_7 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h7;
  wire          compressDataVec_hitReq_36_7 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h7;
  wire          compressDataVec_hitReq_37_7 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h7;
  wire          compressDataVec_hitReq_38_7 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h7;
  wire          compressDataVec_hitReq_39_7 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h7;
  wire          compressDataVec_hitReq_40_7 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h7;
  wire          compressDataVec_hitReq_41_7 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h7;
  wire          compressDataVec_hitReq_42_7 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h7;
  wire          compressDataVec_hitReq_43_7 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h7;
  wire          compressDataVec_hitReq_44_7 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h7;
  wire          compressDataVec_hitReq_45_7 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h7;
  wire          compressDataVec_hitReq_46_7 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h7;
  wire          compressDataVec_hitReq_47_7 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h7;
  wire          compressDataVec_hitReq_48_7 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h7;
  wire          compressDataVec_hitReq_49_7 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h7;
  wire          compressDataVec_hitReq_50_7 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h7;
  wire          compressDataVec_hitReq_51_7 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h7;
  wire          compressDataVec_hitReq_52_7 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h7;
  wire          compressDataVec_hitReq_53_7 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h7;
  wire          compressDataVec_hitReq_54_7 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h7;
  wire          compressDataVec_hitReq_55_7 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h7;
  wire          compressDataVec_hitReq_56_7 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h7;
  wire          compressDataVec_hitReq_57_7 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h7;
  wire          compressDataVec_hitReq_58_7 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h7;
  wire          compressDataVec_hitReq_59_7 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h7;
  wire          compressDataVec_hitReq_60_7 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h7;
  wire          compressDataVec_hitReq_61_7 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h7;
  wire          compressDataVec_hitReq_62_7 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h7;
  wire          compressDataVec_hitReq_63_7 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h7;
  wire [7:0]    compressDataVec_selectReqData_7 =
    (compressDataVec_hitReq_0_7 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_7 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_7 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_7 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_7 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_7 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_7 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_7 ? source2Pipe[63:56] : 8'h0)
    | (compressDataVec_hitReq_8_7 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_7 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_7 ? source2Pipe[87:80] : 8'h0)
    | (compressDataVec_hitReq_11_7 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_7 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_7 ? source2Pipe[111:104] : 8'h0)
    | (compressDataVec_hitReq_14_7 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_7 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_7 ? source2Pipe[135:128] : 8'h0)
    | (compressDataVec_hitReq_17_7 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_7 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_7 ? source2Pipe[159:152] : 8'h0)
    | (compressDataVec_hitReq_20_7 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_7 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_7 ? source2Pipe[183:176] : 8'h0)
    | (compressDataVec_hitReq_23_7 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_7 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_7 ? source2Pipe[207:200] : 8'h0)
    | (compressDataVec_hitReq_26_7 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_7 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_7 ? source2Pipe[231:224] : 8'h0)
    | (compressDataVec_hitReq_29_7 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_7 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_7 ? source2Pipe[255:248] : 8'h0)
    | (compressDataVec_hitReq_32_7 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_7 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_7 ? source2Pipe[279:272] : 8'h0)
    | (compressDataVec_hitReq_35_7 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_7 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_7 ? source2Pipe[303:296] : 8'h0)
    | (compressDataVec_hitReq_38_7 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_7 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_7 ? source2Pipe[327:320] : 8'h0)
    | (compressDataVec_hitReq_41_7 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_7 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_7 ? source2Pipe[351:344] : 8'h0)
    | (compressDataVec_hitReq_44_7 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_7 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_7 ? source2Pipe[375:368] : 8'h0)
    | (compressDataVec_hitReq_47_7 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_7 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_7 ? source2Pipe[399:392] : 8'h0)
    | (compressDataVec_hitReq_50_7 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_7 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_7 ? source2Pipe[423:416] : 8'h0)
    | (compressDataVec_hitReq_53_7 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_7 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_7 ? source2Pipe[447:440] : 8'h0)
    | (compressDataVec_hitReq_56_7 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_7 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_7 ? source2Pipe[471:464] : 8'h0)
    | (compressDataVec_hitReq_59_7 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_7 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_7 ? source2Pipe[495:488] : 8'h0)
    | (compressDataVec_hitReq_62_7 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_7 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_7;
  assign compressDataVec_useTail_7 = |(tailCount[5:3]);
  wire          _GEN_260 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h8;
  wire          compressDataVec_hitReq_0_8;
  assign compressDataVec_hitReq_0_8 = _GEN_260;
  wire          compressDataVec_hitReq_0_136;
  assign compressDataVec_hitReq_0_136 = _GEN_260;
  wire          compressDataVec_hitReq_0_200;
  assign compressDataVec_hitReq_0_200 = _GEN_260;
  wire          _GEN_261 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h8;
  wire          compressDataVec_hitReq_1_8;
  assign compressDataVec_hitReq_1_8 = _GEN_261;
  wire          compressDataVec_hitReq_1_136;
  assign compressDataVec_hitReq_1_136 = _GEN_261;
  wire          compressDataVec_hitReq_1_200;
  assign compressDataVec_hitReq_1_200 = _GEN_261;
  wire          _GEN_262 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h8;
  wire          compressDataVec_hitReq_2_8;
  assign compressDataVec_hitReq_2_8 = _GEN_262;
  wire          compressDataVec_hitReq_2_136;
  assign compressDataVec_hitReq_2_136 = _GEN_262;
  wire          compressDataVec_hitReq_2_200;
  assign compressDataVec_hitReq_2_200 = _GEN_262;
  wire          _GEN_263 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h8;
  wire          compressDataVec_hitReq_3_8;
  assign compressDataVec_hitReq_3_8 = _GEN_263;
  wire          compressDataVec_hitReq_3_136;
  assign compressDataVec_hitReq_3_136 = _GEN_263;
  wire          compressDataVec_hitReq_3_200;
  assign compressDataVec_hitReq_3_200 = _GEN_263;
  wire          _GEN_264 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h8;
  wire          compressDataVec_hitReq_4_8;
  assign compressDataVec_hitReq_4_8 = _GEN_264;
  wire          compressDataVec_hitReq_4_136;
  assign compressDataVec_hitReq_4_136 = _GEN_264;
  wire          compressDataVec_hitReq_4_200;
  assign compressDataVec_hitReq_4_200 = _GEN_264;
  wire          _GEN_265 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h8;
  wire          compressDataVec_hitReq_5_8;
  assign compressDataVec_hitReq_5_8 = _GEN_265;
  wire          compressDataVec_hitReq_5_136;
  assign compressDataVec_hitReq_5_136 = _GEN_265;
  wire          compressDataVec_hitReq_5_200;
  assign compressDataVec_hitReq_5_200 = _GEN_265;
  wire          _GEN_266 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h8;
  wire          compressDataVec_hitReq_6_8;
  assign compressDataVec_hitReq_6_8 = _GEN_266;
  wire          compressDataVec_hitReq_6_136;
  assign compressDataVec_hitReq_6_136 = _GEN_266;
  wire          compressDataVec_hitReq_6_200;
  assign compressDataVec_hitReq_6_200 = _GEN_266;
  wire          _GEN_267 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h8;
  wire          compressDataVec_hitReq_7_8;
  assign compressDataVec_hitReq_7_8 = _GEN_267;
  wire          compressDataVec_hitReq_7_136;
  assign compressDataVec_hitReq_7_136 = _GEN_267;
  wire          compressDataVec_hitReq_7_200;
  assign compressDataVec_hitReq_7_200 = _GEN_267;
  wire          _GEN_268 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h8;
  wire          compressDataVec_hitReq_8_8;
  assign compressDataVec_hitReq_8_8 = _GEN_268;
  wire          compressDataVec_hitReq_8_136;
  assign compressDataVec_hitReq_8_136 = _GEN_268;
  wire          compressDataVec_hitReq_8_200;
  assign compressDataVec_hitReq_8_200 = _GEN_268;
  wire          _GEN_269 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h8;
  wire          compressDataVec_hitReq_9_8;
  assign compressDataVec_hitReq_9_8 = _GEN_269;
  wire          compressDataVec_hitReq_9_136;
  assign compressDataVec_hitReq_9_136 = _GEN_269;
  wire          compressDataVec_hitReq_9_200;
  assign compressDataVec_hitReq_9_200 = _GEN_269;
  wire          _GEN_270 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h8;
  wire          compressDataVec_hitReq_10_8;
  assign compressDataVec_hitReq_10_8 = _GEN_270;
  wire          compressDataVec_hitReq_10_136;
  assign compressDataVec_hitReq_10_136 = _GEN_270;
  wire          compressDataVec_hitReq_10_200;
  assign compressDataVec_hitReq_10_200 = _GEN_270;
  wire          _GEN_271 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h8;
  wire          compressDataVec_hitReq_11_8;
  assign compressDataVec_hitReq_11_8 = _GEN_271;
  wire          compressDataVec_hitReq_11_136;
  assign compressDataVec_hitReq_11_136 = _GEN_271;
  wire          compressDataVec_hitReq_11_200;
  assign compressDataVec_hitReq_11_200 = _GEN_271;
  wire          _GEN_272 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h8;
  wire          compressDataVec_hitReq_12_8;
  assign compressDataVec_hitReq_12_8 = _GEN_272;
  wire          compressDataVec_hitReq_12_136;
  assign compressDataVec_hitReq_12_136 = _GEN_272;
  wire          compressDataVec_hitReq_12_200;
  assign compressDataVec_hitReq_12_200 = _GEN_272;
  wire          _GEN_273 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h8;
  wire          compressDataVec_hitReq_13_8;
  assign compressDataVec_hitReq_13_8 = _GEN_273;
  wire          compressDataVec_hitReq_13_136;
  assign compressDataVec_hitReq_13_136 = _GEN_273;
  wire          compressDataVec_hitReq_13_200;
  assign compressDataVec_hitReq_13_200 = _GEN_273;
  wire          _GEN_274 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h8;
  wire          compressDataVec_hitReq_14_8;
  assign compressDataVec_hitReq_14_8 = _GEN_274;
  wire          compressDataVec_hitReq_14_136;
  assign compressDataVec_hitReq_14_136 = _GEN_274;
  wire          compressDataVec_hitReq_14_200;
  assign compressDataVec_hitReq_14_200 = _GEN_274;
  wire          _GEN_275 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h8;
  wire          compressDataVec_hitReq_15_8;
  assign compressDataVec_hitReq_15_8 = _GEN_275;
  wire          compressDataVec_hitReq_15_136;
  assign compressDataVec_hitReq_15_136 = _GEN_275;
  wire          compressDataVec_hitReq_15_200;
  assign compressDataVec_hitReq_15_200 = _GEN_275;
  wire          _GEN_276 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h8;
  wire          compressDataVec_hitReq_16_8;
  assign compressDataVec_hitReq_16_8 = _GEN_276;
  wire          compressDataVec_hitReq_16_136;
  assign compressDataVec_hitReq_16_136 = _GEN_276;
  wire          _GEN_277 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h8;
  wire          compressDataVec_hitReq_17_8;
  assign compressDataVec_hitReq_17_8 = _GEN_277;
  wire          compressDataVec_hitReq_17_136;
  assign compressDataVec_hitReq_17_136 = _GEN_277;
  wire          _GEN_278 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h8;
  wire          compressDataVec_hitReq_18_8;
  assign compressDataVec_hitReq_18_8 = _GEN_278;
  wire          compressDataVec_hitReq_18_136;
  assign compressDataVec_hitReq_18_136 = _GEN_278;
  wire          _GEN_279 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h8;
  wire          compressDataVec_hitReq_19_8;
  assign compressDataVec_hitReq_19_8 = _GEN_279;
  wire          compressDataVec_hitReq_19_136;
  assign compressDataVec_hitReq_19_136 = _GEN_279;
  wire          _GEN_280 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h8;
  wire          compressDataVec_hitReq_20_8;
  assign compressDataVec_hitReq_20_8 = _GEN_280;
  wire          compressDataVec_hitReq_20_136;
  assign compressDataVec_hitReq_20_136 = _GEN_280;
  wire          _GEN_281 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h8;
  wire          compressDataVec_hitReq_21_8;
  assign compressDataVec_hitReq_21_8 = _GEN_281;
  wire          compressDataVec_hitReq_21_136;
  assign compressDataVec_hitReq_21_136 = _GEN_281;
  wire          _GEN_282 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h8;
  wire          compressDataVec_hitReq_22_8;
  assign compressDataVec_hitReq_22_8 = _GEN_282;
  wire          compressDataVec_hitReq_22_136;
  assign compressDataVec_hitReq_22_136 = _GEN_282;
  wire          _GEN_283 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h8;
  wire          compressDataVec_hitReq_23_8;
  assign compressDataVec_hitReq_23_8 = _GEN_283;
  wire          compressDataVec_hitReq_23_136;
  assign compressDataVec_hitReq_23_136 = _GEN_283;
  wire          _GEN_284 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h8;
  wire          compressDataVec_hitReq_24_8;
  assign compressDataVec_hitReq_24_8 = _GEN_284;
  wire          compressDataVec_hitReq_24_136;
  assign compressDataVec_hitReq_24_136 = _GEN_284;
  wire          _GEN_285 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h8;
  wire          compressDataVec_hitReq_25_8;
  assign compressDataVec_hitReq_25_8 = _GEN_285;
  wire          compressDataVec_hitReq_25_136;
  assign compressDataVec_hitReq_25_136 = _GEN_285;
  wire          _GEN_286 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h8;
  wire          compressDataVec_hitReq_26_8;
  assign compressDataVec_hitReq_26_8 = _GEN_286;
  wire          compressDataVec_hitReq_26_136;
  assign compressDataVec_hitReq_26_136 = _GEN_286;
  wire          _GEN_287 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h8;
  wire          compressDataVec_hitReq_27_8;
  assign compressDataVec_hitReq_27_8 = _GEN_287;
  wire          compressDataVec_hitReq_27_136;
  assign compressDataVec_hitReq_27_136 = _GEN_287;
  wire          _GEN_288 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h8;
  wire          compressDataVec_hitReq_28_8;
  assign compressDataVec_hitReq_28_8 = _GEN_288;
  wire          compressDataVec_hitReq_28_136;
  assign compressDataVec_hitReq_28_136 = _GEN_288;
  wire          _GEN_289 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h8;
  wire          compressDataVec_hitReq_29_8;
  assign compressDataVec_hitReq_29_8 = _GEN_289;
  wire          compressDataVec_hitReq_29_136;
  assign compressDataVec_hitReq_29_136 = _GEN_289;
  wire          _GEN_290 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h8;
  wire          compressDataVec_hitReq_30_8;
  assign compressDataVec_hitReq_30_8 = _GEN_290;
  wire          compressDataVec_hitReq_30_136;
  assign compressDataVec_hitReq_30_136 = _GEN_290;
  wire          _GEN_291 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h8;
  wire          compressDataVec_hitReq_31_8;
  assign compressDataVec_hitReq_31_8 = _GEN_291;
  wire          compressDataVec_hitReq_31_136;
  assign compressDataVec_hitReq_31_136 = _GEN_291;
  wire          compressDataVec_hitReq_32_8 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h8;
  wire          compressDataVec_hitReq_33_8 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h8;
  wire          compressDataVec_hitReq_34_8 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h8;
  wire          compressDataVec_hitReq_35_8 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h8;
  wire          compressDataVec_hitReq_36_8 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h8;
  wire          compressDataVec_hitReq_37_8 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h8;
  wire          compressDataVec_hitReq_38_8 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h8;
  wire          compressDataVec_hitReq_39_8 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h8;
  wire          compressDataVec_hitReq_40_8 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h8;
  wire          compressDataVec_hitReq_41_8 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h8;
  wire          compressDataVec_hitReq_42_8 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h8;
  wire          compressDataVec_hitReq_43_8 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h8;
  wire          compressDataVec_hitReq_44_8 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h8;
  wire          compressDataVec_hitReq_45_8 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h8;
  wire          compressDataVec_hitReq_46_8 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h8;
  wire          compressDataVec_hitReq_47_8 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h8;
  wire          compressDataVec_hitReq_48_8 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h8;
  wire          compressDataVec_hitReq_49_8 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h8;
  wire          compressDataVec_hitReq_50_8 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h8;
  wire          compressDataVec_hitReq_51_8 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h8;
  wire          compressDataVec_hitReq_52_8 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h8;
  wire          compressDataVec_hitReq_53_8 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h8;
  wire          compressDataVec_hitReq_54_8 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h8;
  wire          compressDataVec_hitReq_55_8 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h8;
  wire          compressDataVec_hitReq_56_8 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h8;
  wire          compressDataVec_hitReq_57_8 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h8;
  wire          compressDataVec_hitReq_58_8 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h8;
  wire          compressDataVec_hitReq_59_8 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h8;
  wire          compressDataVec_hitReq_60_8 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h8;
  wire          compressDataVec_hitReq_61_8 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h8;
  wire          compressDataVec_hitReq_62_8 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h8;
  wire          compressDataVec_hitReq_63_8 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h8;
  wire [7:0]    compressDataVec_selectReqData_8 =
    (compressDataVec_hitReq_0_8 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_8 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_8 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_8 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_8 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_8 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_8 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_8 ? source2Pipe[63:56] : 8'h0)
    | (compressDataVec_hitReq_8_8 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_8 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_8 ? source2Pipe[87:80] : 8'h0)
    | (compressDataVec_hitReq_11_8 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_8 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_8 ? source2Pipe[111:104] : 8'h0)
    | (compressDataVec_hitReq_14_8 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_8 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_8 ? source2Pipe[135:128] : 8'h0)
    | (compressDataVec_hitReq_17_8 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_8 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_8 ? source2Pipe[159:152] : 8'h0)
    | (compressDataVec_hitReq_20_8 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_8 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_8 ? source2Pipe[183:176] : 8'h0)
    | (compressDataVec_hitReq_23_8 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_8 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_8 ? source2Pipe[207:200] : 8'h0)
    | (compressDataVec_hitReq_26_8 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_8 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_8 ? source2Pipe[231:224] : 8'h0)
    | (compressDataVec_hitReq_29_8 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_8 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_8 ? source2Pipe[255:248] : 8'h0)
    | (compressDataVec_hitReq_32_8 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_8 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_8 ? source2Pipe[279:272] : 8'h0)
    | (compressDataVec_hitReq_35_8 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_8 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_8 ? source2Pipe[303:296] : 8'h0)
    | (compressDataVec_hitReq_38_8 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_8 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_8 ? source2Pipe[327:320] : 8'h0)
    | (compressDataVec_hitReq_41_8 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_8 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_8 ? source2Pipe[351:344] : 8'h0)
    | (compressDataVec_hitReq_44_8 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_8 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_8 ? source2Pipe[375:368] : 8'h0)
    | (compressDataVec_hitReq_47_8 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_8 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_8 ? source2Pipe[399:392] : 8'h0)
    | (compressDataVec_hitReq_50_8 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_8 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_8 ? source2Pipe[423:416] : 8'h0)
    | (compressDataVec_hitReq_53_8 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_8 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_8 ? source2Pipe[447:440] : 8'h0)
    | (compressDataVec_hitReq_56_8 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_8 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_8 ? source2Pipe[471:464] : 8'h0)
    | (compressDataVec_hitReq_59_8 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_8 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_8 ? source2Pipe[495:488] : 8'h0)
    | (compressDataVec_hitReq_62_8 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_8 ? source2Pipe[511:504] : 8'h0);
  wire          _GEN_292 = tailCount > 6'h8;
  wire          compressDataVec_useTail_8;
  assign compressDataVec_useTail_8 = _GEN_292;
  wire          compressDataVec_useTail_72;
  assign compressDataVec_useTail_72 = _GEN_292;
  wire          compressDataVec_useTail_104;
  assign compressDataVec_useTail_104 = _GEN_292;
  wire          _GEN_293 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h9;
  wire          compressDataVec_hitReq_0_9;
  assign compressDataVec_hitReq_0_9 = _GEN_293;
  wire          compressDataVec_hitReq_0_137;
  assign compressDataVec_hitReq_0_137 = _GEN_293;
  wire          compressDataVec_hitReq_0_201;
  assign compressDataVec_hitReq_0_201 = _GEN_293;
  wire          _GEN_294 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h9;
  wire          compressDataVec_hitReq_1_9;
  assign compressDataVec_hitReq_1_9 = _GEN_294;
  wire          compressDataVec_hitReq_1_137;
  assign compressDataVec_hitReq_1_137 = _GEN_294;
  wire          compressDataVec_hitReq_1_201;
  assign compressDataVec_hitReq_1_201 = _GEN_294;
  wire          _GEN_295 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h9;
  wire          compressDataVec_hitReq_2_9;
  assign compressDataVec_hitReq_2_9 = _GEN_295;
  wire          compressDataVec_hitReq_2_137;
  assign compressDataVec_hitReq_2_137 = _GEN_295;
  wire          compressDataVec_hitReq_2_201;
  assign compressDataVec_hitReq_2_201 = _GEN_295;
  wire          _GEN_296 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h9;
  wire          compressDataVec_hitReq_3_9;
  assign compressDataVec_hitReq_3_9 = _GEN_296;
  wire          compressDataVec_hitReq_3_137;
  assign compressDataVec_hitReq_3_137 = _GEN_296;
  wire          compressDataVec_hitReq_3_201;
  assign compressDataVec_hitReq_3_201 = _GEN_296;
  wire          _GEN_297 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h9;
  wire          compressDataVec_hitReq_4_9;
  assign compressDataVec_hitReq_4_9 = _GEN_297;
  wire          compressDataVec_hitReq_4_137;
  assign compressDataVec_hitReq_4_137 = _GEN_297;
  wire          compressDataVec_hitReq_4_201;
  assign compressDataVec_hitReq_4_201 = _GEN_297;
  wire          _GEN_298 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h9;
  wire          compressDataVec_hitReq_5_9;
  assign compressDataVec_hitReq_5_9 = _GEN_298;
  wire          compressDataVec_hitReq_5_137;
  assign compressDataVec_hitReq_5_137 = _GEN_298;
  wire          compressDataVec_hitReq_5_201;
  assign compressDataVec_hitReq_5_201 = _GEN_298;
  wire          _GEN_299 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h9;
  wire          compressDataVec_hitReq_6_9;
  assign compressDataVec_hitReq_6_9 = _GEN_299;
  wire          compressDataVec_hitReq_6_137;
  assign compressDataVec_hitReq_6_137 = _GEN_299;
  wire          compressDataVec_hitReq_6_201;
  assign compressDataVec_hitReq_6_201 = _GEN_299;
  wire          _GEN_300 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h9;
  wire          compressDataVec_hitReq_7_9;
  assign compressDataVec_hitReq_7_9 = _GEN_300;
  wire          compressDataVec_hitReq_7_137;
  assign compressDataVec_hitReq_7_137 = _GEN_300;
  wire          compressDataVec_hitReq_7_201;
  assign compressDataVec_hitReq_7_201 = _GEN_300;
  wire          _GEN_301 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h9;
  wire          compressDataVec_hitReq_8_9;
  assign compressDataVec_hitReq_8_9 = _GEN_301;
  wire          compressDataVec_hitReq_8_137;
  assign compressDataVec_hitReq_8_137 = _GEN_301;
  wire          compressDataVec_hitReq_8_201;
  assign compressDataVec_hitReq_8_201 = _GEN_301;
  wire          _GEN_302 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h9;
  wire          compressDataVec_hitReq_9_9;
  assign compressDataVec_hitReq_9_9 = _GEN_302;
  wire          compressDataVec_hitReq_9_137;
  assign compressDataVec_hitReq_9_137 = _GEN_302;
  wire          compressDataVec_hitReq_9_201;
  assign compressDataVec_hitReq_9_201 = _GEN_302;
  wire          _GEN_303 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h9;
  wire          compressDataVec_hitReq_10_9;
  assign compressDataVec_hitReq_10_9 = _GEN_303;
  wire          compressDataVec_hitReq_10_137;
  assign compressDataVec_hitReq_10_137 = _GEN_303;
  wire          compressDataVec_hitReq_10_201;
  assign compressDataVec_hitReq_10_201 = _GEN_303;
  wire          _GEN_304 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h9;
  wire          compressDataVec_hitReq_11_9;
  assign compressDataVec_hitReq_11_9 = _GEN_304;
  wire          compressDataVec_hitReq_11_137;
  assign compressDataVec_hitReq_11_137 = _GEN_304;
  wire          compressDataVec_hitReq_11_201;
  assign compressDataVec_hitReq_11_201 = _GEN_304;
  wire          _GEN_305 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h9;
  wire          compressDataVec_hitReq_12_9;
  assign compressDataVec_hitReq_12_9 = _GEN_305;
  wire          compressDataVec_hitReq_12_137;
  assign compressDataVec_hitReq_12_137 = _GEN_305;
  wire          compressDataVec_hitReq_12_201;
  assign compressDataVec_hitReq_12_201 = _GEN_305;
  wire          _GEN_306 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h9;
  wire          compressDataVec_hitReq_13_9;
  assign compressDataVec_hitReq_13_9 = _GEN_306;
  wire          compressDataVec_hitReq_13_137;
  assign compressDataVec_hitReq_13_137 = _GEN_306;
  wire          compressDataVec_hitReq_13_201;
  assign compressDataVec_hitReq_13_201 = _GEN_306;
  wire          _GEN_307 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h9;
  wire          compressDataVec_hitReq_14_9;
  assign compressDataVec_hitReq_14_9 = _GEN_307;
  wire          compressDataVec_hitReq_14_137;
  assign compressDataVec_hitReq_14_137 = _GEN_307;
  wire          compressDataVec_hitReq_14_201;
  assign compressDataVec_hitReq_14_201 = _GEN_307;
  wire          _GEN_308 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h9;
  wire          compressDataVec_hitReq_15_9;
  assign compressDataVec_hitReq_15_9 = _GEN_308;
  wire          compressDataVec_hitReq_15_137;
  assign compressDataVec_hitReq_15_137 = _GEN_308;
  wire          compressDataVec_hitReq_15_201;
  assign compressDataVec_hitReq_15_201 = _GEN_308;
  wire          _GEN_309 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h9;
  wire          compressDataVec_hitReq_16_9;
  assign compressDataVec_hitReq_16_9 = _GEN_309;
  wire          compressDataVec_hitReq_16_137;
  assign compressDataVec_hitReq_16_137 = _GEN_309;
  wire          _GEN_310 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h9;
  wire          compressDataVec_hitReq_17_9;
  assign compressDataVec_hitReq_17_9 = _GEN_310;
  wire          compressDataVec_hitReq_17_137;
  assign compressDataVec_hitReq_17_137 = _GEN_310;
  wire          _GEN_311 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h9;
  wire          compressDataVec_hitReq_18_9;
  assign compressDataVec_hitReq_18_9 = _GEN_311;
  wire          compressDataVec_hitReq_18_137;
  assign compressDataVec_hitReq_18_137 = _GEN_311;
  wire          _GEN_312 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h9;
  wire          compressDataVec_hitReq_19_9;
  assign compressDataVec_hitReq_19_9 = _GEN_312;
  wire          compressDataVec_hitReq_19_137;
  assign compressDataVec_hitReq_19_137 = _GEN_312;
  wire          _GEN_313 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h9;
  wire          compressDataVec_hitReq_20_9;
  assign compressDataVec_hitReq_20_9 = _GEN_313;
  wire          compressDataVec_hitReq_20_137;
  assign compressDataVec_hitReq_20_137 = _GEN_313;
  wire          _GEN_314 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h9;
  wire          compressDataVec_hitReq_21_9;
  assign compressDataVec_hitReq_21_9 = _GEN_314;
  wire          compressDataVec_hitReq_21_137;
  assign compressDataVec_hitReq_21_137 = _GEN_314;
  wire          _GEN_315 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h9;
  wire          compressDataVec_hitReq_22_9;
  assign compressDataVec_hitReq_22_9 = _GEN_315;
  wire          compressDataVec_hitReq_22_137;
  assign compressDataVec_hitReq_22_137 = _GEN_315;
  wire          _GEN_316 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h9;
  wire          compressDataVec_hitReq_23_9;
  assign compressDataVec_hitReq_23_9 = _GEN_316;
  wire          compressDataVec_hitReq_23_137;
  assign compressDataVec_hitReq_23_137 = _GEN_316;
  wire          _GEN_317 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h9;
  wire          compressDataVec_hitReq_24_9;
  assign compressDataVec_hitReq_24_9 = _GEN_317;
  wire          compressDataVec_hitReq_24_137;
  assign compressDataVec_hitReq_24_137 = _GEN_317;
  wire          _GEN_318 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h9;
  wire          compressDataVec_hitReq_25_9;
  assign compressDataVec_hitReq_25_9 = _GEN_318;
  wire          compressDataVec_hitReq_25_137;
  assign compressDataVec_hitReq_25_137 = _GEN_318;
  wire          _GEN_319 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h9;
  wire          compressDataVec_hitReq_26_9;
  assign compressDataVec_hitReq_26_9 = _GEN_319;
  wire          compressDataVec_hitReq_26_137;
  assign compressDataVec_hitReq_26_137 = _GEN_319;
  wire          _GEN_320 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h9;
  wire          compressDataVec_hitReq_27_9;
  assign compressDataVec_hitReq_27_9 = _GEN_320;
  wire          compressDataVec_hitReq_27_137;
  assign compressDataVec_hitReq_27_137 = _GEN_320;
  wire          _GEN_321 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h9;
  wire          compressDataVec_hitReq_28_9;
  assign compressDataVec_hitReq_28_9 = _GEN_321;
  wire          compressDataVec_hitReq_28_137;
  assign compressDataVec_hitReq_28_137 = _GEN_321;
  wire          _GEN_322 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h9;
  wire          compressDataVec_hitReq_29_9;
  assign compressDataVec_hitReq_29_9 = _GEN_322;
  wire          compressDataVec_hitReq_29_137;
  assign compressDataVec_hitReq_29_137 = _GEN_322;
  wire          _GEN_323 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h9;
  wire          compressDataVec_hitReq_30_9;
  assign compressDataVec_hitReq_30_9 = _GEN_323;
  wire          compressDataVec_hitReq_30_137;
  assign compressDataVec_hitReq_30_137 = _GEN_323;
  wire          _GEN_324 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h9;
  wire          compressDataVec_hitReq_31_9;
  assign compressDataVec_hitReq_31_9 = _GEN_324;
  wire          compressDataVec_hitReq_31_137;
  assign compressDataVec_hitReq_31_137 = _GEN_324;
  wire          compressDataVec_hitReq_32_9 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h9;
  wire          compressDataVec_hitReq_33_9 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h9;
  wire          compressDataVec_hitReq_34_9 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h9;
  wire          compressDataVec_hitReq_35_9 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h9;
  wire          compressDataVec_hitReq_36_9 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h9;
  wire          compressDataVec_hitReq_37_9 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h9;
  wire          compressDataVec_hitReq_38_9 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h9;
  wire          compressDataVec_hitReq_39_9 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h9;
  wire          compressDataVec_hitReq_40_9 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h9;
  wire          compressDataVec_hitReq_41_9 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h9;
  wire          compressDataVec_hitReq_42_9 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h9;
  wire          compressDataVec_hitReq_43_9 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h9;
  wire          compressDataVec_hitReq_44_9 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h9;
  wire          compressDataVec_hitReq_45_9 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h9;
  wire          compressDataVec_hitReq_46_9 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h9;
  wire          compressDataVec_hitReq_47_9 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h9;
  wire          compressDataVec_hitReq_48_9 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h9;
  wire          compressDataVec_hitReq_49_9 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h9;
  wire          compressDataVec_hitReq_50_9 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h9;
  wire          compressDataVec_hitReq_51_9 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h9;
  wire          compressDataVec_hitReq_52_9 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h9;
  wire          compressDataVec_hitReq_53_9 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h9;
  wire          compressDataVec_hitReq_54_9 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h9;
  wire          compressDataVec_hitReq_55_9 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h9;
  wire          compressDataVec_hitReq_56_9 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h9;
  wire          compressDataVec_hitReq_57_9 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h9;
  wire          compressDataVec_hitReq_58_9 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h9;
  wire          compressDataVec_hitReq_59_9 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h9;
  wire          compressDataVec_hitReq_60_9 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h9;
  wire          compressDataVec_hitReq_61_9 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h9;
  wire          compressDataVec_hitReq_62_9 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h9;
  wire          compressDataVec_hitReq_63_9 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h9;
  wire [7:0]    compressDataVec_selectReqData_9 =
    (compressDataVec_hitReq_0_9 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_9 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_9 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_9 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_9 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_9 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_9 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_9 ? source2Pipe[63:56] : 8'h0)
    | (compressDataVec_hitReq_8_9 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_9 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_9 ? source2Pipe[87:80] : 8'h0)
    | (compressDataVec_hitReq_11_9 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_9 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_9 ? source2Pipe[111:104] : 8'h0)
    | (compressDataVec_hitReq_14_9 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_9 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_9 ? source2Pipe[135:128] : 8'h0)
    | (compressDataVec_hitReq_17_9 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_9 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_9 ? source2Pipe[159:152] : 8'h0)
    | (compressDataVec_hitReq_20_9 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_9 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_9 ? source2Pipe[183:176] : 8'h0)
    | (compressDataVec_hitReq_23_9 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_9 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_9 ? source2Pipe[207:200] : 8'h0)
    | (compressDataVec_hitReq_26_9 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_9 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_9 ? source2Pipe[231:224] : 8'h0)
    | (compressDataVec_hitReq_29_9 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_9 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_9 ? source2Pipe[255:248] : 8'h0)
    | (compressDataVec_hitReq_32_9 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_9 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_9 ? source2Pipe[279:272] : 8'h0)
    | (compressDataVec_hitReq_35_9 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_9 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_9 ? source2Pipe[303:296] : 8'h0)
    | (compressDataVec_hitReq_38_9 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_9 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_9 ? source2Pipe[327:320] : 8'h0)
    | (compressDataVec_hitReq_41_9 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_9 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_9 ? source2Pipe[351:344] : 8'h0)
    | (compressDataVec_hitReq_44_9 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_9 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_9 ? source2Pipe[375:368] : 8'h0)
    | (compressDataVec_hitReq_47_9 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_9 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_9 ? source2Pipe[399:392] : 8'h0)
    | (compressDataVec_hitReq_50_9 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_9 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_9 ? source2Pipe[423:416] : 8'h0)
    | (compressDataVec_hitReq_53_9 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_9 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_9 ? source2Pipe[447:440] : 8'h0)
    | (compressDataVec_hitReq_56_9 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_9 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_9 ? source2Pipe[471:464] : 8'h0)
    | (compressDataVec_hitReq_59_9 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_9 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_9 ? source2Pipe[495:488] : 8'h0)
    | (compressDataVec_hitReq_62_9 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_9 ? source2Pipe[511:504] : 8'h0);
  wire          _GEN_325 = tailCount > 6'h9;
  wire          compressDataVec_useTail_9;
  assign compressDataVec_useTail_9 = _GEN_325;
  wire          compressDataVec_useTail_73;
  assign compressDataVec_useTail_73 = _GEN_325;
  wire          compressDataVec_useTail_105;
  assign compressDataVec_useTail_105 = _GEN_325;
  wire          _GEN_326 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'hA;
  wire          compressDataVec_hitReq_0_10;
  assign compressDataVec_hitReq_0_10 = _GEN_326;
  wire          compressDataVec_hitReq_0_138;
  assign compressDataVec_hitReq_0_138 = _GEN_326;
  wire          compressDataVec_hitReq_0_202;
  assign compressDataVec_hitReq_0_202 = _GEN_326;
  wire          _GEN_327 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'hA;
  wire          compressDataVec_hitReq_1_10;
  assign compressDataVec_hitReq_1_10 = _GEN_327;
  wire          compressDataVec_hitReq_1_138;
  assign compressDataVec_hitReq_1_138 = _GEN_327;
  wire          compressDataVec_hitReq_1_202;
  assign compressDataVec_hitReq_1_202 = _GEN_327;
  wire          _GEN_328 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'hA;
  wire          compressDataVec_hitReq_2_10;
  assign compressDataVec_hitReq_2_10 = _GEN_328;
  wire          compressDataVec_hitReq_2_138;
  assign compressDataVec_hitReq_2_138 = _GEN_328;
  wire          compressDataVec_hitReq_2_202;
  assign compressDataVec_hitReq_2_202 = _GEN_328;
  wire          _GEN_329 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'hA;
  wire          compressDataVec_hitReq_3_10;
  assign compressDataVec_hitReq_3_10 = _GEN_329;
  wire          compressDataVec_hitReq_3_138;
  assign compressDataVec_hitReq_3_138 = _GEN_329;
  wire          compressDataVec_hitReq_3_202;
  assign compressDataVec_hitReq_3_202 = _GEN_329;
  wire          _GEN_330 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'hA;
  wire          compressDataVec_hitReq_4_10;
  assign compressDataVec_hitReq_4_10 = _GEN_330;
  wire          compressDataVec_hitReq_4_138;
  assign compressDataVec_hitReq_4_138 = _GEN_330;
  wire          compressDataVec_hitReq_4_202;
  assign compressDataVec_hitReq_4_202 = _GEN_330;
  wire          _GEN_331 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'hA;
  wire          compressDataVec_hitReq_5_10;
  assign compressDataVec_hitReq_5_10 = _GEN_331;
  wire          compressDataVec_hitReq_5_138;
  assign compressDataVec_hitReq_5_138 = _GEN_331;
  wire          compressDataVec_hitReq_5_202;
  assign compressDataVec_hitReq_5_202 = _GEN_331;
  wire          _GEN_332 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'hA;
  wire          compressDataVec_hitReq_6_10;
  assign compressDataVec_hitReq_6_10 = _GEN_332;
  wire          compressDataVec_hitReq_6_138;
  assign compressDataVec_hitReq_6_138 = _GEN_332;
  wire          compressDataVec_hitReq_6_202;
  assign compressDataVec_hitReq_6_202 = _GEN_332;
  wire          _GEN_333 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'hA;
  wire          compressDataVec_hitReq_7_10;
  assign compressDataVec_hitReq_7_10 = _GEN_333;
  wire          compressDataVec_hitReq_7_138;
  assign compressDataVec_hitReq_7_138 = _GEN_333;
  wire          compressDataVec_hitReq_7_202;
  assign compressDataVec_hitReq_7_202 = _GEN_333;
  wire          _GEN_334 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'hA;
  wire          compressDataVec_hitReq_8_10;
  assign compressDataVec_hitReq_8_10 = _GEN_334;
  wire          compressDataVec_hitReq_8_138;
  assign compressDataVec_hitReq_8_138 = _GEN_334;
  wire          compressDataVec_hitReq_8_202;
  assign compressDataVec_hitReq_8_202 = _GEN_334;
  wire          _GEN_335 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'hA;
  wire          compressDataVec_hitReq_9_10;
  assign compressDataVec_hitReq_9_10 = _GEN_335;
  wire          compressDataVec_hitReq_9_138;
  assign compressDataVec_hitReq_9_138 = _GEN_335;
  wire          compressDataVec_hitReq_9_202;
  assign compressDataVec_hitReq_9_202 = _GEN_335;
  wire          _GEN_336 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'hA;
  wire          compressDataVec_hitReq_10_10;
  assign compressDataVec_hitReq_10_10 = _GEN_336;
  wire          compressDataVec_hitReq_10_138;
  assign compressDataVec_hitReq_10_138 = _GEN_336;
  wire          compressDataVec_hitReq_10_202;
  assign compressDataVec_hitReq_10_202 = _GEN_336;
  wire          _GEN_337 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'hA;
  wire          compressDataVec_hitReq_11_10;
  assign compressDataVec_hitReq_11_10 = _GEN_337;
  wire          compressDataVec_hitReq_11_138;
  assign compressDataVec_hitReq_11_138 = _GEN_337;
  wire          compressDataVec_hitReq_11_202;
  assign compressDataVec_hitReq_11_202 = _GEN_337;
  wire          _GEN_338 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'hA;
  wire          compressDataVec_hitReq_12_10;
  assign compressDataVec_hitReq_12_10 = _GEN_338;
  wire          compressDataVec_hitReq_12_138;
  assign compressDataVec_hitReq_12_138 = _GEN_338;
  wire          compressDataVec_hitReq_12_202;
  assign compressDataVec_hitReq_12_202 = _GEN_338;
  wire          _GEN_339 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'hA;
  wire          compressDataVec_hitReq_13_10;
  assign compressDataVec_hitReq_13_10 = _GEN_339;
  wire          compressDataVec_hitReq_13_138;
  assign compressDataVec_hitReq_13_138 = _GEN_339;
  wire          compressDataVec_hitReq_13_202;
  assign compressDataVec_hitReq_13_202 = _GEN_339;
  wire          _GEN_340 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'hA;
  wire          compressDataVec_hitReq_14_10;
  assign compressDataVec_hitReq_14_10 = _GEN_340;
  wire          compressDataVec_hitReq_14_138;
  assign compressDataVec_hitReq_14_138 = _GEN_340;
  wire          compressDataVec_hitReq_14_202;
  assign compressDataVec_hitReq_14_202 = _GEN_340;
  wire          _GEN_341 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'hA;
  wire          compressDataVec_hitReq_15_10;
  assign compressDataVec_hitReq_15_10 = _GEN_341;
  wire          compressDataVec_hitReq_15_138;
  assign compressDataVec_hitReq_15_138 = _GEN_341;
  wire          compressDataVec_hitReq_15_202;
  assign compressDataVec_hitReq_15_202 = _GEN_341;
  wire          _GEN_342 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'hA;
  wire          compressDataVec_hitReq_16_10;
  assign compressDataVec_hitReq_16_10 = _GEN_342;
  wire          compressDataVec_hitReq_16_138;
  assign compressDataVec_hitReq_16_138 = _GEN_342;
  wire          _GEN_343 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'hA;
  wire          compressDataVec_hitReq_17_10;
  assign compressDataVec_hitReq_17_10 = _GEN_343;
  wire          compressDataVec_hitReq_17_138;
  assign compressDataVec_hitReq_17_138 = _GEN_343;
  wire          _GEN_344 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'hA;
  wire          compressDataVec_hitReq_18_10;
  assign compressDataVec_hitReq_18_10 = _GEN_344;
  wire          compressDataVec_hitReq_18_138;
  assign compressDataVec_hitReq_18_138 = _GEN_344;
  wire          _GEN_345 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'hA;
  wire          compressDataVec_hitReq_19_10;
  assign compressDataVec_hitReq_19_10 = _GEN_345;
  wire          compressDataVec_hitReq_19_138;
  assign compressDataVec_hitReq_19_138 = _GEN_345;
  wire          _GEN_346 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'hA;
  wire          compressDataVec_hitReq_20_10;
  assign compressDataVec_hitReq_20_10 = _GEN_346;
  wire          compressDataVec_hitReq_20_138;
  assign compressDataVec_hitReq_20_138 = _GEN_346;
  wire          _GEN_347 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'hA;
  wire          compressDataVec_hitReq_21_10;
  assign compressDataVec_hitReq_21_10 = _GEN_347;
  wire          compressDataVec_hitReq_21_138;
  assign compressDataVec_hitReq_21_138 = _GEN_347;
  wire          _GEN_348 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'hA;
  wire          compressDataVec_hitReq_22_10;
  assign compressDataVec_hitReq_22_10 = _GEN_348;
  wire          compressDataVec_hitReq_22_138;
  assign compressDataVec_hitReq_22_138 = _GEN_348;
  wire          _GEN_349 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'hA;
  wire          compressDataVec_hitReq_23_10;
  assign compressDataVec_hitReq_23_10 = _GEN_349;
  wire          compressDataVec_hitReq_23_138;
  assign compressDataVec_hitReq_23_138 = _GEN_349;
  wire          _GEN_350 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'hA;
  wire          compressDataVec_hitReq_24_10;
  assign compressDataVec_hitReq_24_10 = _GEN_350;
  wire          compressDataVec_hitReq_24_138;
  assign compressDataVec_hitReq_24_138 = _GEN_350;
  wire          _GEN_351 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'hA;
  wire          compressDataVec_hitReq_25_10;
  assign compressDataVec_hitReq_25_10 = _GEN_351;
  wire          compressDataVec_hitReq_25_138;
  assign compressDataVec_hitReq_25_138 = _GEN_351;
  wire          _GEN_352 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'hA;
  wire          compressDataVec_hitReq_26_10;
  assign compressDataVec_hitReq_26_10 = _GEN_352;
  wire          compressDataVec_hitReq_26_138;
  assign compressDataVec_hitReq_26_138 = _GEN_352;
  wire          _GEN_353 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'hA;
  wire          compressDataVec_hitReq_27_10;
  assign compressDataVec_hitReq_27_10 = _GEN_353;
  wire          compressDataVec_hitReq_27_138;
  assign compressDataVec_hitReq_27_138 = _GEN_353;
  wire          _GEN_354 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'hA;
  wire          compressDataVec_hitReq_28_10;
  assign compressDataVec_hitReq_28_10 = _GEN_354;
  wire          compressDataVec_hitReq_28_138;
  assign compressDataVec_hitReq_28_138 = _GEN_354;
  wire          _GEN_355 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'hA;
  wire          compressDataVec_hitReq_29_10;
  assign compressDataVec_hitReq_29_10 = _GEN_355;
  wire          compressDataVec_hitReq_29_138;
  assign compressDataVec_hitReq_29_138 = _GEN_355;
  wire          _GEN_356 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'hA;
  wire          compressDataVec_hitReq_30_10;
  assign compressDataVec_hitReq_30_10 = _GEN_356;
  wire          compressDataVec_hitReq_30_138;
  assign compressDataVec_hitReq_30_138 = _GEN_356;
  wire          _GEN_357 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'hA;
  wire          compressDataVec_hitReq_31_10;
  assign compressDataVec_hitReq_31_10 = _GEN_357;
  wire          compressDataVec_hitReq_31_138;
  assign compressDataVec_hitReq_31_138 = _GEN_357;
  wire          compressDataVec_hitReq_32_10 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'hA;
  wire          compressDataVec_hitReq_33_10 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'hA;
  wire          compressDataVec_hitReq_34_10 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'hA;
  wire          compressDataVec_hitReq_35_10 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'hA;
  wire          compressDataVec_hitReq_36_10 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'hA;
  wire          compressDataVec_hitReq_37_10 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'hA;
  wire          compressDataVec_hitReq_38_10 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'hA;
  wire          compressDataVec_hitReq_39_10 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'hA;
  wire          compressDataVec_hitReq_40_10 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'hA;
  wire          compressDataVec_hitReq_41_10 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'hA;
  wire          compressDataVec_hitReq_42_10 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'hA;
  wire          compressDataVec_hitReq_43_10 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'hA;
  wire          compressDataVec_hitReq_44_10 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'hA;
  wire          compressDataVec_hitReq_45_10 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'hA;
  wire          compressDataVec_hitReq_46_10 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'hA;
  wire          compressDataVec_hitReq_47_10 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'hA;
  wire          compressDataVec_hitReq_48_10 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'hA;
  wire          compressDataVec_hitReq_49_10 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'hA;
  wire          compressDataVec_hitReq_50_10 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'hA;
  wire          compressDataVec_hitReq_51_10 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'hA;
  wire          compressDataVec_hitReq_52_10 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'hA;
  wire          compressDataVec_hitReq_53_10 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'hA;
  wire          compressDataVec_hitReq_54_10 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'hA;
  wire          compressDataVec_hitReq_55_10 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'hA;
  wire          compressDataVec_hitReq_56_10 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'hA;
  wire          compressDataVec_hitReq_57_10 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'hA;
  wire          compressDataVec_hitReq_58_10 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'hA;
  wire          compressDataVec_hitReq_59_10 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'hA;
  wire          compressDataVec_hitReq_60_10 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'hA;
  wire          compressDataVec_hitReq_61_10 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'hA;
  wire          compressDataVec_hitReq_62_10 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'hA;
  wire          compressDataVec_hitReq_63_10 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'hA;
  wire [7:0]    compressDataVec_selectReqData_10 =
    (compressDataVec_hitReq_0_10 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_10 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_10 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_10 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_10 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_10 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_10 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_10 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_10 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_10 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_10 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_10 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_10 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_10 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_10 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_10 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_10 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_10 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_10 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_10 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_10 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_10 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_10 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_10 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_10 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_10 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_10 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_10 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_10 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_10 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_10 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_10 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_10 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_10 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_10 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_10 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_10 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_10 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_10 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_10 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_10 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_10 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_10 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_10 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_10 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_10 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_10 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_10 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_10 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_10 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_10 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_10 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_10 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_10 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_10 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_10 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_10 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_10 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_10 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_10 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_10 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_10 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_10 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_10 ? source2Pipe[511:504] : 8'h0);
  wire          _GEN_358 = tailCount > 6'hA;
  wire          compressDataVec_useTail_10;
  assign compressDataVec_useTail_10 = _GEN_358;
  wire          compressDataVec_useTail_74;
  assign compressDataVec_useTail_74 = _GEN_358;
  wire          compressDataVec_useTail_106;
  assign compressDataVec_useTail_106 = _GEN_358;
  wire          _GEN_359 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'hB;
  wire          compressDataVec_hitReq_0_11;
  assign compressDataVec_hitReq_0_11 = _GEN_359;
  wire          compressDataVec_hitReq_0_139;
  assign compressDataVec_hitReq_0_139 = _GEN_359;
  wire          compressDataVec_hitReq_0_203;
  assign compressDataVec_hitReq_0_203 = _GEN_359;
  wire          _GEN_360 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'hB;
  wire          compressDataVec_hitReq_1_11;
  assign compressDataVec_hitReq_1_11 = _GEN_360;
  wire          compressDataVec_hitReq_1_139;
  assign compressDataVec_hitReq_1_139 = _GEN_360;
  wire          compressDataVec_hitReq_1_203;
  assign compressDataVec_hitReq_1_203 = _GEN_360;
  wire          _GEN_361 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'hB;
  wire          compressDataVec_hitReq_2_11;
  assign compressDataVec_hitReq_2_11 = _GEN_361;
  wire          compressDataVec_hitReq_2_139;
  assign compressDataVec_hitReq_2_139 = _GEN_361;
  wire          compressDataVec_hitReq_2_203;
  assign compressDataVec_hitReq_2_203 = _GEN_361;
  wire          _GEN_362 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'hB;
  wire          compressDataVec_hitReq_3_11;
  assign compressDataVec_hitReq_3_11 = _GEN_362;
  wire          compressDataVec_hitReq_3_139;
  assign compressDataVec_hitReq_3_139 = _GEN_362;
  wire          compressDataVec_hitReq_3_203;
  assign compressDataVec_hitReq_3_203 = _GEN_362;
  wire          _GEN_363 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'hB;
  wire          compressDataVec_hitReq_4_11;
  assign compressDataVec_hitReq_4_11 = _GEN_363;
  wire          compressDataVec_hitReq_4_139;
  assign compressDataVec_hitReq_4_139 = _GEN_363;
  wire          compressDataVec_hitReq_4_203;
  assign compressDataVec_hitReq_4_203 = _GEN_363;
  wire          _GEN_364 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'hB;
  wire          compressDataVec_hitReq_5_11;
  assign compressDataVec_hitReq_5_11 = _GEN_364;
  wire          compressDataVec_hitReq_5_139;
  assign compressDataVec_hitReq_5_139 = _GEN_364;
  wire          compressDataVec_hitReq_5_203;
  assign compressDataVec_hitReq_5_203 = _GEN_364;
  wire          _GEN_365 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'hB;
  wire          compressDataVec_hitReq_6_11;
  assign compressDataVec_hitReq_6_11 = _GEN_365;
  wire          compressDataVec_hitReq_6_139;
  assign compressDataVec_hitReq_6_139 = _GEN_365;
  wire          compressDataVec_hitReq_6_203;
  assign compressDataVec_hitReq_6_203 = _GEN_365;
  wire          _GEN_366 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'hB;
  wire          compressDataVec_hitReq_7_11;
  assign compressDataVec_hitReq_7_11 = _GEN_366;
  wire          compressDataVec_hitReq_7_139;
  assign compressDataVec_hitReq_7_139 = _GEN_366;
  wire          compressDataVec_hitReq_7_203;
  assign compressDataVec_hitReq_7_203 = _GEN_366;
  wire          _GEN_367 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'hB;
  wire          compressDataVec_hitReq_8_11;
  assign compressDataVec_hitReq_8_11 = _GEN_367;
  wire          compressDataVec_hitReq_8_139;
  assign compressDataVec_hitReq_8_139 = _GEN_367;
  wire          compressDataVec_hitReq_8_203;
  assign compressDataVec_hitReq_8_203 = _GEN_367;
  wire          _GEN_368 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'hB;
  wire          compressDataVec_hitReq_9_11;
  assign compressDataVec_hitReq_9_11 = _GEN_368;
  wire          compressDataVec_hitReq_9_139;
  assign compressDataVec_hitReq_9_139 = _GEN_368;
  wire          compressDataVec_hitReq_9_203;
  assign compressDataVec_hitReq_9_203 = _GEN_368;
  wire          _GEN_369 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'hB;
  wire          compressDataVec_hitReq_10_11;
  assign compressDataVec_hitReq_10_11 = _GEN_369;
  wire          compressDataVec_hitReq_10_139;
  assign compressDataVec_hitReq_10_139 = _GEN_369;
  wire          compressDataVec_hitReq_10_203;
  assign compressDataVec_hitReq_10_203 = _GEN_369;
  wire          _GEN_370 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'hB;
  wire          compressDataVec_hitReq_11_11;
  assign compressDataVec_hitReq_11_11 = _GEN_370;
  wire          compressDataVec_hitReq_11_139;
  assign compressDataVec_hitReq_11_139 = _GEN_370;
  wire          compressDataVec_hitReq_11_203;
  assign compressDataVec_hitReq_11_203 = _GEN_370;
  wire          _GEN_371 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'hB;
  wire          compressDataVec_hitReq_12_11;
  assign compressDataVec_hitReq_12_11 = _GEN_371;
  wire          compressDataVec_hitReq_12_139;
  assign compressDataVec_hitReq_12_139 = _GEN_371;
  wire          compressDataVec_hitReq_12_203;
  assign compressDataVec_hitReq_12_203 = _GEN_371;
  wire          _GEN_372 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'hB;
  wire          compressDataVec_hitReq_13_11;
  assign compressDataVec_hitReq_13_11 = _GEN_372;
  wire          compressDataVec_hitReq_13_139;
  assign compressDataVec_hitReq_13_139 = _GEN_372;
  wire          compressDataVec_hitReq_13_203;
  assign compressDataVec_hitReq_13_203 = _GEN_372;
  wire          _GEN_373 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'hB;
  wire          compressDataVec_hitReq_14_11;
  assign compressDataVec_hitReq_14_11 = _GEN_373;
  wire          compressDataVec_hitReq_14_139;
  assign compressDataVec_hitReq_14_139 = _GEN_373;
  wire          compressDataVec_hitReq_14_203;
  assign compressDataVec_hitReq_14_203 = _GEN_373;
  wire          _GEN_374 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'hB;
  wire          compressDataVec_hitReq_15_11;
  assign compressDataVec_hitReq_15_11 = _GEN_374;
  wire          compressDataVec_hitReq_15_139;
  assign compressDataVec_hitReq_15_139 = _GEN_374;
  wire          compressDataVec_hitReq_15_203;
  assign compressDataVec_hitReq_15_203 = _GEN_374;
  wire          _GEN_375 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'hB;
  wire          compressDataVec_hitReq_16_11;
  assign compressDataVec_hitReq_16_11 = _GEN_375;
  wire          compressDataVec_hitReq_16_139;
  assign compressDataVec_hitReq_16_139 = _GEN_375;
  wire          _GEN_376 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'hB;
  wire          compressDataVec_hitReq_17_11;
  assign compressDataVec_hitReq_17_11 = _GEN_376;
  wire          compressDataVec_hitReq_17_139;
  assign compressDataVec_hitReq_17_139 = _GEN_376;
  wire          _GEN_377 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'hB;
  wire          compressDataVec_hitReq_18_11;
  assign compressDataVec_hitReq_18_11 = _GEN_377;
  wire          compressDataVec_hitReq_18_139;
  assign compressDataVec_hitReq_18_139 = _GEN_377;
  wire          _GEN_378 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'hB;
  wire          compressDataVec_hitReq_19_11;
  assign compressDataVec_hitReq_19_11 = _GEN_378;
  wire          compressDataVec_hitReq_19_139;
  assign compressDataVec_hitReq_19_139 = _GEN_378;
  wire          _GEN_379 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'hB;
  wire          compressDataVec_hitReq_20_11;
  assign compressDataVec_hitReq_20_11 = _GEN_379;
  wire          compressDataVec_hitReq_20_139;
  assign compressDataVec_hitReq_20_139 = _GEN_379;
  wire          _GEN_380 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'hB;
  wire          compressDataVec_hitReq_21_11;
  assign compressDataVec_hitReq_21_11 = _GEN_380;
  wire          compressDataVec_hitReq_21_139;
  assign compressDataVec_hitReq_21_139 = _GEN_380;
  wire          _GEN_381 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'hB;
  wire          compressDataVec_hitReq_22_11;
  assign compressDataVec_hitReq_22_11 = _GEN_381;
  wire          compressDataVec_hitReq_22_139;
  assign compressDataVec_hitReq_22_139 = _GEN_381;
  wire          _GEN_382 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'hB;
  wire          compressDataVec_hitReq_23_11;
  assign compressDataVec_hitReq_23_11 = _GEN_382;
  wire          compressDataVec_hitReq_23_139;
  assign compressDataVec_hitReq_23_139 = _GEN_382;
  wire          _GEN_383 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'hB;
  wire          compressDataVec_hitReq_24_11;
  assign compressDataVec_hitReq_24_11 = _GEN_383;
  wire          compressDataVec_hitReq_24_139;
  assign compressDataVec_hitReq_24_139 = _GEN_383;
  wire          _GEN_384 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'hB;
  wire          compressDataVec_hitReq_25_11;
  assign compressDataVec_hitReq_25_11 = _GEN_384;
  wire          compressDataVec_hitReq_25_139;
  assign compressDataVec_hitReq_25_139 = _GEN_384;
  wire          _GEN_385 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'hB;
  wire          compressDataVec_hitReq_26_11;
  assign compressDataVec_hitReq_26_11 = _GEN_385;
  wire          compressDataVec_hitReq_26_139;
  assign compressDataVec_hitReq_26_139 = _GEN_385;
  wire          _GEN_386 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'hB;
  wire          compressDataVec_hitReq_27_11;
  assign compressDataVec_hitReq_27_11 = _GEN_386;
  wire          compressDataVec_hitReq_27_139;
  assign compressDataVec_hitReq_27_139 = _GEN_386;
  wire          _GEN_387 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'hB;
  wire          compressDataVec_hitReq_28_11;
  assign compressDataVec_hitReq_28_11 = _GEN_387;
  wire          compressDataVec_hitReq_28_139;
  assign compressDataVec_hitReq_28_139 = _GEN_387;
  wire          _GEN_388 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'hB;
  wire          compressDataVec_hitReq_29_11;
  assign compressDataVec_hitReq_29_11 = _GEN_388;
  wire          compressDataVec_hitReq_29_139;
  assign compressDataVec_hitReq_29_139 = _GEN_388;
  wire          _GEN_389 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'hB;
  wire          compressDataVec_hitReq_30_11;
  assign compressDataVec_hitReq_30_11 = _GEN_389;
  wire          compressDataVec_hitReq_30_139;
  assign compressDataVec_hitReq_30_139 = _GEN_389;
  wire          _GEN_390 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'hB;
  wire          compressDataVec_hitReq_31_11;
  assign compressDataVec_hitReq_31_11 = _GEN_390;
  wire          compressDataVec_hitReq_31_139;
  assign compressDataVec_hitReq_31_139 = _GEN_390;
  wire          compressDataVec_hitReq_32_11 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'hB;
  wire          compressDataVec_hitReq_33_11 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'hB;
  wire          compressDataVec_hitReq_34_11 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'hB;
  wire          compressDataVec_hitReq_35_11 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'hB;
  wire          compressDataVec_hitReq_36_11 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'hB;
  wire          compressDataVec_hitReq_37_11 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'hB;
  wire          compressDataVec_hitReq_38_11 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'hB;
  wire          compressDataVec_hitReq_39_11 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'hB;
  wire          compressDataVec_hitReq_40_11 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'hB;
  wire          compressDataVec_hitReq_41_11 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'hB;
  wire          compressDataVec_hitReq_42_11 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'hB;
  wire          compressDataVec_hitReq_43_11 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'hB;
  wire          compressDataVec_hitReq_44_11 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'hB;
  wire          compressDataVec_hitReq_45_11 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'hB;
  wire          compressDataVec_hitReq_46_11 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'hB;
  wire          compressDataVec_hitReq_47_11 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'hB;
  wire          compressDataVec_hitReq_48_11 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'hB;
  wire          compressDataVec_hitReq_49_11 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'hB;
  wire          compressDataVec_hitReq_50_11 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'hB;
  wire          compressDataVec_hitReq_51_11 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'hB;
  wire          compressDataVec_hitReq_52_11 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'hB;
  wire          compressDataVec_hitReq_53_11 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'hB;
  wire          compressDataVec_hitReq_54_11 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'hB;
  wire          compressDataVec_hitReq_55_11 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'hB;
  wire          compressDataVec_hitReq_56_11 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'hB;
  wire          compressDataVec_hitReq_57_11 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'hB;
  wire          compressDataVec_hitReq_58_11 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'hB;
  wire          compressDataVec_hitReq_59_11 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'hB;
  wire          compressDataVec_hitReq_60_11 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'hB;
  wire          compressDataVec_hitReq_61_11 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'hB;
  wire          compressDataVec_hitReq_62_11 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'hB;
  wire          compressDataVec_hitReq_63_11 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'hB;
  wire [7:0]    compressDataVec_selectReqData_11 =
    (compressDataVec_hitReq_0_11 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_11 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_11 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_11 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_11 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_11 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_11 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_11 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_11 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_11 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_11 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_11 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_11 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_11 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_11 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_11 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_11 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_11 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_11 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_11 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_11 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_11 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_11 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_11 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_11 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_11 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_11 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_11 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_11 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_11 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_11 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_11 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_11 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_11 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_11 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_11 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_11 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_11 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_11 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_11 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_11 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_11 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_11 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_11 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_11 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_11 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_11 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_11 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_11 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_11 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_11 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_11 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_11 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_11 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_11 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_11 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_11 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_11 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_11 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_11 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_11 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_11 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_11 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_11 ? source2Pipe[511:504] : 8'h0);
  wire          _GEN_391 = tailCount > 6'hB;
  wire          compressDataVec_useTail_11;
  assign compressDataVec_useTail_11 = _GEN_391;
  wire          compressDataVec_useTail_75;
  assign compressDataVec_useTail_75 = _GEN_391;
  wire          compressDataVec_useTail_107;
  assign compressDataVec_useTail_107 = _GEN_391;
  wire          _GEN_392 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'hC;
  wire          compressDataVec_hitReq_0_12;
  assign compressDataVec_hitReq_0_12 = _GEN_392;
  wire          compressDataVec_hitReq_0_140;
  assign compressDataVec_hitReq_0_140 = _GEN_392;
  wire          compressDataVec_hitReq_0_204;
  assign compressDataVec_hitReq_0_204 = _GEN_392;
  wire          _GEN_393 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'hC;
  wire          compressDataVec_hitReq_1_12;
  assign compressDataVec_hitReq_1_12 = _GEN_393;
  wire          compressDataVec_hitReq_1_140;
  assign compressDataVec_hitReq_1_140 = _GEN_393;
  wire          compressDataVec_hitReq_1_204;
  assign compressDataVec_hitReq_1_204 = _GEN_393;
  wire          _GEN_394 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'hC;
  wire          compressDataVec_hitReq_2_12;
  assign compressDataVec_hitReq_2_12 = _GEN_394;
  wire          compressDataVec_hitReq_2_140;
  assign compressDataVec_hitReq_2_140 = _GEN_394;
  wire          compressDataVec_hitReq_2_204;
  assign compressDataVec_hitReq_2_204 = _GEN_394;
  wire          _GEN_395 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'hC;
  wire          compressDataVec_hitReq_3_12;
  assign compressDataVec_hitReq_3_12 = _GEN_395;
  wire          compressDataVec_hitReq_3_140;
  assign compressDataVec_hitReq_3_140 = _GEN_395;
  wire          compressDataVec_hitReq_3_204;
  assign compressDataVec_hitReq_3_204 = _GEN_395;
  wire          _GEN_396 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'hC;
  wire          compressDataVec_hitReq_4_12;
  assign compressDataVec_hitReq_4_12 = _GEN_396;
  wire          compressDataVec_hitReq_4_140;
  assign compressDataVec_hitReq_4_140 = _GEN_396;
  wire          compressDataVec_hitReq_4_204;
  assign compressDataVec_hitReq_4_204 = _GEN_396;
  wire          _GEN_397 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'hC;
  wire          compressDataVec_hitReq_5_12;
  assign compressDataVec_hitReq_5_12 = _GEN_397;
  wire          compressDataVec_hitReq_5_140;
  assign compressDataVec_hitReq_5_140 = _GEN_397;
  wire          compressDataVec_hitReq_5_204;
  assign compressDataVec_hitReq_5_204 = _GEN_397;
  wire          _GEN_398 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'hC;
  wire          compressDataVec_hitReq_6_12;
  assign compressDataVec_hitReq_6_12 = _GEN_398;
  wire          compressDataVec_hitReq_6_140;
  assign compressDataVec_hitReq_6_140 = _GEN_398;
  wire          compressDataVec_hitReq_6_204;
  assign compressDataVec_hitReq_6_204 = _GEN_398;
  wire          _GEN_399 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'hC;
  wire          compressDataVec_hitReq_7_12;
  assign compressDataVec_hitReq_7_12 = _GEN_399;
  wire          compressDataVec_hitReq_7_140;
  assign compressDataVec_hitReq_7_140 = _GEN_399;
  wire          compressDataVec_hitReq_7_204;
  assign compressDataVec_hitReq_7_204 = _GEN_399;
  wire          _GEN_400 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'hC;
  wire          compressDataVec_hitReq_8_12;
  assign compressDataVec_hitReq_8_12 = _GEN_400;
  wire          compressDataVec_hitReq_8_140;
  assign compressDataVec_hitReq_8_140 = _GEN_400;
  wire          compressDataVec_hitReq_8_204;
  assign compressDataVec_hitReq_8_204 = _GEN_400;
  wire          _GEN_401 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'hC;
  wire          compressDataVec_hitReq_9_12;
  assign compressDataVec_hitReq_9_12 = _GEN_401;
  wire          compressDataVec_hitReq_9_140;
  assign compressDataVec_hitReq_9_140 = _GEN_401;
  wire          compressDataVec_hitReq_9_204;
  assign compressDataVec_hitReq_9_204 = _GEN_401;
  wire          _GEN_402 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'hC;
  wire          compressDataVec_hitReq_10_12;
  assign compressDataVec_hitReq_10_12 = _GEN_402;
  wire          compressDataVec_hitReq_10_140;
  assign compressDataVec_hitReq_10_140 = _GEN_402;
  wire          compressDataVec_hitReq_10_204;
  assign compressDataVec_hitReq_10_204 = _GEN_402;
  wire          _GEN_403 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'hC;
  wire          compressDataVec_hitReq_11_12;
  assign compressDataVec_hitReq_11_12 = _GEN_403;
  wire          compressDataVec_hitReq_11_140;
  assign compressDataVec_hitReq_11_140 = _GEN_403;
  wire          compressDataVec_hitReq_11_204;
  assign compressDataVec_hitReq_11_204 = _GEN_403;
  wire          _GEN_404 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'hC;
  wire          compressDataVec_hitReq_12_12;
  assign compressDataVec_hitReq_12_12 = _GEN_404;
  wire          compressDataVec_hitReq_12_140;
  assign compressDataVec_hitReq_12_140 = _GEN_404;
  wire          compressDataVec_hitReq_12_204;
  assign compressDataVec_hitReq_12_204 = _GEN_404;
  wire          _GEN_405 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'hC;
  wire          compressDataVec_hitReq_13_12;
  assign compressDataVec_hitReq_13_12 = _GEN_405;
  wire          compressDataVec_hitReq_13_140;
  assign compressDataVec_hitReq_13_140 = _GEN_405;
  wire          compressDataVec_hitReq_13_204;
  assign compressDataVec_hitReq_13_204 = _GEN_405;
  wire          _GEN_406 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'hC;
  wire          compressDataVec_hitReq_14_12;
  assign compressDataVec_hitReq_14_12 = _GEN_406;
  wire          compressDataVec_hitReq_14_140;
  assign compressDataVec_hitReq_14_140 = _GEN_406;
  wire          compressDataVec_hitReq_14_204;
  assign compressDataVec_hitReq_14_204 = _GEN_406;
  wire          _GEN_407 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'hC;
  wire          compressDataVec_hitReq_15_12;
  assign compressDataVec_hitReq_15_12 = _GEN_407;
  wire          compressDataVec_hitReq_15_140;
  assign compressDataVec_hitReq_15_140 = _GEN_407;
  wire          compressDataVec_hitReq_15_204;
  assign compressDataVec_hitReq_15_204 = _GEN_407;
  wire          _GEN_408 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'hC;
  wire          compressDataVec_hitReq_16_12;
  assign compressDataVec_hitReq_16_12 = _GEN_408;
  wire          compressDataVec_hitReq_16_140;
  assign compressDataVec_hitReq_16_140 = _GEN_408;
  wire          _GEN_409 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'hC;
  wire          compressDataVec_hitReq_17_12;
  assign compressDataVec_hitReq_17_12 = _GEN_409;
  wire          compressDataVec_hitReq_17_140;
  assign compressDataVec_hitReq_17_140 = _GEN_409;
  wire          _GEN_410 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'hC;
  wire          compressDataVec_hitReq_18_12;
  assign compressDataVec_hitReq_18_12 = _GEN_410;
  wire          compressDataVec_hitReq_18_140;
  assign compressDataVec_hitReq_18_140 = _GEN_410;
  wire          _GEN_411 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'hC;
  wire          compressDataVec_hitReq_19_12;
  assign compressDataVec_hitReq_19_12 = _GEN_411;
  wire          compressDataVec_hitReq_19_140;
  assign compressDataVec_hitReq_19_140 = _GEN_411;
  wire          _GEN_412 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'hC;
  wire          compressDataVec_hitReq_20_12;
  assign compressDataVec_hitReq_20_12 = _GEN_412;
  wire          compressDataVec_hitReq_20_140;
  assign compressDataVec_hitReq_20_140 = _GEN_412;
  wire          _GEN_413 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'hC;
  wire          compressDataVec_hitReq_21_12;
  assign compressDataVec_hitReq_21_12 = _GEN_413;
  wire          compressDataVec_hitReq_21_140;
  assign compressDataVec_hitReq_21_140 = _GEN_413;
  wire          _GEN_414 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'hC;
  wire          compressDataVec_hitReq_22_12;
  assign compressDataVec_hitReq_22_12 = _GEN_414;
  wire          compressDataVec_hitReq_22_140;
  assign compressDataVec_hitReq_22_140 = _GEN_414;
  wire          _GEN_415 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'hC;
  wire          compressDataVec_hitReq_23_12;
  assign compressDataVec_hitReq_23_12 = _GEN_415;
  wire          compressDataVec_hitReq_23_140;
  assign compressDataVec_hitReq_23_140 = _GEN_415;
  wire          _GEN_416 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'hC;
  wire          compressDataVec_hitReq_24_12;
  assign compressDataVec_hitReq_24_12 = _GEN_416;
  wire          compressDataVec_hitReq_24_140;
  assign compressDataVec_hitReq_24_140 = _GEN_416;
  wire          _GEN_417 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'hC;
  wire          compressDataVec_hitReq_25_12;
  assign compressDataVec_hitReq_25_12 = _GEN_417;
  wire          compressDataVec_hitReq_25_140;
  assign compressDataVec_hitReq_25_140 = _GEN_417;
  wire          _GEN_418 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'hC;
  wire          compressDataVec_hitReq_26_12;
  assign compressDataVec_hitReq_26_12 = _GEN_418;
  wire          compressDataVec_hitReq_26_140;
  assign compressDataVec_hitReq_26_140 = _GEN_418;
  wire          _GEN_419 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'hC;
  wire          compressDataVec_hitReq_27_12;
  assign compressDataVec_hitReq_27_12 = _GEN_419;
  wire          compressDataVec_hitReq_27_140;
  assign compressDataVec_hitReq_27_140 = _GEN_419;
  wire          _GEN_420 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'hC;
  wire          compressDataVec_hitReq_28_12;
  assign compressDataVec_hitReq_28_12 = _GEN_420;
  wire          compressDataVec_hitReq_28_140;
  assign compressDataVec_hitReq_28_140 = _GEN_420;
  wire          _GEN_421 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'hC;
  wire          compressDataVec_hitReq_29_12;
  assign compressDataVec_hitReq_29_12 = _GEN_421;
  wire          compressDataVec_hitReq_29_140;
  assign compressDataVec_hitReq_29_140 = _GEN_421;
  wire          _GEN_422 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'hC;
  wire          compressDataVec_hitReq_30_12;
  assign compressDataVec_hitReq_30_12 = _GEN_422;
  wire          compressDataVec_hitReq_30_140;
  assign compressDataVec_hitReq_30_140 = _GEN_422;
  wire          _GEN_423 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'hC;
  wire          compressDataVec_hitReq_31_12;
  assign compressDataVec_hitReq_31_12 = _GEN_423;
  wire          compressDataVec_hitReq_31_140;
  assign compressDataVec_hitReq_31_140 = _GEN_423;
  wire          compressDataVec_hitReq_32_12 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'hC;
  wire          compressDataVec_hitReq_33_12 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'hC;
  wire          compressDataVec_hitReq_34_12 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'hC;
  wire          compressDataVec_hitReq_35_12 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'hC;
  wire          compressDataVec_hitReq_36_12 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'hC;
  wire          compressDataVec_hitReq_37_12 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'hC;
  wire          compressDataVec_hitReq_38_12 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'hC;
  wire          compressDataVec_hitReq_39_12 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'hC;
  wire          compressDataVec_hitReq_40_12 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'hC;
  wire          compressDataVec_hitReq_41_12 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'hC;
  wire          compressDataVec_hitReq_42_12 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'hC;
  wire          compressDataVec_hitReq_43_12 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'hC;
  wire          compressDataVec_hitReq_44_12 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'hC;
  wire          compressDataVec_hitReq_45_12 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'hC;
  wire          compressDataVec_hitReq_46_12 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'hC;
  wire          compressDataVec_hitReq_47_12 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'hC;
  wire          compressDataVec_hitReq_48_12 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'hC;
  wire          compressDataVec_hitReq_49_12 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'hC;
  wire          compressDataVec_hitReq_50_12 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'hC;
  wire          compressDataVec_hitReq_51_12 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'hC;
  wire          compressDataVec_hitReq_52_12 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'hC;
  wire          compressDataVec_hitReq_53_12 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'hC;
  wire          compressDataVec_hitReq_54_12 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'hC;
  wire          compressDataVec_hitReq_55_12 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'hC;
  wire          compressDataVec_hitReq_56_12 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'hC;
  wire          compressDataVec_hitReq_57_12 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'hC;
  wire          compressDataVec_hitReq_58_12 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'hC;
  wire          compressDataVec_hitReq_59_12 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'hC;
  wire          compressDataVec_hitReq_60_12 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'hC;
  wire          compressDataVec_hitReq_61_12 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'hC;
  wire          compressDataVec_hitReq_62_12 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'hC;
  wire          compressDataVec_hitReq_63_12 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'hC;
  wire [7:0]    compressDataVec_selectReqData_12 =
    (compressDataVec_hitReq_0_12 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_12 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_12 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_12 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_12 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_12 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_12 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_12 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_12 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_12 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_12 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_12 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_12 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_12 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_12 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_12 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_12 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_12 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_12 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_12 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_12 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_12 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_12 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_12 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_12 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_12 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_12 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_12 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_12 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_12 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_12 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_12 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_12 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_12 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_12 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_12 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_12 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_12 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_12 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_12 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_12 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_12 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_12 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_12 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_12 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_12 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_12 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_12 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_12 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_12 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_12 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_12 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_12 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_12 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_12 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_12 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_12 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_12 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_12 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_12 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_12 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_12 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_12 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_12 ? source2Pipe[511:504] : 8'h0);
  wire          _GEN_424 = tailCount > 6'hC;
  wire          compressDataVec_useTail_12;
  assign compressDataVec_useTail_12 = _GEN_424;
  wire          compressDataVec_useTail_76;
  assign compressDataVec_useTail_76 = _GEN_424;
  wire          compressDataVec_useTail_108;
  assign compressDataVec_useTail_108 = _GEN_424;
  wire          _GEN_425 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'hD;
  wire          compressDataVec_hitReq_0_13;
  assign compressDataVec_hitReq_0_13 = _GEN_425;
  wire          compressDataVec_hitReq_0_141;
  assign compressDataVec_hitReq_0_141 = _GEN_425;
  wire          compressDataVec_hitReq_0_205;
  assign compressDataVec_hitReq_0_205 = _GEN_425;
  wire          _GEN_426 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'hD;
  wire          compressDataVec_hitReq_1_13;
  assign compressDataVec_hitReq_1_13 = _GEN_426;
  wire          compressDataVec_hitReq_1_141;
  assign compressDataVec_hitReq_1_141 = _GEN_426;
  wire          compressDataVec_hitReq_1_205;
  assign compressDataVec_hitReq_1_205 = _GEN_426;
  wire          _GEN_427 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'hD;
  wire          compressDataVec_hitReq_2_13;
  assign compressDataVec_hitReq_2_13 = _GEN_427;
  wire          compressDataVec_hitReq_2_141;
  assign compressDataVec_hitReq_2_141 = _GEN_427;
  wire          compressDataVec_hitReq_2_205;
  assign compressDataVec_hitReq_2_205 = _GEN_427;
  wire          _GEN_428 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'hD;
  wire          compressDataVec_hitReq_3_13;
  assign compressDataVec_hitReq_3_13 = _GEN_428;
  wire          compressDataVec_hitReq_3_141;
  assign compressDataVec_hitReq_3_141 = _GEN_428;
  wire          compressDataVec_hitReq_3_205;
  assign compressDataVec_hitReq_3_205 = _GEN_428;
  wire          _GEN_429 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'hD;
  wire          compressDataVec_hitReq_4_13;
  assign compressDataVec_hitReq_4_13 = _GEN_429;
  wire          compressDataVec_hitReq_4_141;
  assign compressDataVec_hitReq_4_141 = _GEN_429;
  wire          compressDataVec_hitReq_4_205;
  assign compressDataVec_hitReq_4_205 = _GEN_429;
  wire          _GEN_430 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'hD;
  wire          compressDataVec_hitReq_5_13;
  assign compressDataVec_hitReq_5_13 = _GEN_430;
  wire          compressDataVec_hitReq_5_141;
  assign compressDataVec_hitReq_5_141 = _GEN_430;
  wire          compressDataVec_hitReq_5_205;
  assign compressDataVec_hitReq_5_205 = _GEN_430;
  wire          _GEN_431 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'hD;
  wire          compressDataVec_hitReq_6_13;
  assign compressDataVec_hitReq_6_13 = _GEN_431;
  wire          compressDataVec_hitReq_6_141;
  assign compressDataVec_hitReq_6_141 = _GEN_431;
  wire          compressDataVec_hitReq_6_205;
  assign compressDataVec_hitReq_6_205 = _GEN_431;
  wire          _GEN_432 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'hD;
  wire          compressDataVec_hitReq_7_13;
  assign compressDataVec_hitReq_7_13 = _GEN_432;
  wire          compressDataVec_hitReq_7_141;
  assign compressDataVec_hitReq_7_141 = _GEN_432;
  wire          compressDataVec_hitReq_7_205;
  assign compressDataVec_hitReq_7_205 = _GEN_432;
  wire          _GEN_433 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'hD;
  wire          compressDataVec_hitReq_8_13;
  assign compressDataVec_hitReq_8_13 = _GEN_433;
  wire          compressDataVec_hitReq_8_141;
  assign compressDataVec_hitReq_8_141 = _GEN_433;
  wire          compressDataVec_hitReq_8_205;
  assign compressDataVec_hitReq_8_205 = _GEN_433;
  wire          _GEN_434 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'hD;
  wire          compressDataVec_hitReq_9_13;
  assign compressDataVec_hitReq_9_13 = _GEN_434;
  wire          compressDataVec_hitReq_9_141;
  assign compressDataVec_hitReq_9_141 = _GEN_434;
  wire          compressDataVec_hitReq_9_205;
  assign compressDataVec_hitReq_9_205 = _GEN_434;
  wire          _GEN_435 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'hD;
  wire          compressDataVec_hitReq_10_13;
  assign compressDataVec_hitReq_10_13 = _GEN_435;
  wire          compressDataVec_hitReq_10_141;
  assign compressDataVec_hitReq_10_141 = _GEN_435;
  wire          compressDataVec_hitReq_10_205;
  assign compressDataVec_hitReq_10_205 = _GEN_435;
  wire          _GEN_436 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'hD;
  wire          compressDataVec_hitReq_11_13;
  assign compressDataVec_hitReq_11_13 = _GEN_436;
  wire          compressDataVec_hitReq_11_141;
  assign compressDataVec_hitReq_11_141 = _GEN_436;
  wire          compressDataVec_hitReq_11_205;
  assign compressDataVec_hitReq_11_205 = _GEN_436;
  wire          _GEN_437 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'hD;
  wire          compressDataVec_hitReq_12_13;
  assign compressDataVec_hitReq_12_13 = _GEN_437;
  wire          compressDataVec_hitReq_12_141;
  assign compressDataVec_hitReq_12_141 = _GEN_437;
  wire          compressDataVec_hitReq_12_205;
  assign compressDataVec_hitReq_12_205 = _GEN_437;
  wire          _GEN_438 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'hD;
  wire          compressDataVec_hitReq_13_13;
  assign compressDataVec_hitReq_13_13 = _GEN_438;
  wire          compressDataVec_hitReq_13_141;
  assign compressDataVec_hitReq_13_141 = _GEN_438;
  wire          compressDataVec_hitReq_13_205;
  assign compressDataVec_hitReq_13_205 = _GEN_438;
  wire          _GEN_439 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'hD;
  wire          compressDataVec_hitReq_14_13;
  assign compressDataVec_hitReq_14_13 = _GEN_439;
  wire          compressDataVec_hitReq_14_141;
  assign compressDataVec_hitReq_14_141 = _GEN_439;
  wire          compressDataVec_hitReq_14_205;
  assign compressDataVec_hitReq_14_205 = _GEN_439;
  wire          _GEN_440 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'hD;
  wire          compressDataVec_hitReq_15_13;
  assign compressDataVec_hitReq_15_13 = _GEN_440;
  wire          compressDataVec_hitReq_15_141;
  assign compressDataVec_hitReq_15_141 = _GEN_440;
  wire          compressDataVec_hitReq_15_205;
  assign compressDataVec_hitReq_15_205 = _GEN_440;
  wire          _GEN_441 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'hD;
  wire          compressDataVec_hitReq_16_13;
  assign compressDataVec_hitReq_16_13 = _GEN_441;
  wire          compressDataVec_hitReq_16_141;
  assign compressDataVec_hitReq_16_141 = _GEN_441;
  wire          _GEN_442 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'hD;
  wire          compressDataVec_hitReq_17_13;
  assign compressDataVec_hitReq_17_13 = _GEN_442;
  wire          compressDataVec_hitReq_17_141;
  assign compressDataVec_hitReq_17_141 = _GEN_442;
  wire          _GEN_443 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'hD;
  wire          compressDataVec_hitReq_18_13;
  assign compressDataVec_hitReq_18_13 = _GEN_443;
  wire          compressDataVec_hitReq_18_141;
  assign compressDataVec_hitReq_18_141 = _GEN_443;
  wire          _GEN_444 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'hD;
  wire          compressDataVec_hitReq_19_13;
  assign compressDataVec_hitReq_19_13 = _GEN_444;
  wire          compressDataVec_hitReq_19_141;
  assign compressDataVec_hitReq_19_141 = _GEN_444;
  wire          _GEN_445 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'hD;
  wire          compressDataVec_hitReq_20_13;
  assign compressDataVec_hitReq_20_13 = _GEN_445;
  wire          compressDataVec_hitReq_20_141;
  assign compressDataVec_hitReq_20_141 = _GEN_445;
  wire          _GEN_446 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'hD;
  wire          compressDataVec_hitReq_21_13;
  assign compressDataVec_hitReq_21_13 = _GEN_446;
  wire          compressDataVec_hitReq_21_141;
  assign compressDataVec_hitReq_21_141 = _GEN_446;
  wire          _GEN_447 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'hD;
  wire          compressDataVec_hitReq_22_13;
  assign compressDataVec_hitReq_22_13 = _GEN_447;
  wire          compressDataVec_hitReq_22_141;
  assign compressDataVec_hitReq_22_141 = _GEN_447;
  wire          _GEN_448 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'hD;
  wire          compressDataVec_hitReq_23_13;
  assign compressDataVec_hitReq_23_13 = _GEN_448;
  wire          compressDataVec_hitReq_23_141;
  assign compressDataVec_hitReq_23_141 = _GEN_448;
  wire          _GEN_449 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'hD;
  wire          compressDataVec_hitReq_24_13;
  assign compressDataVec_hitReq_24_13 = _GEN_449;
  wire          compressDataVec_hitReq_24_141;
  assign compressDataVec_hitReq_24_141 = _GEN_449;
  wire          _GEN_450 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'hD;
  wire          compressDataVec_hitReq_25_13;
  assign compressDataVec_hitReq_25_13 = _GEN_450;
  wire          compressDataVec_hitReq_25_141;
  assign compressDataVec_hitReq_25_141 = _GEN_450;
  wire          _GEN_451 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'hD;
  wire          compressDataVec_hitReq_26_13;
  assign compressDataVec_hitReq_26_13 = _GEN_451;
  wire          compressDataVec_hitReq_26_141;
  assign compressDataVec_hitReq_26_141 = _GEN_451;
  wire          _GEN_452 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'hD;
  wire          compressDataVec_hitReq_27_13;
  assign compressDataVec_hitReq_27_13 = _GEN_452;
  wire          compressDataVec_hitReq_27_141;
  assign compressDataVec_hitReq_27_141 = _GEN_452;
  wire          _GEN_453 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'hD;
  wire          compressDataVec_hitReq_28_13;
  assign compressDataVec_hitReq_28_13 = _GEN_453;
  wire          compressDataVec_hitReq_28_141;
  assign compressDataVec_hitReq_28_141 = _GEN_453;
  wire          _GEN_454 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'hD;
  wire          compressDataVec_hitReq_29_13;
  assign compressDataVec_hitReq_29_13 = _GEN_454;
  wire          compressDataVec_hitReq_29_141;
  assign compressDataVec_hitReq_29_141 = _GEN_454;
  wire          _GEN_455 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'hD;
  wire          compressDataVec_hitReq_30_13;
  assign compressDataVec_hitReq_30_13 = _GEN_455;
  wire          compressDataVec_hitReq_30_141;
  assign compressDataVec_hitReq_30_141 = _GEN_455;
  wire          _GEN_456 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'hD;
  wire          compressDataVec_hitReq_31_13;
  assign compressDataVec_hitReq_31_13 = _GEN_456;
  wire          compressDataVec_hitReq_31_141;
  assign compressDataVec_hitReq_31_141 = _GEN_456;
  wire          compressDataVec_hitReq_32_13 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'hD;
  wire          compressDataVec_hitReq_33_13 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'hD;
  wire          compressDataVec_hitReq_34_13 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'hD;
  wire          compressDataVec_hitReq_35_13 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'hD;
  wire          compressDataVec_hitReq_36_13 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'hD;
  wire          compressDataVec_hitReq_37_13 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'hD;
  wire          compressDataVec_hitReq_38_13 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'hD;
  wire          compressDataVec_hitReq_39_13 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'hD;
  wire          compressDataVec_hitReq_40_13 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'hD;
  wire          compressDataVec_hitReq_41_13 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'hD;
  wire          compressDataVec_hitReq_42_13 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'hD;
  wire          compressDataVec_hitReq_43_13 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'hD;
  wire          compressDataVec_hitReq_44_13 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'hD;
  wire          compressDataVec_hitReq_45_13 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'hD;
  wire          compressDataVec_hitReq_46_13 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'hD;
  wire          compressDataVec_hitReq_47_13 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'hD;
  wire          compressDataVec_hitReq_48_13 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'hD;
  wire          compressDataVec_hitReq_49_13 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'hD;
  wire          compressDataVec_hitReq_50_13 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'hD;
  wire          compressDataVec_hitReq_51_13 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'hD;
  wire          compressDataVec_hitReq_52_13 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'hD;
  wire          compressDataVec_hitReq_53_13 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'hD;
  wire          compressDataVec_hitReq_54_13 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'hD;
  wire          compressDataVec_hitReq_55_13 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'hD;
  wire          compressDataVec_hitReq_56_13 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'hD;
  wire          compressDataVec_hitReq_57_13 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'hD;
  wire          compressDataVec_hitReq_58_13 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'hD;
  wire          compressDataVec_hitReq_59_13 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'hD;
  wire          compressDataVec_hitReq_60_13 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'hD;
  wire          compressDataVec_hitReq_61_13 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'hD;
  wire          compressDataVec_hitReq_62_13 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'hD;
  wire          compressDataVec_hitReq_63_13 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'hD;
  wire [7:0]    compressDataVec_selectReqData_13 =
    (compressDataVec_hitReq_0_13 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_13 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_13 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_13 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_13 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_13 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_13 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_13 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_13 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_13 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_13 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_13 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_13 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_13 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_13 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_13 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_13 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_13 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_13 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_13 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_13 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_13 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_13 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_13 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_13 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_13 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_13 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_13 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_13 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_13 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_13 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_13 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_13 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_13 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_13 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_13 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_13 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_13 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_13 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_13 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_13 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_13 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_13 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_13 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_13 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_13 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_13 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_13 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_13 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_13 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_13 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_13 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_13 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_13 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_13 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_13 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_13 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_13 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_13 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_13 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_13 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_13 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_13 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_13 ? source2Pipe[511:504] : 8'h0);
  wire          _GEN_457 = tailCount > 6'hD;
  wire          compressDataVec_useTail_13;
  assign compressDataVec_useTail_13 = _GEN_457;
  wire          compressDataVec_useTail_77;
  assign compressDataVec_useTail_77 = _GEN_457;
  wire          compressDataVec_useTail_109;
  assign compressDataVec_useTail_109 = _GEN_457;
  wire          _GEN_458 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'hE;
  wire          compressDataVec_hitReq_0_14;
  assign compressDataVec_hitReq_0_14 = _GEN_458;
  wire          compressDataVec_hitReq_0_142;
  assign compressDataVec_hitReq_0_142 = _GEN_458;
  wire          compressDataVec_hitReq_0_206;
  assign compressDataVec_hitReq_0_206 = _GEN_458;
  wire          _GEN_459 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'hE;
  wire          compressDataVec_hitReq_1_14;
  assign compressDataVec_hitReq_1_14 = _GEN_459;
  wire          compressDataVec_hitReq_1_142;
  assign compressDataVec_hitReq_1_142 = _GEN_459;
  wire          compressDataVec_hitReq_1_206;
  assign compressDataVec_hitReq_1_206 = _GEN_459;
  wire          _GEN_460 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'hE;
  wire          compressDataVec_hitReq_2_14;
  assign compressDataVec_hitReq_2_14 = _GEN_460;
  wire          compressDataVec_hitReq_2_142;
  assign compressDataVec_hitReq_2_142 = _GEN_460;
  wire          compressDataVec_hitReq_2_206;
  assign compressDataVec_hitReq_2_206 = _GEN_460;
  wire          _GEN_461 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'hE;
  wire          compressDataVec_hitReq_3_14;
  assign compressDataVec_hitReq_3_14 = _GEN_461;
  wire          compressDataVec_hitReq_3_142;
  assign compressDataVec_hitReq_3_142 = _GEN_461;
  wire          compressDataVec_hitReq_3_206;
  assign compressDataVec_hitReq_3_206 = _GEN_461;
  wire          _GEN_462 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'hE;
  wire          compressDataVec_hitReq_4_14;
  assign compressDataVec_hitReq_4_14 = _GEN_462;
  wire          compressDataVec_hitReq_4_142;
  assign compressDataVec_hitReq_4_142 = _GEN_462;
  wire          compressDataVec_hitReq_4_206;
  assign compressDataVec_hitReq_4_206 = _GEN_462;
  wire          _GEN_463 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'hE;
  wire          compressDataVec_hitReq_5_14;
  assign compressDataVec_hitReq_5_14 = _GEN_463;
  wire          compressDataVec_hitReq_5_142;
  assign compressDataVec_hitReq_5_142 = _GEN_463;
  wire          compressDataVec_hitReq_5_206;
  assign compressDataVec_hitReq_5_206 = _GEN_463;
  wire          _GEN_464 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'hE;
  wire          compressDataVec_hitReq_6_14;
  assign compressDataVec_hitReq_6_14 = _GEN_464;
  wire          compressDataVec_hitReq_6_142;
  assign compressDataVec_hitReq_6_142 = _GEN_464;
  wire          compressDataVec_hitReq_6_206;
  assign compressDataVec_hitReq_6_206 = _GEN_464;
  wire          _GEN_465 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'hE;
  wire          compressDataVec_hitReq_7_14;
  assign compressDataVec_hitReq_7_14 = _GEN_465;
  wire          compressDataVec_hitReq_7_142;
  assign compressDataVec_hitReq_7_142 = _GEN_465;
  wire          compressDataVec_hitReq_7_206;
  assign compressDataVec_hitReq_7_206 = _GEN_465;
  wire          _GEN_466 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'hE;
  wire          compressDataVec_hitReq_8_14;
  assign compressDataVec_hitReq_8_14 = _GEN_466;
  wire          compressDataVec_hitReq_8_142;
  assign compressDataVec_hitReq_8_142 = _GEN_466;
  wire          compressDataVec_hitReq_8_206;
  assign compressDataVec_hitReq_8_206 = _GEN_466;
  wire          _GEN_467 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'hE;
  wire          compressDataVec_hitReq_9_14;
  assign compressDataVec_hitReq_9_14 = _GEN_467;
  wire          compressDataVec_hitReq_9_142;
  assign compressDataVec_hitReq_9_142 = _GEN_467;
  wire          compressDataVec_hitReq_9_206;
  assign compressDataVec_hitReq_9_206 = _GEN_467;
  wire          _GEN_468 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'hE;
  wire          compressDataVec_hitReq_10_14;
  assign compressDataVec_hitReq_10_14 = _GEN_468;
  wire          compressDataVec_hitReq_10_142;
  assign compressDataVec_hitReq_10_142 = _GEN_468;
  wire          compressDataVec_hitReq_10_206;
  assign compressDataVec_hitReq_10_206 = _GEN_468;
  wire          _GEN_469 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'hE;
  wire          compressDataVec_hitReq_11_14;
  assign compressDataVec_hitReq_11_14 = _GEN_469;
  wire          compressDataVec_hitReq_11_142;
  assign compressDataVec_hitReq_11_142 = _GEN_469;
  wire          compressDataVec_hitReq_11_206;
  assign compressDataVec_hitReq_11_206 = _GEN_469;
  wire          _GEN_470 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'hE;
  wire          compressDataVec_hitReq_12_14;
  assign compressDataVec_hitReq_12_14 = _GEN_470;
  wire          compressDataVec_hitReq_12_142;
  assign compressDataVec_hitReq_12_142 = _GEN_470;
  wire          compressDataVec_hitReq_12_206;
  assign compressDataVec_hitReq_12_206 = _GEN_470;
  wire          _GEN_471 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'hE;
  wire          compressDataVec_hitReq_13_14;
  assign compressDataVec_hitReq_13_14 = _GEN_471;
  wire          compressDataVec_hitReq_13_142;
  assign compressDataVec_hitReq_13_142 = _GEN_471;
  wire          compressDataVec_hitReq_13_206;
  assign compressDataVec_hitReq_13_206 = _GEN_471;
  wire          _GEN_472 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'hE;
  wire          compressDataVec_hitReq_14_14;
  assign compressDataVec_hitReq_14_14 = _GEN_472;
  wire          compressDataVec_hitReq_14_142;
  assign compressDataVec_hitReq_14_142 = _GEN_472;
  wire          compressDataVec_hitReq_14_206;
  assign compressDataVec_hitReq_14_206 = _GEN_472;
  wire          _GEN_473 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'hE;
  wire          compressDataVec_hitReq_15_14;
  assign compressDataVec_hitReq_15_14 = _GEN_473;
  wire          compressDataVec_hitReq_15_142;
  assign compressDataVec_hitReq_15_142 = _GEN_473;
  wire          compressDataVec_hitReq_15_206;
  assign compressDataVec_hitReq_15_206 = _GEN_473;
  wire          _GEN_474 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'hE;
  wire          compressDataVec_hitReq_16_14;
  assign compressDataVec_hitReq_16_14 = _GEN_474;
  wire          compressDataVec_hitReq_16_142;
  assign compressDataVec_hitReq_16_142 = _GEN_474;
  wire          _GEN_475 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'hE;
  wire          compressDataVec_hitReq_17_14;
  assign compressDataVec_hitReq_17_14 = _GEN_475;
  wire          compressDataVec_hitReq_17_142;
  assign compressDataVec_hitReq_17_142 = _GEN_475;
  wire          _GEN_476 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'hE;
  wire          compressDataVec_hitReq_18_14;
  assign compressDataVec_hitReq_18_14 = _GEN_476;
  wire          compressDataVec_hitReq_18_142;
  assign compressDataVec_hitReq_18_142 = _GEN_476;
  wire          _GEN_477 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'hE;
  wire          compressDataVec_hitReq_19_14;
  assign compressDataVec_hitReq_19_14 = _GEN_477;
  wire          compressDataVec_hitReq_19_142;
  assign compressDataVec_hitReq_19_142 = _GEN_477;
  wire          _GEN_478 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'hE;
  wire          compressDataVec_hitReq_20_14;
  assign compressDataVec_hitReq_20_14 = _GEN_478;
  wire          compressDataVec_hitReq_20_142;
  assign compressDataVec_hitReq_20_142 = _GEN_478;
  wire          _GEN_479 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'hE;
  wire          compressDataVec_hitReq_21_14;
  assign compressDataVec_hitReq_21_14 = _GEN_479;
  wire          compressDataVec_hitReq_21_142;
  assign compressDataVec_hitReq_21_142 = _GEN_479;
  wire          _GEN_480 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'hE;
  wire          compressDataVec_hitReq_22_14;
  assign compressDataVec_hitReq_22_14 = _GEN_480;
  wire          compressDataVec_hitReq_22_142;
  assign compressDataVec_hitReq_22_142 = _GEN_480;
  wire          _GEN_481 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'hE;
  wire          compressDataVec_hitReq_23_14;
  assign compressDataVec_hitReq_23_14 = _GEN_481;
  wire          compressDataVec_hitReq_23_142;
  assign compressDataVec_hitReq_23_142 = _GEN_481;
  wire          _GEN_482 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'hE;
  wire          compressDataVec_hitReq_24_14;
  assign compressDataVec_hitReq_24_14 = _GEN_482;
  wire          compressDataVec_hitReq_24_142;
  assign compressDataVec_hitReq_24_142 = _GEN_482;
  wire          _GEN_483 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'hE;
  wire          compressDataVec_hitReq_25_14;
  assign compressDataVec_hitReq_25_14 = _GEN_483;
  wire          compressDataVec_hitReq_25_142;
  assign compressDataVec_hitReq_25_142 = _GEN_483;
  wire          _GEN_484 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'hE;
  wire          compressDataVec_hitReq_26_14;
  assign compressDataVec_hitReq_26_14 = _GEN_484;
  wire          compressDataVec_hitReq_26_142;
  assign compressDataVec_hitReq_26_142 = _GEN_484;
  wire          _GEN_485 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'hE;
  wire          compressDataVec_hitReq_27_14;
  assign compressDataVec_hitReq_27_14 = _GEN_485;
  wire          compressDataVec_hitReq_27_142;
  assign compressDataVec_hitReq_27_142 = _GEN_485;
  wire          _GEN_486 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'hE;
  wire          compressDataVec_hitReq_28_14;
  assign compressDataVec_hitReq_28_14 = _GEN_486;
  wire          compressDataVec_hitReq_28_142;
  assign compressDataVec_hitReq_28_142 = _GEN_486;
  wire          _GEN_487 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'hE;
  wire          compressDataVec_hitReq_29_14;
  assign compressDataVec_hitReq_29_14 = _GEN_487;
  wire          compressDataVec_hitReq_29_142;
  assign compressDataVec_hitReq_29_142 = _GEN_487;
  wire          _GEN_488 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'hE;
  wire          compressDataVec_hitReq_30_14;
  assign compressDataVec_hitReq_30_14 = _GEN_488;
  wire          compressDataVec_hitReq_30_142;
  assign compressDataVec_hitReq_30_142 = _GEN_488;
  wire          _GEN_489 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'hE;
  wire          compressDataVec_hitReq_31_14;
  assign compressDataVec_hitReq_31_14 = _GEN_489;
  wire          compressDataVec_hitReq_31_142;
  assign compressDataVec_hitReq_31_142 = _GEN_489;
  wire          compressDataVec_hitReq_32_14 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'hE;
  wire          compressDataVec_hitReq_33_14 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'hE;
  wire          compressDataVec_hitReq_34_14 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'hE;
  wire          compressDataVec_hitReq_35_14 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'hE;
  wire          compressDataVec_hitReq_36_14 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'hE;
  wire          compressDataVec_hitReq_37_14 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'hE;
  wire          compressDataVec_hitReq_38_14 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'hE;
  wire          compressDataVec_hitReq_39_14 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'hE;
  wire          compressDataVec_hitReq_40_14 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'hE;
  wire          compressDataVec_hitReq_41_14 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'hE;
  wire          compressDataVec_hitReq_42_14 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'hE;
  wire          compressDataVec_hitReq_43_14 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'hE;
  wire          compressDataVec_hitReq_44_14 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'hE;
  wire          compressDataVec_hitReq_45_14 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'hE;
  wire          compressDataVec_hitReq_46_14 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'hE;
  wire          compressDataVec_hitReq_47_14 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'hE;
  wire          compressDataVec_hitReq_48_14 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'hE;
  wire          compressDataVec_hitReq_49_14 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'hE;
  wire          compressDataVec_hitReq_50_14 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'hE;
  wire          compressDataVec_hitReq_51_14 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'hE;
  wire          compressDataVec_hitReq_52_14 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'hE;
  wire          compressDataVec_hitReq_53_14 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'hE;
  wire          compressDataVec_hitReq_54_14 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'hE;
  wire          compressDataVec_hitReq_55_14 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'hE;
  wire          compressDataVec_hitReq_56_14 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'hE;
  wire          compressDataVec_hitReq_57_14 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'hE;
  wire          compressDataVec_hitReq_58_14 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'hE;
  wire          compressDataVec_hitReq_59_14 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'hE;
  wire          compressDataVec_hitReq_60_14 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'hE;
  wire          compressDataVec_hitReq_61_14 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'hE;
  wire          compressDataVec_hitReq_62_14 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'hE;
  wire          compressDataVec_hitReq_63_14 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'hE;
  wire [7:0]    compressDataVec_selectReqData_14 =
    (compressDataVec_hitReq_0_14 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_14 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_14 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_14 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_14 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_14 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_14 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_14 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_14 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_14 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_14 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_14 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_14 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_14 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_14 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_14 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_14 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_14 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_14 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_14 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_14 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_14 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_14 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_14 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_14 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_14 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_14 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_14 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_14 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_14 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_14 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_14 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_14 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_14 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_14 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_14 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_14 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_14 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_14 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_14 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_14 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_14 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_14 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_14 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_14 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_14 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_14 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_14 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_14 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_14 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_14 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_14 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_14 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_14 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_14 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_14 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_14 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_14 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_14 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_14 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_14 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_14 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_14 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_14 ? source2Pipe[511:504] : 8'h0);
  wire          _GEN_490 = tailCount > 6'hE;
  wire          compressDataVec_useTail_14;
  assign compressDataVec_useTail_14 = _GEN_490;
  wire          compressDataVec_useTail_78;
  assign compressDataVec_useTail_78 = _GEN_490;
  wire          compressDataVec_useTail_110;
  assign compressDataVec_useTail_110 = _GEN_490;
  wire          _GEN_491 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'hF;
  wire          compressDataVec_hitReq_0_15;
  assign compressDataVec_hitReq_0_15 = _GEN_491;
  wire          compressDataVec_hitReq_0_143;
  assign compressDataVec_hitReq_0_143 = _GEN_491;
  wire          compressDataVec_hitReq_0_207;
  assign compressDataVec_hitReq_0_207 = _GEN_491;
  wire          _GEN_492 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'hF;
  wire          compressDataVec_hitReq_1_15;
  assign compressDataVec_hitReq_1_15 = _GEN_492;
  wire          compressDataVec_hitReq_1_143;
  assign compressDataVec_hitReq_1_143 = _GEN_492;
  wire          compressDataVec_hitReq_1_207;
  assign compressDataVec_hitReq_1_207 = _GEN_492;
  wire          _GEN_493 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'hF;
  wire          compressDataVec_hitReq_2_15;
  assign compressDataVec_hitReq_2_15 = _GEN_493;
  wire          compressDataVec_hitReq_2_143;
  assign compressDataVec_hitReq_2_143 = _GEN_493;
  wire          compressDataVec_hitReq_2_207;
  assign compressDataVec_hitReq_2_207 = _GEN_493;
  wire          _GEN_494 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'hF;
  wire          compressDataVec_hitReq_3_15;
  assign compressDataVec_hitReq_3_15 = _GEN_494;
  wire          compressDataVec_hitReq_3_143;
  assign compressDataVec_hitReq_3_143 = _GEN_494;
  wire          compressDataVec_hitReq_3_207;
  assign compressDataVec_hitReq_3_207 = _GEN_494;
  wire          _GEN_495 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'hF;
  wire          compressDataVec_hitReq_4_15;
  assign compressDataVec_hitReq_4_15 = _GEN_495;
  wire          compressDataVec_hitReq_4_143;
  assign compressDataVec_hitReq_4_143 = _GEN_495;
  wire          compressDataVec_hitReq_4_207;
  assign compressDataVec_hitReq_4_207 = _GEN_495;
  wire          _GEN_496 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'hF;
  wire          compressDataVec_hitReq_5_15;
  assign compressDataVec_hitReq_5_15 = _GEN_496;
  wire          compressDataVec_hitReq_5_143;
  assign compressDataVec_hitReq_5_143 = _GEN_496;
  wire          compressDataVec_hitReq_5_207;
  assign compressDataVec_hitReq_5_207 = _GEN_496;
  wire          _GEN_497 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'hF;
  wire          compressDataVec_hitReq_6_15;
  assign compressDataVec_hitReq_6_15 = _GEN_497;
  wire          compressDataVec_hitReq_6_143;
  assign compressDataVec_hitReq_6_143 = _GEN_497;
  wire          compressDataVec_hitReq_6_207;
  assign compressDataVec_hitReq_6_207 = _GEN_497;
  wire          _GEN_498 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'hF;
  wire          compressDataVec_hitReq_7_15;
  assign compressDataVec_hitReq_7_15 = _GEN_498;
  wire          compressDataVec_hitReq_7_143;
  assign compressDataVec_hitReq_7_143 = _GEN_498;
  wire          compressDataVec_hitReq_7_207;
  assign compressDataVec_hitReq_7_207 = _GEN_498;
  wire          _GEN_499 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'hF;
  wire          compressDataVec_hitReq_8_15;
  assign compressDataVec_hitReq_8_15 = _GEN_499;
  wire          compressDataVec_hitReq_8_143;
  assign compressDataVec_hitReq_8_143 = _GEN_499;
  wire          compressDataVec_hitReq_8_207;
  assign compressDataVec_hitReq_8_207 = _GEN_499;
  wire          _GEN_500 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'hF;
  wire          compressDataVec_hitReq_9_15;
  assign compressDataVec_hitReq_9_15 = _GEN_500;
  wire          compressDataVec_hitReq_9_143;
  assign compressDataVec_hitReq_9_143 = _GEN_500;
  wire          compressDataVec_hitReq_9_207;
  assign compressDataVec_hitReq_9_207 = _GEN_500;
  wire          _GEN_501 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'hF;
  wire          compressDataVec_hitReq_10_15;
  assign compressDataVec_hitReq_10_15 = _GEN_501;
  wire          compressDataVec_hitReq_10_143;
  assign compressDataVec_hitReq_10_143 = _GEN_501;
  wire          compressDataVec_hitReq_10_207;
  assign compressDataVec_hitReq_10_207 = _GEN_501;
  wire          _GEN_502 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'hF;
  wire          compressDataVec_hitReq_11_15;
  assign compressDataVec_hitReq_11_15 = _GEN_502;
  wire          compressDataVec_hitReq_11_143;
  assign compressDataVec_hitReq_11_143 = _GEN_502;
  wire          compressDataVec_hitReq_11_207;
  assign compressDataVec_hitReq_11_207 = _GEN_502;
  wire          _GEN_503 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'hF;
  wire          compressDataVec_hitReq_12_15;
  assign compressDataVec_hitReq_12_15 = _GEN_503;
  wire          compressDataVec_hitReq_12_143;
  assign compressDataVec_hitReq_12_143 = _GEN_503;
  wire          compressDataVec_hitReq_12_207;
  assign compressDataVec_hitReq_12_207 = _GEN_503;
  wire          _GEN_504 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'hF;
  wire          compressDataVec_hitReq_13_15;
  assign compressDataVec_hitReq_13_15 = _GEN_504;
  wire          compressDataVec_hitReq_13_143;
  assign compressDataVec_hitReq_13_143 = _GEN_504;
  wire          compressDataVec_hitReq_13_207;
  assign compressDataVec_hitReq_13_207 = _GEN_504;
  wire          _GEN_505 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'hF;
  wire          compressDataVec_hitReq_14_15;
  assign compressDataVec_hitReq_14_15 = _GEN_505;
  wire          compressDataVec_hitReq_14_143;
  assign compressDataVec_hitReq_14_143 = _GEN_505;
  wire          compressDataVec_hitReq_14_207;
  assign compressDataVec_hitReq_14_207 = _GEN_505;
  wire          _GEN_506 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'hF;
  wire          compressDataVec_hitReq_15_15;
  assign compressDataVec_hitReq_15_15 = _GEN_506;
  wire          compressDataVec_hitReq_15_143;
  assign compressDataVec_hitReq_15_143 = _GEN_506;
  wire          compressDataVec_hitReq_15_207;
  assign compressDataVec_hitReq_15_207 = _GEN_506;
  wire          _GEN_507 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'hF;
  wire          compressDataVec_hitReq_16_15;
  assign compressDataVec_hitReq_16_15 = _GEN_507;
  wire          compressDataVec_hitReq_16_143;
  assign compressDataVec_hitReq_16_143 = _GEN_507;
  wire          _GEN_508 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'hF;
  wire          compressDataVec_hitReq_17_15;
  assign compressDataVec_hitReq_17_15 = _GEN_508;
  wire          compressDataVec_hitReq_17_143;
  assign compressDataVec_hitReq_17_143 = _GEN_508;
  wire          _GEN_509 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'hF;
  wire          compressDataVec_hitReq_18_15;
  assign compressDataVec_hitReq_18_15 = _GEN_509;
  wire          compressDataVec_hitReq_18_143;
  assign compressDataVec_hitReq_18_143 = _GEN_509;
  wire          _GEN_510 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'hF;
  wire          compressDataVec_hitReq_19_15;
  assign compressDataVec_hitReq_19_15 = _GEN_510;
  wire          compressDataVec_hitReq_19_143;
  assign compressDataVec_hitReq_19_143 = _GEN_510;
  wire          _GEN_511 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'hF;
  wire          compressDataVec_hitReq_20_15;
  assign compressDataVec_hitReq_20_15 = _GEN_511;
  wire          compressDataVec_hitReq_20_143;
  assign compressDataVec_hitReq_20_143 = _GEN_511;
  wire          _GEN_512 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'hF;
  wire          compressDataVec_hitReq_21_15;
  assign compressDataVec_hitReq_21_15 = _GEN_512;
  wire          compressDataVec_hitReq_21_143;
  assign compressDataVec_hitReq_21_143 = _GEN_512;
  wire          _GEN_513 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'hF;
  wire          compressDataVec_hitReq_22_15;
  assign compressDataVec_hitReq_22_15 = _GEN_513;
  wire          compressDataVec_hitReq_22_143;
  assign compressDataVec_hitReq_22_143 = _GEN_513;
  wire          _GEN_514 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'hF;
  wire          compressDataVec_hitReq_23_15;
  assign compressDataVec_hitReq_23_15 = _GEN_514;
  wire          compressDataVec_hitReq_23_143;
  assign compressDataVec_hitReq_23_143 = _GEN_514;
  wire          _GEN_515 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'hF;
  wire          compressDataVec_hitReq_24_15;
  assign compressDataVec_hitReq_24_15 = _GEN_515;
  wire          compressDataVec_hitReq_24_143;
  assign compressDataVec_hitReq_24_143 = _GEN_515;
  wire          _GEN_516 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'hF;
  wire          compressDataVec_hitReq_25_15;
  assign compressDataVec_hitReq_25_15 = _GEN_516;
  wire          compressDataVec_hitReq_25_143;
  assign compressDataVec_hitReq_25_143 = _GEN_516;
  wire          _GEN_517 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'hF;
  wire          compressDataVec_hitReq_26_15;
  assign compressDataVec_hitReq_26_15 = _GEN_517;
  wire          compressDataVec_hitReq_26_143;
  assign compressDataVec_hitReq_26_143 = _GEN_517;
  wire          _GEN_518 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'hF;
  wire          compressDataVec_hitReq_27_15;
  assign compressDataVec_hitReq_27_15 = _GEN_518;
  wire          compressDataVec_hitReq_27_143;
  assign compressDataVec_hitReq_27_143 = _GEN_518;
  wire          _GEN_519 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'hF;
  wire          compressDataVec_hitReq_28_15;
  assign compressDataVec_hitReq_28_15 = _GEN_519;
  wire          compressDataVec_hitReq_28_143;
  assign compressDataVec_hitReq_28_143 = _GEN_519;
  wire          _GEN_520 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'hF;
  wire          compressDataVec_hitReq_29_15;
  assign compressDataVec_hitReq_29_15 = _GEN_520;
  wire          compressDataVec_hitReq_29_143;
  assign compressDataVec_hitReq_29_143 = _GEN_520;
  wire          _GEN_521 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'hF;
  wire          compressDataVec_hitReq_30_15;
  assign compressDataVec_hitReq_30_15 = _GEN_521;
  wire          compressDataVec_hitReq_30_143;
  assign compressDataVec_hitReq_30_143 = _GEN_521;
  wire          _GEN_522 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'hF;
  wire          compressDataVec_hitReq_31_15;
  assign compressDataVec_hitReq_31_15 = _GEN_522;
  wire          compressDataVec_hitReq_31_143;
  assign compressDataVec_hitReq_31_143 = _GEN_522;
  wire          compressDataVec_hitReq_32_15 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'hF;
  wire          compressDataVec_hitReq_33_15 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'hF;
  wire          compressDataVec_hitReq_34_15 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'hF;
  wire          compressDataVec_hitReq_35_15 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'hF;
  wire          compressDataVec_hitReq_36_15 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'hF;
  wire          compressDataVec_hitReq_37_15 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'hF;
  wire          compressDataVec_hitReq_38_15 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'hF;
  wire          compressDataVec_hitReq_39_15 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'hF;
  wire          compressDataVec_hitReq_40_15 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'hF;
  wire          compressDataVec_hitReq_41_15 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'hF;
  wire          compressDataVec_hitReq_42_15 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'hF;
  wire          compressDataVec_hitReq_43_15 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'hF;
  wire          compressDataVec_hitReq_44_15 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'hF;
  wire          compressDataVec_hitReq_45_15 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'hF;
  wire          compressDataVec_hitReq_46_15 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'hF;
  wire          compressDataVec_hitReq_47_15 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'hF;
  wire          compressDataVec_hitReq_48_15 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'hF;
  wire          compressDataVec_hitReq_49_15 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'hF;
  wire          compressDataVec_hitReq_50_15 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'hF;
  wire          compressDataVec_hitReq_51_15 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'hF;
  wire          compressDataVec_hitReq_52_15 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'hF;
  wire          compressDataVec_hitReq_53_15 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'hF;
  wire          compressDataVec_hitReq_54_15 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'hF;
  wire          compressDataVec_hitReq_55_15 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'hF;
  wire          compressDataVec_hitReq_56_15 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'hF;
  wire          compressDataVec_hitReq_57_15 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'hF;
  wire          compressDataVec_hitReq_58_15 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'hF;
  wire          compressDataVec_hitReq_59_15 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'hF;
  wire          compressDataVec_hitReq_60_15 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'hF;
  wire          compressDataVec_hitReq_61_15 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'hF;
  wire          compressDataVec_hitReq_62_15 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'hF;
  wire          compressDataVec_hitReq_63_15 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'hF;
  wire [7:0]    compressDataVec_selectReqData_15 =
    (compressDataVec_hitReq_0_15 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_15 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_15 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_15 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_15 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_15 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_15 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_15 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_15 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_15 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_15 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_15 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_15 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_15 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_15 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_15 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_15 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_15 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_15 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_15 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_15 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_15 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_15 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_15 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_15 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_15 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_15 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_15 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_15 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_15 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_15 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_15 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_15 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_15 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_15 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_15 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_15 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_15 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_15 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_15 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_15 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_15 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_15 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_15 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_15 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_15 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_15 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_15 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_15 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_15 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_15 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_15 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_15 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_15 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_15 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_15 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_15 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_15 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_15 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_15 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_15 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_15 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_15 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_15 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_15;
  assign compressDataVec_useTail_15 = |(tailCount[5:4]);
  wire          _GEN_523 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h10;
  wire          compressDataVec_hitReq_0_16;
  assign compressDataVec_hitReq_0_16 = _GEN_523;
  wire          compressDataVec_hitReq_0_144;
  assign compressDataVec_hitReq_0_144 = _GEN_523;
  wire          compressDataVec_hitReq_0_208;
  assign compressDataVec_hitReq_0_208 = _GEN_523;
  wire          _GEN_524 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h10;
  wire          compressDataVec_hitReq_1_16;
  assign compressDataVec_hitReq_1_16 = _GEN_524;
  wire          compressDataVec_hitReq_1_144;
  assign compressDataVec_hitReq_1_144 = _GEN_524;
  wire          compressDataVec_hitReq_1_208;
  assign compressDataVec_hitReq_1_208 = _GEN_524;
  wire          _GEN_525 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h10;
  wire          compressDataVec_hitReq_2_16;
  assign compressDataVec_hitReq_2_16 = _GEN_525;
  wire          compressDataVec_hitReq_2_144;
  assign compressDataVec_hitReq_2_144 = _GEN_525;
  wire          compressDataVec_hitReq_2_208;
  assign compressDataVec_hitReq_2_208 = _GEN_525;
  wire          _GEN_526 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h10;
  wire          compressDataVec_hitReq_3_16;
  assign compressDataVec_hitReq_3_16 = _GEN_526;
  wire          compressDataVec_hitReq_3_144;
  assign compressDataVec_hitReq_3_144 = _GEN_526;
  wire          compressDataVec_hitReq_3_208;
  assign compressDataVec_hitReq_3_208 = _GEN_526;
  wire          _GEN_527 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h10;
  wire          compressDataVec_hitReq_4_16;
  assign compressDataVec_hitReq_4_16 = _GEN_527;
  wire          compressDataVec_hitReq_4_144;
  assign compressDataVec_hitReq_4_144 = _GEN_527;
  wire          compressDataVec_hitReq_4_208;
  assign compressDataVec_hitReq_4_208 = _GEN_527;
  wire          _GEN_528 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h10;
  wire          compressDataVec_hitReq_5_16;
  assign compressDataVec_hitReq_5_16 = _GEN_528;
  wire          compressDataVec_hitReq_5_144;
  assign compressDataVec_hitReq_5_144 = _GEN_528;
  wire          compressDataVec_hitReq_5_208;
  assign compressDataVec_hitReq_5_208 = _GEN_528;
  wire          _GEN_529 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h10;
  wire          compressDataVec_hitReq_6_16;
  assign compressDataVec_hitReq_6_16 = _GEN_529;
  wire          compressDataVec_hitReq_6_144;
  assign compressDataVec_hitReq_6_144 = _GEN_529;
  wire          compressDataVec_hitReq_6_208;
  assign compressDataVec_hitReq_6_208 = _GEN_529;
  wire          _GEN_530 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h10;
  wire          compressDataVec_hitReq_7_16;
  assign compressDataVec_hitReq_7_16 = _GEN_530;
  wire          compressDataVec_hitReq_7_144;
  assign compressDataVec_hitReq_7_144 = _GEN_530;
  wire          compressDataVec_hitReq_7_208;
  assign compressDataVec_hitReq_7_208 = _GEN_530;
  wire          _GEN_531 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h10;
  wire          compressDataVec_hitReq_8_16;
  assign compressDataVec_hitReq_8_16 = _GEN_531;
  wire          compressDataVec_hitReq_8_144;
  assign compressDataVec_hitReq_8_144 = _GEN_531;
  wire          compressDataVec_hitReq_8_208;
  assign compressDataVec_hitReq_8_208 = _GEN_531;
  wire          _GEN_532 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h10;
  wire          compressDataVec_hitReq_9_16;
  assign compressDataVec_hitReq_9_16 = _GEN_532;
  wire          compressDataVec_hitReq_9_144;
  assign compressDataVec_hitReq_9_144 = _GEN_532;
  wire          compressDataVec_hitReq_9_208;
  assign compressDataVec_hitReq_9_208 = _GEN_532;
  wire          _GEN_533 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h10;
  wire          compressDataVec_hitReq_10_16;
  assign compressDataVec_hitReq_10_16 = _GEN_533;
  wire          compressDataVec_hitReq_10_144;
  assign compressDataVec_hitReq_10_144 = _GEN_533;
  wire          compressDataVec_hitReq_10_208;
  assign compressDataVec_hitReq_10_208 = _GEN_533;
  wire          _GEN_534 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h10;
  wire          compressDataVec_hitReq_11_16;
  assign compressDataVec_hitReq_11_16 = _GEN_534;
  wire          compressDataVec_hitReq_11_144;
  assign compressDataVec_hitReq_11_144 = _GEN_534;
  wire          compressDataVec_hitReq_11_208;
  assign compressDataVec_hitReq_11_208 = _GEN_534;
  wire          _GEN_535 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h10;
  wire          compressDataVec_hitReq_12_16;
  assign compressDataVec_hitReq_12_16 = _GEN_535;
  wire          compressDataVec_hitReq_12_144;
  assign compressDataVec_hitReq_12_144 = _GEN_535;
  wire          compressDataVec_hitReq_12_208;
  assign compressDataVec_hitReq_12_208 = _GEN_535;
  wire          _GEN_536 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h10;
  wire          compressDataVec_hitReq_13_16;
  assign compressDataVec_hitReq_13_16 = _GEN_536;
  wire          compressDataVec_hitReq_13_144;
  assign compressDataVec_hitReq_13_144 = _GEN_536;
  wire          compressDataVec_hitReq_13_208;
  assign compressDataVec_hitReq_13_208 = _GEN_536;
  wire          _GEN_537 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h10;
  wire          compressDataVec_hitReq_14_16;
  assign compressDataVec_hitReq_14_16 = _GEN_537;
  wire          compressDataVec_hitReq_14_144;
  assign compressDataVec_hitReq_14_144 = _GEN_537;
  wire          compressDataVec_hitReq_14_208;
  assign compressDataVec_hitReq_14_208 = _GEN_537;
  wire          _GEN_538 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h10;
  wire          compressDataVec_hitReq_15_16;
  assign compressDataVec_hitReq_15_16 = _GEN_538;
  wire          compressDataVec_hitReq_15_144;
  assign compressDataVec_hitReq_15_144 = _GEN_538;
  wire          compressDataVec_hitReq_15_208;
  assign compressDataVec_hitReq_15_208 = _GEN_538;
  wire          _GEN_539 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h10;
  wire          compressDataVec_hitReq_16_16;
  assign compressDataVec_hitReq_16_16 = _GEN_539;
  wire          compressDataVec_hitReq_16_144;
  assign compressDataVec_hitReq_16_144 = _GEN_539;
  wire          _GEN_540 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h10;
  wire          compressDataVec_hitReq_17_16;
  assign compressDataVec_hitReq_17_16 = _GEN_540;
  wire          compressDataVec_hitReq_17_144;
  assign compressDataVec_hitReq_17_144 = _GEN_540;
  wire          _GEN_541 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h10;
  wire          compressDataVec_hitReq_18_16;
  assign compressDataVec_hitReq_18_16 = _GEN_541;
  wire          compressDataVec_hitReq_18_144;
  assign compressDataVec_hitReq_18_144 = _GEN_541;
  wire          _GEN_542 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h10;
  wire          compressDataVec_hitReq_19_16;
  assign compressDataVec_hitReq_19_16 = _GEN_542;
  wire          compressDataVec_hitReq_19_144;
  assign compressDataVec_hitReq_19_144 = _GEN_542;
  wire          _GEN_543 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h10;
  wire          compressDataVec_hitReq_20_16;
  assign compressDataVec_hitReq_20_16 = _GEN_543;
  wire          compressDataVec_hitReq_20_144;
  assign compressDataVec_hitReq_20_144 = _GEN_543;
  wire          _GEN_544 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h10;
  wire          compressDataVec_hitReq_21_16;
  assign compressDataVec_hitReq_21_16 = _GEN_544;
  wire          compressDataVec_hitReq_21_144;
  assign compressDataVec_hitReq_21_144 = _GEN_544;
  wire          _GEN_545 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h10;
  wire          compressDataVec_hitReq_22_16;
  assign compressDataVec_hitReq_22_16 = _GEN_545;
  wire          compressDataVec_hitReq_22_144;
  assign compressDataVec_hitReq_22_144 = _GEN_545;
  wire          _GEN_546 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h10;
  wire          compressDataVec_hitReq_23_16;
  assign compressDataVec_hitReq_23_16 = _GEN_546;
  wire          compressDataVec_hitReq_23_144;
  assign compressDataVec_hitReq_23_144 = _GEN_546;
  wire          _GEN_547 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h10;
  wire          compressDataVec_hitReq_24_16;
  assign compressDataVec_hitReq_24_16 = _GEN_547;
  wire          compressDataVec_hitReq_24_144;
  assign compressDataVec_hitReq_24_144 = _GEN_547;
  wire          _GEN_548 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h10;
  wire          compressDataVec_hitReq_25_16;
  assign compressDataVec_hitReq_25_16 = _GEN_548;
  wire          compressDataVec_hitReq_25_144;
  assign compressDataVec_hitReq_25_144 = _GEN_548;
  wire          _GEN_549 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h10;
  wire          compressDataVec_hitReq_26_16;
  assign compressDataVec_hitReq_26_16 = _GEN_549;
  wire          compressDataVec_hitReq_26_144;
  assign compressDataVec_hitReq_26_144 = _GEN_549;
  wire          _GEN_550 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h10;
  wire          compressDataVec_hitReq_27_16;
  assign compressDataVec_hitReq_27_16 = _GEN_550;
  wire          compressDataVec_hitReq_27_144;
  assign compressDataVec_hitReq_27_144 = _GEN_550;
  wire          _GEN_551 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h10;
  wire          compressDataVec_hitReq_28_16;
  assign compressDataVec_hitReq_28_16 = _GEN_551;
  wire          compressDataVec_hitReq_28_144;
  assign compressDataVec_hitReq_28_144 = _GEN_551;
  wire          _GEN_552 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h10;
  wire          compressDataVec_hitReq_29_16;
  assign compressDataVec_hitReq_29_16 = _GEN_552;
  wire          compressDataVec_hitReq_29_144;
  assign compressDataVec_hitReq_29_144 = _GEN_552;
  wire          _GEN_553 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h10;
  wire          compressDataVec_hitReq_30_16;
  assign compressDataVec_hitReq_30_16 = _GEN_553;
  wire          compressDataVec_hitReq_30_144;
  assign compressDataVec_hitReq_30_144 = _GEN_553;
  wire          _GEN_554 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h10;
  wire          compressDataVec_hitReq_31_16;
  assign compressDataVec_hitReq_31_16 = _GEN_554;
  wire          compressDataVec_hitReq_31_144;
  assign compressDataVec_hitReq_31_144 = _GEN_554;
  wire          compressDataVec_hitReq_32_16 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h10;
  wire          compressDataVec_hitReq_33_16 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h10;
  wire          compressDataVec_hitReq_34_16 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h10;
  wire          compressDataVec_hitReq_35_16 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h10;
  wire          compressDataVec_hitReq_36_16 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h10;
  wire          compressDataVec_hitReq_37_16 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h10;
  wire          compressDataVec_hitReq_38_16 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h10;
  wire          compressDataVec_hitReq_39_16 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h10;
  wire          compressDataVec_hitReq_40_16 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h10;
  wire          compressDataVec_hitReq_41_16 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h10;
  wire          compressDataVec_hitReq_42_16 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h10;
  wire          compressDataVec_hitReq_43_16 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h10;
  wire          compressDataVec_hitReq_44_16 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h10;
  wire          compressDataVec_hitReq_45_16 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h10;
  wire          compressDataVec_hitReq_46_16 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h10;
  wire          compressDataVec_hitReq_47_16 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h10;
  wire          compressDataVec_hitReq_48_16 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h10;
  wire          compressDataVec_hitReq_49_16 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h10;
  wire          compressDataVec_hitReq_50_16 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h10;
  wire          compressDataVec_hitReq_51_16 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h10;
  wire          compressDataVec_hitReq_52_16 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h10;
  wire          compressDataVec_hitReq_53_16 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h10;
  wire          compressDataVec_hitReq_54_16 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h10;
  wire          compressDataVec_hitReq_55_16 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h10;
  wire          compressDataVec_hitReq_56_16 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h10;
  wire          compressDataVec_hitReq_57_16 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h10;
  wire          compressDataVec_hitReq_58_16 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h10;
  wire          compressDataVec_hitReq_59_16 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h10;
  wire          compressDataVec_hitReq_60_16 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h10;
  wire          compressDataVec_hitReq_61_16 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h10;
  wire          compressDataVec_hitReq_62_16 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h10;
  wire          compressDataVec_hitReq_63_16 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h10;
  wire [7:0]    compressDataVec_selectReqData_16 =
    (compressDataVec_hitReq_0_16 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_16 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_16 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_16 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_16 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_16 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_16 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_16 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_16 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_16 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_16 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_16 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_16 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_16 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_16 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_16 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_16 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_16 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_16 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_16 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_16 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_16 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_16 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_16 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_16 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_16 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_16 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_16 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_16 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_16 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_16 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_16 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_16 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_16 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_16 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_16 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_16 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_16 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_16 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_16 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_16 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_16 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_16 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_16 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_16 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_16 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_16 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_16 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_16 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_16 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_16 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_16 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_16 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_16 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_16 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_16 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_16 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_16 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_16 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_16 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_16 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_16 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_16 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_16 ? source2Pipe[511:504] : 8'h0);
  wire          _GEN_555 = tailCount > 6'h10;
  wire          compressDataVec_useTail_16;
  assign compressDataVec_useTail_16 = _GEN_555;
  wire          compressDataVec_useTail_80;
  assign compressDataVec_useTail_80 = _GEN_555;
  wire          _GEN_556 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h11;
  wire          compressDataVec_hitReq_0_17;
  assign compressDataVec_hitReq_0_17 = _GEN_556;
  wire          compressDataVec_hitReq_0_145;
  assign compressDataVec_hitReq_0_145 = _GEN_556;
  wire          compressDataVec_hitReq_0_209;
  assign compressDataVec_hitReq_0_209 = _GEN_556;
  wire          _GEN_557 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h11;
  wire          compressDataVec_hitReq_1_17;
  assign compressDataVec_hitReq_1_17 = _GEN_557;
  wire          compressDataVec_hitReq_1_145;
  assign compressDataVec_hitReq_1_145 = _GEN_557;
  wire          compressDataVec_hitReq_1_209;
  assign compressDataVec_hitReq_1_209 = _GEN_557;
  wire          _GEN_558 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h11;
  wire          compressDataVec_hitReq_2_17;
  assign compressDataVec_hitReq_2_17 = _GEN_558;
  wire          compressDataVec_hitReq_2_145;
  assign compressDataVec_hitReq_2_145 = _GEN_558;
  wire          compressDataVec_hitReq_2_209;
  assign compressDataVec_hitReq_2_209 = _GEN_558;
  wire          _GEN_559 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h11;
  wire          compressDataVec_hitReq_3_17;
  assign compressDataVec_hitReq_3_17 = _GEN_559;
  wire          compressDataVec_hitReq_3_145;
  assign compressDataVec_hitReq_3_145 = _GEN_559;
  wire          compressDataVec_hitReq_3_209;
  assign compressDataVec_hitReq_3_209 = _GEN_559;
  wire          _GEN_560 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h11;
  wire          compressDataVec_hitReq_4_17;
  assign compressDataVec_hitReq_4_17 = _GEN_560;
  wire          compressDataVec_hitReq_4_145;
  assign compressDataVec_hitReq_4_145 = _GEN_560;
  wire          compressDataVec_hitReq_4_209;
  assign compressDataVec_hitReq_4_209 = _GEN_560;
  wire          _GEN_561 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h11;
  wire          compressDataVec_hitReq_5_17;
  assign compressDataVec_hitReq_5_17 = _GEN_561;
  wire          compressDataVec_hitReq_5_145;
  assign compressDataVec_hitReq_5_145 = _GEN_561;
  wire          compressDataVec_hitReq_5_209;
  assign compressDataVec_hitReq_5_209 = _GEN_561;
  wire          _GEN_562 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h11;
  wire          compressDataVec_hitReq_6_17;
  assign compressDataVec_hitReq_6_17 = _GEN_562;
  wire          compressDataVec_hitReq_6_145;
  assign compressDataVec_hitReq_6_145 = _GEN_562;
  wire          compressDataVec_hitReq_6_209;
  assign compressDataVec_hitReq_6_209 = _GEN_562;
  wire          _GEN_563 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h11;
  wire          compressDataVec_hitReq_7_17;
  assign compressDataVec_hitReq_7_17 = _GEN_563;
  wire          compressDataVec_hitReq_7_145;
  assign compressDataVec_hitReq_7_145 = _GEN_563;
  wire          compressDataVec_hitReq_7_209;
  assign compressDataVec_hitReq_7_209 = _GEN_563;
  wire          _GEN_564 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h11;
  wire          compressDataVec_hitReq_8_17;
  assign compressDataVec_hitReq_8_17 = _GEN_564;
  wire          compressDataVec_hitReq_8_145;
  assign compressDataVec_hitReq_8_145 = _GEN_564;
  wire          compressDataVec_hitReq_8_209;
  assign compressDataVec_hitReq_8_209 = _GEN_564;
  wire          _GEN_565 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h11;
  wire          compressDataVec_hitReq_9_17;
  assign compressDataVec_hitReq_9_17 = _GEN_565;
  wire          compressDataVec_hitReq_9_145;
  assign compressDataVec_hitReq_9_145 = _GEN_565;
  wire          compressDataVec_hitReq_9_209;
  assign compressDataVec_hitReq_9_209 = _GEN_565;
  wire          _GEN_566 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h11;
  wire          compressDataVec_hitReq_10_17;
  assign compressDataVec_hitReq_10_17 = _GEN_566;
  wire          compressDataVec_hitReq_10_145;
  assign compressDataVec_hitReq_10_145 = _GEN_566;
  wire          compressDataVec_hitReq_10_209;
  assign compressDataVec_hitReq_10_209 = _GEN_566;
  wire          _GEN_567 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h11;
  wire          compressDataVec_hitReq_11_17;
  assign compressDataVec_hitReq_11_17 = _GEN_567;
  wire          compressDataVec_hitReq_11_145;
  assign compressDataVec_hitReq_11_145 = _GEN_567;
  wire          compressDataVec_hitReq_11_209;
  assign compressDataVec_hitReq_11_209 = _GEN_567;
  wire          _GEN_568 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h11;
  wire          compressDataVec_hitReq_12_17;
  assign compressDataVec_hitReq_12_17 = _GEN_568;
  wire          compressDataVec_hitReq_12_145;
  assign compressDataVec_hitReq_12_145 = _GEN_568;
  wire          compressDataVec_hitReq_12_209;
  assign compressDataVec_hitReq_12_209 = _GEN_568;
  wire          _GEN_569 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h11;
  wire          compressDataVec_hitReq_13_17;
  assign compressDataVec_hitReq_13_17 = _GEN_569;
  wire          compressDataVec_hitReq_13_145;
  assign compressDataVec_hitReq_13_145 = _GEN_569;
  wire          compressDataVec_hitReq_13_209;
  assign compressDataVec_hitReq_13_209 = _GEN_569;
  wire          _GEN_570 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h11;
  wire          compressDataVec_hitReq_14_17;
  assign compressDataVec_hitReq_14_17 = _GEN_570;
  wire          compressDataVec_hitReq_14_145;
  assign compressDataVec_hitReq_14_145 = _GEN_570;
  wire          compressDataVec_hitReq_14_209;
  assign compressDataVec_hitReq_14_209 = _GEN_570;
  wire          _GEN_571 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h11;
  wire          compressDataVec_hitReq_15_17;
  assign compressDataVec_hitReq_15_17 = _GEN_571;
  wire          compressDataVec_hitReq_15_145;
  assign compressDataVec_hitReq_15_145 = _GEN_571;
  wire          compressDataVec_hitReq_15_209;
  assign compressDataVec_hitReq_15_209 = _GEN_571;
  wire          _GEN_572 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h11;
  wire          compressDataVec_hitReq_16_17;
  assign compressDataVec_hitReq_16_17 = _GEN_572;
  wire          compressDataVec_hitReq_16_145;
  assign compressDataVec_hitReq_16_145 = _GEN_572;
  wire          _GEN_573 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h11;
  wire          compressDataVec_hitReq_17_17;
  assign compressDataVec_hitReq_17_17 = _GEN_573;
  wire          compressDataVec_hitReq_17_145;
  assign compressDataVec_hitReq_17_145 = _GEN_573;
  wire          _GEN_574 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h11;
  wire          compressDataVec_hitReq_18_17;
  assign compressDataVec_hitReq_18_17 = _GEN_574;
  wire          compressDataVec_hitReq_18_145;
  assign compressDataVec_hitReq_18_145 = _GEN_574;
  wire          _GEN_575 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h11;
  wire          compressDataVec_hitReq_19_17;
  assign compressDataVec_hitReq_19_17 = _GEN_575;
  wire          compressDataVec_hitReq_19_145;
  assign compressDataVec_hitReq_19_145 = _GEN_575;
  wire          _GEN_576 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h11;
  wire          compressDataVec_hitReq_20_17;
  assign compressDataVec_hitReq_20_17 = _GEN_576;
  wire          compressDataVec_hitReq_20_145;
  assign compressDataVec_hitReq_20_145 = _GEN_576;
  wire          _GEN_577 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h11;
  wire          compressDataVec_hitReq_21_17;
  assign compressDataVec_hitReq_21_17 = _GEN_577;
  wire          compressDataVec_hitReq_21_145;
  assign compressDataVec_hitReq_21_145 = _GEN_577;
  wire          _GEN_578 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h11;
  wire          compressDataVec_hitReq_22_17;
  assign compressDataVec_hitReq_22_17 = _GEN_578;
  wire          compressDataVec_hitReq_22_145;
  assign compressDataVec_hitReq_22_145 = _GEN_578;
  wire          _GEN_579 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h11;
  wire          compressDataVec_hitReq_23_17;
  assign compressDataVec_hitReq_23_17 = _GEN_579;
  wire          compressDataVec_hitReq_23_145;
  assign compressDataVec_hitReq_23_145 = _GEN_579;
  wire          _GEN_580 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h11;
  wire          compressDataVec_hitReq_24_17;
  assign compressDataVec_hitReq_24_17 = _GEN_580;
  wire          compressDataVec_hitReq_24_145;
  assign compressDataVec_hitReq_24_145 = _GEN_580;
  wire          _GEN_581 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h11;
  wire          compressDataVec_hitReq_25_17;
  assign compressDataVec_hitReq_25_17 = _GEN_581;
  wire          compressDataVec_hitReq_25_145;
  assign compressDataVec_hitReq_25_145 = _GEN_581;
  wire          _GEN_582 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h11;
  wire          compressDataVec_hitReq_26_17;
  assign compressDataVec_hitReq_26_17 = _GEN_582;
  wire          compressDataVec_hitReq_26_145;
  assign compressDataVec_hitReq_26_145 = _GEN_582;
  wire          _GEN_583 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h11;
  wire          compressDataVec_hitReq_27_17;
  assign compressDataVec_hitReq_27_17 = _GEN_583;
  wire          compressDataVec_hitReq_27_145;
  assign compressDataVec_hitReq_27_145 = _GEN_583;
  wire          _GEN_584 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h11;
  wire          compressDataVec_hitReq_28_17;
  assign compressDataVec_hitReq_28_17 = _GEN_584;
  wire          compressDataVec_hitReq_28_145;
  assign compressDataVec_hitReq_28_145 = _GEN_584;
  wire          _GEN_585 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h11;
  wire          compressDataVec_hitReq_29_17;
  assign compressDataVec_hitReq_29_17 = _GEN_585;
  wire          compressDataVec_hitReq_29_145;
  assign compressDataVec_hitReq_29_145 = _GEN_585;
  wire          _GEN_586 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h11;
  wire          compressDataVec_hitReq_30_17;
  assign compressDataVec_hitReq_30_17 = _GEN_586;
  wire          compressDataVec_hitReq_30_145;
  assign compressDataVec_hitReq_30_145 = _GEN_586;
  wire          _GEN_587 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h11;
  wire          compressDataVec_hitReq_31_17;
  assign compressDataVec_hitReq_31_17 = _GEN_587;
  wire          compressDataVec_hitReq_31_145;
  assign compressDataVec_hitReq_31_145 = _GEN_587;
  wire          compressDataVec_hitReq_32_17 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h11;
  wire          compressDataVec_hitReq_33_17 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h11;
  wire          compressDataVec_hitReq_34_17 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h11;
  wire          compressDataVec_hitReq_35_17 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h11;
  wire          compressDataVec_hitReq_36_17 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h11;
  wire          compressDataVec_hitReq_37_17 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h11;
  wire          compressDataVec_hitReq_38_17 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h11;
  wire          compressDataVec_hitReq_39_17 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h11;
  wire          compressDataVec_hitReq_40_17 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h11;
  wire          compressDataVec_hitReq_41_17 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h11;
  wire          compressDataVec_hitReq_42_17 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h11;
  wire          compressDataVec_hitReq_43_17 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h11;
  wire          compressDataVec_hitReq_44_17 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h11;
  wire          compressDataVec_hitReq_45_17 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h11;
  wire          compressDataVec_hitReq_46_17 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h11;
  wire          compressDataVec_hitReq_47_17 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h11;
  wire          compressDataVec_hitReq_48_17 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h11;
  wire          compressDataVec_hitReq_49_17 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h11;
  wire          compressDataVec_hitReq_50_17 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h11;
  wire          compressDataVec_hitReq_51_17 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h11;
  wire          compressDataVec_hitReq_52_17 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h11;
  wire          compressDataVec_hitReq_53_17 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h11;
  wire          compressDataVec_hitReq_54_17 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h11;
  wire          compressDataVec_hitReq_55_17 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h11;
  wire          compressDataVec_hitReq_56_17 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h11;
  wire          compressDataVec_hitReq_57_17 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h11;
  wire          compressDataVec_hitReq_58_17 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h11;
  wire          compressDataVec_hitReq_59_17 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h11;
  wire          compressDataVec_hitReq_60_17 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h11;
  wire          compressDataVec_hitReq_61_17 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h11;
  wire          compressDataVec_hitReq_62_17 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h11;
  wire          compressDataVec_hitReq_63_17 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h11;
  wire [7:0]    compressDataVec_selectReqData_17 =
    (compressDataVec_hitReq_0_17 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_17 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_17 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_17 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_17 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_17 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_17 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_17 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_17 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_17 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_17 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_17 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_17 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_17 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_17 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_17 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_17 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_17 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_17 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_17 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_17 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_17 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_17 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_17 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_17 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_17 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_17 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_17 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_17 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_17 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_17 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_17 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_17 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_17 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_17 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_17 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_17 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_17 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_17 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_17 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_17 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_17 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_17 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_17 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_17 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_17 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_17 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_17 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_17 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_17 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_17 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_17 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_17 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_17 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_17 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_17 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_17 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_17 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_17 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_17 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_17 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_17 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_17 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_17 ? source2Pipe[511:504] : 8'h0);
  wire          _GEN_588 = tailCount > 6'h11;
  wire          compressDataVec_useTail_17;
  assign compressDataVec_useTail_17 = _GEN_588;
  wire          compressDataVec_useTail_81;
  assign compressDataVec_useTail_81 = _GEN_588;
  wire          _GEN_589 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h12;
  wire          compressDataVec_hitReq_0_18;
  assign compressDataVec_hitReq_0_18 = _GEN_589;
  wire          compressDataVec_hitReq_0_146;
  assign compressDataVec_hitReq_0_146 = _GEN_589;
  wire          compressDataVec_hitReq_0_210;
  assign compressDataVec_hitReq_0_210 = _GEN_589;
  wire          _GEN_590 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h12;
  wire          compressDataVec_hitReq_1_18;
  assign compressDataVec_hitReq_1_18 = _GEN_590;
  wire          compressDataVec_hitReq_1_146;
  assign compressDataVec_hitReq_1_146 = _GEN_590;
  wire          compressDataVec_hitReq_1_210;
  assign compressDataVec_hitReq_1_210 = _GEN_590;
  wire          _GEN_591 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h12;
  wire          compressDataVec_hitReq_2_18;
  assign compressDataVec_hitReq_2_18 = _GEN_591;
  wire          compressDataVec_hitReq_2_146;
  assign compressDataVec_hitReq_2_146 = _GEN_591;
  wire          compressDataVec_hitReq_2_210;
  assign compressDataVec_hitReq_2_210 = _GEN_591;
  wire          _GEN_592 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h12;
  wire          compressDataVec_hitReq_3_18;
  assign compressDataVec_hitReq_3_18 = _GEN_592;
  wire          compressDataVec_hitReq_3_146;
  assign compressDataVec_hitReq_3_146 = _GEN_592;
  wire          compressDataVec_hitReq_3_210;
  assign compressDataVec_hitReq_3_210 = _GEN_592;
  wire          _GEN_593 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h12;
  wire          compressDataVec_hitReq_4_18;
  assign compressDataVec_hitReq_4_18 = _GEN_593;
  wire          compressDataVec_hitReq_4_146;
  assign compressDataVec_hitReq_4_146 = _GEN_593;
  wire          compressDataVec_hitReq_4_210;
  assign compressDataVec_hitReq_4_210 = _GEN_593;
  wire          _GEN_594 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h12;
  wire          compressDataVec_hitReq_5_18;
  assign compressDataVec_hitReq_5_18 = _GEN_594;
  wire          compressDataVec_hitReq_5_146;
  assign compressDataVec_hitReq_5_146 = _GEN_594;
  wire          compressDataVec_hitReq_5_210;
  assign compressDataVec_hitReq_5_210 = _GEN_594;
  wire          _GEN_595 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h12;
  wire          compressDataVec_hitReq_6_18;
  assign compressDataVec_hitReq_6_18 = _GEN_595;
  wire          compressDataVec_hitReq_6_146;
  assign compressDataVec_hitReq_6_146 = _GEN_595;
  wire          compressDataVec_hitReq_6_210;
  assign compressDataVec_hitReq_6_210 = _GEN_595;
  wire          _GEN_596 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h12;
  wire          compressDataVec_hitReq_7_18;
  assign compressDataVec_hitReq_7_18 = _GEN_596;
  wire          compressDataVec_hitReq_7_146;
  assign compressDataVec_hitReq_7_146 = _GEN_596;
  wire          compressDataVec_hitReq_7_210;
  assign compressDataVec_hitReq_7_210 = _GEN_596;
  wire          _GEN_597 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h12;
  wire          compressDataVec_hitReq_8_18;
  assign compressDataVec_hitReq_8_18 = _GEN_597;
  wire          compressDataVec_hitReq_8_146;
  assign compressDataVec_hitReq_8_146 = _GEN_597;
  wire          compressDataVec_hitReq_8_210;
  assign compressDataVec_hitReq_8_210 = _GEN_597;
  wire          _GEN_598 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h12;
  wire          compressDataVec_hitReq_9_18;
  assign compressDataVec_hitReq_9_18 = _GEN_598;
  wire          compressDataVec_hitReq_9_146;
  assign compressDataVec_hitReq_9_146 = _GEN_598;
  wire          compressDataVec_hitReq_9_210;
  assign compressDataVec_hitReq_9_210 = _GEN_598;
  wire          _GEN_599 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h12;
  wire          compressDataVec_hitReq_10_18;
  assign compressDataVec_hitReq_10_18 = _GEN_599;
  wire          compressDataVec_hitReq_10_146;
  assign compressDataVec_hitReq_10_146 = _GEN_599;
  wire          compressDataVec_hitReq_10_210;
  assign compressDataVec_hitReq_10_210 = _GEN_599;
  wire          _GEN_600 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h12;
  wire          compressDataVec_hitReq_11_18;
  assign compressDataVec_hitReq_11_18 = _GEN_600;
  wire          compressDataVec_hitReq_11_146;
  assign compressDataVec_hitReq_11_146 = _GEN_600;
  wire          compressDataVec_hitReq_11_210;
  assign compressDataVec_hitReq_11_210 = _GEN_600;
  wire          _GEN_601 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h12;
  wire          compressDataVec_hitReq_12_18;
  assign compressDataVec_hitReq_12_18 = _GEN_601;
  wire          compressDataVec_hitReq_12_146;
  assign compressDataVec_hitReq_12_146 = _GEN_601;
  wire          compressDataVec_hitReq_12_210;
  assign compressDataVec_hitReq_12_210 = _GEN_601;
  wire          _GEN_602 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h12;
  wire          compressDataVec_hitReq_13_18;
  assign compressDataVec_hitReq_13_18 = _GEN_602;
  wire          compressDataVec_hitReq_13_146;
  assign compressDataVec_hitReq_13_146 = _GEN_602;
  wire          compressDataVec_hitReq_13_210;
  assign compressDataVec_hitReq_13_210 = _GEN_602;
  wire          _GEN_603 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h12;
  wire          compressDataVec_hitReq_14_18;
  assign compressDataVec_hitReq_14_18 = _GEN_603;
  wire          compressDataVec_hitReq_14_146;
  assign compressDataVec_hitReq_14_146 = _GEN_603;
  wire          compressDataVec_hitReq_14_210;
  assign compressDataVec_hitReq_14_210 = _GEN_603;
  wire          _GEN_604 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h12;
  wire          compressDataVec_hitReq_15_18;
  assign compressDataVec_hitReq_15_18 = _GEN_604;
  wire          compressDataVec_hitReq_15_146;
  assign compressDataVec_hitReq_15_146 = _GEN_604;
  wire          compressDataVec_hitReq_15_210;
  assign compressDataVec_hitReq_15_210 = _GEN_604;
  wire          _GEN_605 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h12;
  wire          compressDataVec_hitReq_16_18;
  assign compressDataVec_hitReq_16_18 = _GEN_605;
  wire          compressDataVec_hitReq_16_146;
  assign compressDataVec_hitReq_16_146 = _GEN_605;
  wire          _GEN_606 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h12;
  wire          compressDataVec_hitReq_17_18;
  assign compressDataVec_hitReq_17_18 = _GEN_606;
  wire          compressDataVec_hitReq_17_146;
  assign compressDataVec_hitReq_17_146 = _GEN_606;
  wire          _GEN_607 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h12;
  wire          compressDataVec_hitReq_18_18;
  assign compressDataVec_hitReq_18_18 = _GEN_607;
  wire          compressDataVec_hitReq_18_146;
  assign compressDataVec_hitReq_18_146 = _GEN_607;
  wire          _GEN_608 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h12;
  wire          compressDataVec_hitReq_19_18;
  assign compressDataVec_hitReq_19_18 = _GEN_608;
  wire          compressDataVec_hitReq_19_146;
  assign compressDataVec_hitReq_19_146 = _GEN_608;
  wire          _GEN_609 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h12;
  wire          compressDataVec_hitReq_20_18;
  assign compressDataVec_hitReq_20_18 = _GEN_609;
  wire          compressDataVec_hitReq_20_146;
  assign compressDataVec_hitReq_20_146 = _GEN_609;
  wire          _GEN_610 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h12;
  wire          compressDataVec_hitReq_21_18;
  assign compressDataVec_hitReq_21_18 = _GEN_610;
  wire          compressDataVec_hitReq_21_146;
  assign compressDataVec_hitReq_21_146 = _GEN_610;
  wire          _GEN_611 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h12;
  wire          compressDataVec_hitReq_22_18;
  assign compressDataVec_hitReq_22_18 = _GEN_611;
  wire          compressDataVec_hitReq_22_146;
  assign compressDataVec_hitReq_22_146 = _GEN_611;
  wire          _GEN_612 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h12;
  wire          compressDataVec_hitReq_23_18;
  assign compressDataVec_hitReq_23_18 = _GEN_612;
  wire          compressDataVec_hitReq_23_146;
  assign compressDataVec_hitReq_23_146 = _GEN_612;
  wire          _GEN_613 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h12;
  wire          compressDataVec_hitReq_24_18;
  assign compressDataVec_hitReq_24_18 = _GEN_613;
  wire          compressDataVec_hitReq_24_146;
  assign compressDataVec_hitReq_24_146 = _GEN_613;
  wire          _GEN_614 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h12;
  wire          compressDataVec_hitReq_25_18;
  assign compressDataVec_hitReq_25_18 = _GEN_614;
  wire          compressDataVec_hitReq_25_146;
  assign compressDataVec_hitReq_25_146 = _GEN_614;
  wire          _GEN_615 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h12;
  wire          compressDataVec_hitReq_26_18;
  assign compressDataVec_hitReq_26_18 = _GEN_615;
  wire          compressDataVec_hitReq_26_146;
  assign compressDataVec_hitReq_26_146 = _GEN_615;
  wire          _GEN_616 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h12;
  wire          compressDataVec_hitReq_27_18;
  assign compressDataVec_hitReq_27_18 = _GEN_616;
  wire          compressDataVec_hitReq_27_146;
  assign compressDataVec_hitReq_27_146 = _GEN_616;
  wire          _GEN_617 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h12;
  wire          compressDataVec_hitReq_28_18;
  assign compressDataVec_hitReq_28_18 = _GEN_617;
  wire          compressDataVec_hitReq_28_146;
  assign compressDataVec_hitReq_28_146 = _GEN_617;
  wire          _GEN_618 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h12;
  wire          compressDataVec_hitReq_29_18;
  assign compressDataVec_hitReq_29_18 = _GEN_618;
  wire          compressDataVec_hitReq_29_146;
  assign compressDataVec_hitReq_29_146 = _GEN_618;
  wire          _GEN_619 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h12;
  wire          compressDataVec_hitReq_30_18;
  assign compressDataVec_hitReq_30_18 = _GEN_619;
  wire          compressDataVec_hitReq_30_146;
  assign compressDataVec_hitReq_30_146 = _GEN_619;
  wire          _GEN_620 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h12;
  wire          compressDataVec_hitReq_31_18;
  assign compressDataVec_hitReq_31_18 = _GEN_620;
  wire          compressDataVec_hitReq_31_146;
  assign compressDataVec_hitReq_31_146 = _GEN_620;
  wire          compressDataVec_hitReq_32_18 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h12;
  wire          compressDataVec_hitReq_33_18 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h12;
  wire          compressDataVec_hitReq_34_18 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h12;
  wire          compressDataVec_hitReq_35_18 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h12;
  wire          compressDataVec_hitReq_36_18 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h12;
  wire          compressDataVec_hitReq_37_18 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h12;
  wire          compressDataVec_hitReq_38_18 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h12;
  wire          compressDataVec_hitReq_39_18 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h12;
  wire          compressDataVec_hitReq_40_18 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h12;
  wire          compressDataVec_hitReq_41_18 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h12;
  wire          compressDataVec_hitReq_42_18 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h12;
  wire          compressDataVec_hitReq_43_18 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h12;
  wire          compressDataVec_hitReq_44_18 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h12;
  wire          compressDataVec_hitReq_45_18 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h12;
  wire          compressDataVec_hitReq_46_18 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h12;
  wire          compressDataVec_hitReq_47_18 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h12;
  wire          compressDataVec_hitReq_48_18 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h12;
  wire          compressDataVec_hitReq_49_18 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h12;
  wire          compressDataVec_hitReq_50_18 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h12;
  wire          compressDataVec_hitReq_51_18 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h12;
  wire          compressDataVec_hitReq_52_18 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h12;
  wire          compressDataVec_hitReq_53_18 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h12;
  wire          compressDataVec_hitReq_54_18 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h12;
  wire          compressDataVec_hitReq_55_18 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h12;
  wire          compressDataVec_hitReq_56_18 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h12;
  wire          compressDataVec_hitReq_57_18 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h12;
  wire          compressDataVec_hitReq_58_18 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h12;
  wire          compressDataVec_hitReq_59_18 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h12;
  wire          compressDataVec_hitReq_60_18 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h12;
  wire          compressDataVec_hitReq_61_18 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h12;
  wire          compressDataVec_hitReq_62_18 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h12;
  wire          compressDataVec_hitReq_63_18 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h12;
  wire [7:0]    compressDataVec_selectReqData_18 =
    (compressDataVec_hitReq_0_18 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_18 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_18 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_18 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_18 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_18 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_18 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_18 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_18 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_18 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_18 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_18 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_18 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_18 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_18 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_18 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_18 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_18 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_18 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_18 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_18 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_18 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_18 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_18 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_18 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_18 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_18 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_18 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_18 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_18 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_18 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_18 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_18 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_18 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_18 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_18 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_18 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_18 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_18 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_18 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_18 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_18 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_18 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_18 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_18 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_18 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_18 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_18 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_18 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_18 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_18 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_18 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_18 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_18 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_18 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_18 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_18 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_18 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_18 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_18 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_18 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_18 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_18 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_18 ? source2Pipe[511:504] : 8'h0);
  wire          _GEN_621 = tailCount > 6'h12;
  wire          compressDataVec_useTail_18;
  assign compressDataVec_useTail_18 = _GEN_621;
  wire          compressDataVec_useTail_82;
  assign compressDataVec_useTail_82 = _GEN_621;
  wire          _GEN_622 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h13;
  wire          compressDataVec_hitReq_0_19;
  assign compressDataVec_hitReq_0_19 = _GEN_622;
  wire          compressDataVec_hitReq_0_147;
  assign compressDataVec_hitReq_0_147 = _GEN_622;
  wire          compressDataVec_hitReq_0_211;
  assign compressDataVec_hitReq_0_211 = _GEN_622;
  wire          _GEN_623 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h13;
  wire          compressDataVec_hitReq_1_19;
  assign compressDataVec_hitReq_1_19 = _GEN_623;
  wire          compressDataVec_hitReq_1_147;
  assign compressDataVec_hitReq_1_147 = _GEN_623;
  wire          compressDataVec_hitReq_1_211;
  assign compressDataVec_hitReq_1_211 = _GEN_623;
  wire          _GEN_624 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h13;
  wire          compressDataVec_hitReq_2_19;
  assign compressDataVec_hitReq_2_19 = _GEN_624;
  wire          compressDataVec_hitReq_2_147;
  assign compressDataVec_hitReq_2_147 = _GEN_624;
  wire          compressDataVec_hitReq_2_211;
  assign compressDataVec_hitReq_2_211 = _GEN_624;
  wire          _GEN_625 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h13;
  wire          compressDataVec_hitReq_3_19;
  assign compressDataVec_hitReq_3_19 = _GEN_625;
  wire          compressDataVec_hitReq_3_147;
  assign compressDataVec_hitReq_3_147 = _GEN_625;
  wire          compressDataVec_hitReq_3_211;
  assign compressDataVec_hitReq_3_211 = _GEN_625;
  wire          _GEN_626 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h13;
  wire          compressDataVec_hitReq_4_19;
  assign compressDataVec_hitReq_4_19 = _GEN_626;
  wire          compressDataVec_hitReq_4_147;
  assign compressDataVec_hitReq_4_147 = _GEN_626;
  wire          compressDataVec_hitReq_4_211;
  assign compressDataVec_hitReq_4_211 = _GEN_626;
  wire          _GEN_627 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h13;
  wire          compressDataVec_hitReq_5_19;
  assign compressDataVec_hitReq_5_19 = _GEN_627;
  wire          compressDataVec_hitReq_5_147;
  assign compressDataVec_hitReq_5_147 = _GEN_627;
  wire          compressDataVec_hitReq_5_211;
  assign compressDataVec_hitReq_5_211 = _GEN_627;
  wire          _GEN_628 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h13;
  wire          compressDataVec_hitReq_6_19;
  assign compressDataVec_hitReq_6_19 = _GEN_628;
  wire          compressDataVec_hitReq_6_147;
  assign compressDataVec_hitReq_6_147 = _GEN_628;
  wire          compressDataVec_hitReq_6_211;
  assign compressDataVec_hitReq_6_211 = _GEN_628;
  wire          _GEN_629 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h13;
  wire          compressDataVec_hitReq_7_19;
  assign compressDataVec_hitReq_7_19 = _GEN_629;
  wire          compressDataVec_hitReq_7_147;
  assign compressDataVec_hitReq_7_147 = _GEN_629;
  wire          compressDataVec_hitReq_7_211;
  assign compressDataVec_hitReq_7_211 = _GEN_629;
  wire          _GEN_630 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h13;
  wire          compressDataVec_hitReq_8_19;
  assign compressDataVec_hitReq_8_19 = _GEN_630;
  wire          compressDataVec_hitReq_8_147;
  assign compressDataVec_hitReq_8_147 = _GEN_630;
  wire          compressDataVec_hitReq_8_211;
  assign compressDataVec_hitReq_8_211 = _GEN_630;
  wire          _GEN_631 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h13;
  wire          compressDataVec_hitReq_9_19;
  assign compressDataVec_hitReq_9_19 = _GEN_631;
  wire          compressDataVec_hitReq_9_147;
  assign compressDataVec_hitReq_9_147 = _GEN_631;
  wire          compressDataVec_hitReq_9_211;
  assign compressDataVec_hitReq_9_211 = _GEN_631;
  wire          _GEN_632 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h13;
  wire          compressDataVec_hitReq_10_19;
  assign compressDataVec_hitReq_10_19 = _GEN_632;
  wire          compressDataVec_hitReq_10_147;
  assign compressDataVec_hitReq_10_147 = _GEN_632;
  wire          compressDataVec_hitReq_10_211;
  assign compressDataVec_hitReq_10_211 = _GEN_632;
  wire          _GEN_633 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h13;
  wire          compressDataVec_hitReq_11_19;
  assign compressDataVec_hitReq_11_19 = _GEN_633;
  wire          compressDataVec_hitReq_11_147;
  assign compressDataVec_hitReq_11_147 = _GEN_633;
  wire          compressDataVec_hitReq_11_211;
  assign compressDataVec_hitReq_11_211 = _GEN_633;
  wire          _GEN_634 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h13;
  wire          compressDataVec_hitReq_12_19;
  assign compressDataVec_hitReq_12_19 = _GEN_634;
  wire          compressDataVec_hitReq_12_147;
  assign compressDataVec_hitReq_12_147 = _GEN_634;
  wire          compressDataVec_hitReq_12_211;
  assign compressDataVec_hitReq_12_211 = _GEN_634;
  wire          _GEN_635 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h13;
  wire          compressDataVec_hitReq_13_19;
  assign compressDataVec_hitReq_13_19 = _GEN_635;
  wire          compressDataVec_hitReq_13_147;
  assign compressDataVec_hitReq_13_147 = _GEN_635;
  wire          compressDataVec_hitReq_13_211;
  assign compressDataVec_hitReq_13_211 = _GEN_635;
  wire          _GEN_636 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h13;
  wire          compressDataVec_hitReq_14_19;
  assign compressDataVec_hitReq_14_19 = _GEN_636;
  wire          compressDataVec_hitReq_14_147;
  assign compressDataVec_hitReq_14_147 = _GEN_636;
  wire          compressDataVec_hitReq_14_211;
  assign compressDataVec_hitReq_14_211 = _GEN_636;
  wire          _GEN_637 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h13;
  wire          compressDataVec_hitReq_15_19;
  assign compressDataVec_hitReq_15_19 = _GEN_637;
  wire          compressDataVec_hitReq_15_147;
  assign compressDataVec_hitReq_15_147 = _GEN_637;
  wire          compressDataVec_hitReq_15_211;
  assign compressDataVec_hitReq_15_211 = _GEN_637;
  wire          _GEN_638 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h13;
  wire          compressDataVec_hitReq_16_19;
  assign compressDataVec_hitReq_16_19 = _GEN_638;
  wire          compressDataVec_hitReq_16_147;
  assign compressDataVec_hitReq_16_147 = _GEN_638;
  wire          _GEN_639 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h13;
  wire          compressDataVec_hitReq_17_19;
  assign compressDataVec_hitReq_17_19 = _GEN_639;
  wire          compressDataVec_hitReq_17_147;
  assign compressDataVec_hitReq_17_147 = _GEN_639;
  wire          _GEN_640 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h13;
  wire          compressDataVec_hitReq_18_19;
  assign compressDataVec_hitReq_18_19 = _GEN_640;
  wire          compressDataVec_hitReq_18_147;
  assign compressDataVec_hitReq_18_147 = _GEN_640;
  wire          _GEN_641 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h13;
  wire          compressDataVec_hitReq_19_19;
  assign compressDataVec_hitReq_19_19 = _GEN_641;
  wire          compressDataVec_hitReq_19_147;
  assign compressDataVec_hitReq_19_147 = _GEN_641;
  wire          _GEN_642 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h13;
  wire          compressDataVec_hitReq_20_19;
  assign compressDataVec_hitReq_20_19 = _GEN_642;
  wire          compressDataVec_hitReq_20_147;
  assign compressDataVec_hitReq_20_147 = _GEN_642;
  wire          _GEN_643 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h13;
  wire          compressDataVec_hitReq_21_19;
  assign compressDataVec_hitReq_21_19 = _GEN_643;
  wire          compressDataVec_hitReq_21_147;
  assign compressDataVec_hitReq_21_147 = _GEN_643;
  wire          _GEN_644 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h13;
  wire          compressDataVec_hitReq_22_19;
  assign compressDataVec_hitReq_22_19 = _GEN_644;
  wire          compressDataVec_hitReq_22_147;
  assign compressDataVec_hitReq_22_147 = _GEN_644;
  wire          _GEN_645 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h13;
  wire          compressDataVec_hitReq_23_19;
  assign compressDataVec_hitReq_23_19 = _GEN_645;
  wire          compressDataVec_hitReq_23_147;
  assign compressDataVec_hitReq_23_147 = _GEN_645;
  wire          _GEN_646 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h13;
  wire          compressDataVec_hitReq_24_19;
  assign compressDataVec_hitReq_24_19 = _GEN_646;
  wire          compressDataVec_hitReq_24_147;
  assign compressDataVec_hitReq_24_147 = _GEN_646;
  wire          _GEN_647 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h13;
  wire          compressDataVec_hitReq_25_19;
  assign compressDataVec_hitReq_25_19 = _GEN_647;
  wire          compressDataVec_hitReq_25_147;
  assign compressDataVec_hitReq_25_147 = _GEN_647;
  wire          _GEN_648 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h13;
  wire          compressDataVec_hitReq_26_19;
  assign compressDataVec_hitReq_26_19 = _GEN_648;
  wire          compressDataVec_hitReq_26_147;
  assign compressDataVec_hitReq_26_147 = _GEN_648;
  wire          _GEN_649 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h13;
  wire          compressDataVec_hitReq_27_19;
  assign compressDataVec_hitReq_27_19 = _GEN_649;
  wire          compressDataVec_hitReq_27_147;
  assign compressDataVec_hitReq_27_147 = _GEN_649;
  wire          _GEN_650 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h13;
  wire          compressDataVec_hitReq_28_19;
  assign compressDataVec_hitReq_28_19 = _GEN_650;
  wire          compressDataVec_hitReq_28_147;
  assign compressDataVec_hitReq_28_147 = _GEN_650;
  wire          _GEN_651 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h13;
  wire          compressDataVec_hitReq_29_19;
  assign compressDataVec_hitReq_29_19 = _GEN_651;
  wire          compressDataVec_hitReq_29_147;
  assign compressDataVec_hitReq_29_147 = _GEN_651;
  wire          _GEN_652 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h13;
  wire          compressDataVec_hitReq_30_19;
  assign compressDataVec_hitReq_30_19 = _GEN_652;
  wire          compressDataVec_hitReq_30_147;
  assign compressDataVec_hitReq_30_147 = _GEN_652;
  wire          _GEN_653 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h13;
  wire          compressDataVec_hitReq_31_19;
  assign compressDataVec_hitReq_31_19 = _GEN_653;
  wire          compressDataVec_hitReq_31_147;
  assign compressDataVec_hitReq_31_147 = _GEN_653;
  wire          compressDataVec_hitReq_32_19 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h13;
  wire          compressDataVec_hitReq_33_19 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h13;
  wire          compressDataVec_hitReq_34_19 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h13;
  wire          compressDataVec_hitReq_35_19 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h13;
  wire          compressDataVec_hitReq_36_19 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h13;
  wire          compressDataVec_hitReq_37_19 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h13;
  wire          compressDataVec_hitReq_38_19 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h13;
  wire          compressDataVec_hitReq_39_19 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h13;
  wire          compressDataVec_hitReq_40_19 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h13;
  wire          compressDataVec_hitReq_41_19 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h13;
  wire          compressDataVec_hitReq_42_19 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h13;
  wire          compressDataVec_hitReq_43_19 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h13;
  wire          compressDataVec_hitReq_44_19 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h13;
  wire          compressDataVec_hitReq_45_19 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h13;
  wire          compressDataVec_hitReq_46_19 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h13;
  wire          compressDataVec_hitReq_47_19 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h13;
  wire          compressDataVec_hitReq_48_19 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h13;
  wire          compressDataVec_hitReq_49_19 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h13;
  wire          compressDataVec_hitReq_50_19 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h13;
  wire          compressDataVec_hitReq_51_19 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h13;
  wire          compressDataVec_hitReq_52_19 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h13;
  wire          compressDataVec_hitReq_53_19 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h13;
  wire          compressDataVec_hitReq_54_19 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h13;
  wire          compressDataVec_hitReq_55_19 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h13;
  wire          compressDataVec_hitReq_56_19 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h13;
  wire          compressDataVec_hitReq_57_19 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h13;
  wire          compressDataVec_hitReq_58_19 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h13;
  wire          compressDataVec_hitReq_59_19 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h13;
  wire          compressDataVec_hitReq_60_19 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h13;
  wire          compressDataVec_hitReq_61_19 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h13;
  wire          compressDataVec_hitReq_62_19 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h13;
  wire          compressDataVec_hitReq_63_19 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h13;
  wire [7:0]    compressDataVec_selectReqData_19 =
    (compressDataVec_hitReq_0_19 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_19 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_19 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_19 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_19 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_19 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_19 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_19 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_19 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_19 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_19 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_19 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_19 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_19 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_19 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_19 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_19 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_19 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_19 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_19 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_19 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_19 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_19 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_19 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_19 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_19 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_19 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_19 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_19 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_19 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_19 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_19 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_19 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_19 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_19 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_19 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_19 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_19 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_19 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_19 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_19 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_19 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_19 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_19 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_19 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_19 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_19 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_19 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_19 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_19 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_19 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_19 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_19 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_19 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_19 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_19 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_19 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_19 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_19 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_19 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_19 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_19 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_19 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_19 ? source2Pipe[511:504] : 8'h0);
  wire          _GEN_654 = tailCount > 6'h13;
  wire          compressDataVec_useTail_19;
  assign compressDataVec_useTail_19 = _GEN_654;
  wire          compressDataVec_useTail_83;
  assign compressDataVec_useTail_83 = _GEN_654;
  wire          _GEN_655 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h14;
  wire          compressDataVec_hitReq_0_20;
  assign compressDataVec_hitReq_0_20 = _GEN_655;
  wire          compressDataVec_hitReq_0_148;
  assign compressDataVec_hitReq_0_148 = _GEN_655;
  wire          compressDataVec_hitReq_0_212;
  assign compressDataVec_hitReq_0_212 = _GEN_655;
  wire          _GEN_656 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h14;
  wire          compressDataVec_hitReq_1_20;
  assign compressDataVec_hitReq_1_20 = _GEN_656;
  wire          compressDataVec_hitReq_1_148;
  assign compressDataVec_hitReq_1_148 = _GEN_656;
  wire          compressDataVec_hitReq_1_212;
  assign compressDataVec_hitReq_1_212 = _GEN_656;
  wire          _GEN_657 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h14;
  wire          compressDataVec_hitReq_2_20;
  assign compressDataVec_hitReq_2_20 = _GEN_657;
  wire          compressDataVec_hitReq_2_148;
  assign compressDataVec_hitReq_2_148 = _GEN_657;
  wire          compressDataVec_hitReq_2_212;
  assign compressDataVec_hitReq_2_212 = _GEN_657;
  wire          _GEN_658 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h14;
  wire          compressDataVec_hitReq_3_20;
  assign compressDataVec_hitReq_3_20 = _GEN_658;
  wire          compressDataVec_hitReq_3_148;
  assign compressDataVec_hitReq_3_148 = _GEN_658;
  wire          compressDataVec_hitReq_3_212;
  assign compressDataVec_hitReq_3_212 = _GEN_658;
  wire          _GEN_659 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h14;
  wire          compressDataVec_hitReq_4_20;
  assign compressDataVec_hitReq_4_20 = _GEN_659;
  wire          compressDataVec_hitReq_4_148;
  assign compressDataVec_hitReq_4_148 = _GEN_659;
  wire          compressDataVec_hitReq_4_212;
  assign compressDataVec_hitReq_4_212 = _GEN_659;
  wire          _GEN_660 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h14;
  wire          compressDataVec_hitReq_5_20;
  assign compressDataVec_hitReq_5_20 = _GEN_660;
  wire          compressDataVec_hitReq_5_148;
  assign compressDataVec_hitReq_5_148 = _GEN_660;
  wire          compressDataVec_hitReq_5_212;
  assign compressDataVec_hitReq_5_212 = _GEN_660;
  wire          _GEN_661 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h14;
  wire          compressDataVec_hitReq_6_20;
  assign compressDataVec_hitReq_6_20 = _GEN_661;
  wire          compressDataVec_hitReq_6_148;
  assign compressDataVec_hitReq_6_148 = _GEN_661;
  wire          compressDataVec_hitReq_6_212;
  assign compressDataVec_hitReq_6_212 = _GEN_661;
  wire          _GEN_662 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h14;
  wire          compressDataVec_hitReq_7_20;
  assign compressDataVec_hitReq_7_20 = _GEN_662;
  wire          compressDataVec_hitReq_7_148;
  assign compressDataVec_hitReq_7_148 = _GEN_662;
  wire          compressDataVec_hitReq_7_212;
  assign compressDataVec_hitReq_7_212 = _GEN_662;
  wire          _GEN_663 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h14;
  wire          compressDataVec_hitReq_8_20;
  assign compressDataVec_hitReq_8_20 = _GEN_663;
  wire          compressDataVec_hitReq_8_148;
  assign compressDataVec_hitReq_8_148 = _GEN_663;
  wire          compressDataVec_hitReq_8_212;
  assign compressDataVec_hitReq_8_212 = _GEN_663;
  wire          _GEN_664 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h14;
  wire          compressDataVec_hitReq_9_20;
  assign compressDataVec_hitReq_9_20 = _GEN_664;
  wire          compressDataVec_hitReq_9_148;
  assign compressDataVec_hitReq_9_148 = _GEN_664;
  wire          compressDataVec_hitReq_9_212;
  assign compressDataVec_hitReq_9_212 = _GEN_664;
  wire          _GEN_665 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h14;
  wire          compressDataVec_hitReq_10_20;
  assign compressDataVec_hitReq_10_20 = _GEN_665;
  wire          compressDataVec_hitReq_10_148;
  assign compressDataVec_hitReq_10_148 = _GEN_665;
  wire          compressDataVec_hitReq_10_212;
  assign compressDataVec_hitReq_10_212 = _GEN_665;
  wire          _GEN_666 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h14;
  wire          compressDataVec_hitReq_11_20;
  assign compressDataVec_hitReq_11_20 = _GEN_666;
  wire          compressDataVec_hitReq_11_148;
  assign compressDataVec_hitReq_11_148 = _GEN_666;
  wire          compressDataVec_hitReq_11_212;
  assign compressDataVec_hitReq_11_212 = _GEN_666;
  wire          _GEN_667 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h14;
  wire          compressDataVec_hitReq_12_20;
  assign compressDataVec_hitReq_12_20 = _GEN_667;
  wire          compressDataVec_hitReq_12_148;
  assign compressDataVec_hitReq_12_148 = _GEN_667;
  wire          compressDataVec_hitReq_12_212;
  assign compressDataVec_hitReq_12_212 = _GEN_667;
  wire          _GEN_668 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h14;
  wire          compressDataVec_hitReq_13_20;
  assign compressDataVec_hitReq_13_20 = _GEN_668;
  wire          compressDataVec_hitReq_13_148;
  assign compressDataVec_hitReq_13_148 = _GEN_668;
  wire          compressDataVec_hitReq_13_212;
  assign compressDataVec_hitReq_13_212 = _GEN_668;
  wire          _GEN_669 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h14;
  wire          compressDataVec_hitReq_14_20;
  assign compressDataVec_hitReq_14_20 = _GEN_669;
  wire          compressDataVec_hitReq_14_148;
  assign compressDataVec_hitReq_14_148 = _GEN_669;
  wire          compressDataVec_hitReq_14_212;
  assign compressDataVec_hitReq_14_212 = _GEN_669;
  wire          _GEN_670 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h14;
  wire          compressDataVec_hitReq_15_20;
  assign compressDataVec_hitReq_15_20 = _GEN_670;
  wire          compressDataVec_hitReq_15_148;
  assign compressDataVec_hitReq_15_148 = _GEN_670;
  wire          compressDataVec_hitReq_15_212;
  assign compressDataVec_hitReq_15_212 = _GEN_670;
  wire          _GEN_671 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h14;
  wire          compressDataVec_hitReq_16_20;
  assign compressDataVec_hitReq_16_20 = _GEN_671;
  wire          compressDataVec_hitReq_16_148;
  assign compressDataVec_hitReq_16_148 = _GEN_671;
  wire          _GEN_672 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h14;
  wire          compressDataVec_hitReq_17_20;
  assign compressDataVec_hitReq_17_20 = _GEN_672;
  wire          compressDataVec_hitReq_17_148;
  assign compressDataVec_hitReq_17_148 = _GEN_672;
  wire          _GEN_673 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h14;
  wire          compressDataVec_hitReq_18_20;
  assign compressDataVec_hitReq_18_20 = _GEN_673;
  wire          compressDataVec_hitReq_18_148;
  assign compressDataVec_hitReq_18_148 = _GEN_673;
  wire          _GEN_674 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h14;
  wire          compressDataVec_hitReq_19_20;
  assign compressDataVec_hitReq_19_20 = _GEN_674;
  wire          compressDataVec_hitReq_19_148;
  assign compressDataVec_hitReq_19_148 = _GEN_674;
  wire          _GEN_675 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h14;
  wire          compressDataVec_hitReq_20_20;
  assign compressDataVec_hitReq_20_20 = _GEN_675;
  wire          compressDataVec_hitReq_20_148;
  assign compressDataVec_hitReq_20_148 = _GEN_675;
  wire          _GEN_676 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h14;
  wire          compressDataVec_hitReq_21_20;
  assign compressDataVec_hitReq_21_20 = _GEN_676;
  wire          compressDataVec_hitReq_21_148;
  assign compressDataVec_hitReq_21_148 = _GEN_676;
  wire          _GEN_677 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h14;
  wire          compressDataVec_hitReq_22_20;
  assign compressDataVec_hitReq_22_20 = _GEN_677;
  wire          compressDataVec_hitReq_22_148;
  assign compressDataVec_hitReq_22_148 = _GEN_677;
  wire          _GEN_678 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h14;
  wire          compressDataVec_hitReq_23_20;
  assign compressDataVec_hitReq_23_20 = _GEN_678;
  wire          compressDataVec_hitReq_23_148;
  assign compressDataVec_hitReq_23_148 = _GEN_678;
  wire          _GEN_679 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h14;
  wire          compressDataVec_hitReq_24_20;
  assign compressDataVec_hitReq_24_20 = _GEN_679;
  wire          compressDataVec_hitReq_24_148;
  assign compressDataVec_hitReq_24_148 = _GEN_679;
  wire          _GEN_680 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h14;
  wire          compressDataVec_hitReq_25_20;
  assign compressDataVec_hitReq_25_20 = _GEN_680;
  wire          compressDataVec_hitReq_25_148;
  assign compressDataVec_hitReq_25_148 = _GEN_680;
  wire          _GEN_681 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h14;
  wire          compressDataVec_hitReq_26_20;
  assign compressDataVec_hitReq_26_20 = _GEN_681;
  wire          compressDataVec_hitReq_26_148;
  assign compressDataVec_hitReq_26_148 = _GEN_681;
  wire          _GEN_682 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h14;
  wire          compressDataVec_hitReq_27_20;
  assign compressDataVec_hitReq_27_20 = _GEN_682;
  wire          compressDataVec_hitReq_27_148;
  assign compressDataVec_hitReq_27_148 = _GEN_682;
  wire          _GEN_683 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h14;
  wire          compressDataVec_hitReq_28_20;
  assign compressDataVec_hitReq_28_20 = _GEN_683;
  wire          compressDataVec_hitReq_28_148;
  assign compressDataVec_hitReq_28_148 = _GEN_683;
  wire          _GEN_684 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h14;
  wire          compressDataVec_hitReq_29_20;
  assign compressDataVec_hitReq_29_20 = _GEN_684;
  wire          compressDataVec_hitReq_29_148;
  assign compressDataVec_hitReq_29_148 = _GEN_684;
  wire          _GEN_685 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h14;
  wire          compressDataVec_hitReq_30_20;
  assign compressDataVec_hitReq_30_20 = _GEN_685;
  wire          compressDataVec_hitReq_30_148;
  assign compressDataVec_hitReq_30_148 = _GEN_685;
  wire          _GEN_686 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h14;
  wire          compressDataVec_hitReq_31_20;
  assign compressDataVec_hitReq_31_20 = _GEN_686;
  wire          compressDataVec_hitReq_31_148;
  assign compressDataVec_hitReq_31_148 = _GEN_686;
  wire          compressDataVec_hitReq_32_20 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h14;
  wire          compressDataVec_hitReq_33_20 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h14;
  wire          compressDataVec_hitReq_34_20 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h14;
  wire          compressDataVec_hitReq_35_20 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h14;
  wire          compressDataVec_hitReq_36_20 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h14;
  wire          compressDataVec_hitReq_37_20 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h14;
  wire          compressDataVec_hitReq_38_20 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h14;
  wire          compressDataVec_hitReq_39_20 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h14;
  wire          compressDataVec_hitReq_40_20 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h14;
  wire          compressDataVec_hitReq_41_20 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h14;
  wire          compressDataVec_hitReq_42_20 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h14;
  wire          compressDataVec_hitReq_43_20 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h14;
  wire          compressDataVec_hitReq_44_20 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h14;
  wire          compressDataVec_hitReq_45_20 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h14;
  wire          compressDataVec_hitReq_46_20 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h14;
  wire          compressDataVec_hitReq_47_20 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h14;
  wire          compressDataVec_hitReq_48_20 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h14;
  wire          compressDataVec_hitReq_49_20 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h14;
  wire          compressDataVec_hitReq_50_20 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h14;
  wire          compressDataVec_hitReq_51_20 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h14;
  wire          compressDataVec_hitReq_52_20 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h14;
  wire          compressDataVec_hitReq_53_20 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h14;
  wire          compressDataVec_hitReq_54_20 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h14;
  wire          compressDataVec_hitReq_55_20 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h14;
  wire          compressDataVec_hitReq_56_20 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h14;
  wire          compressDataVec_hitReq_57_20 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h14;
  wire          compressDataVec_hitReq_58_20 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h14;
  wire          compressDataVec_hitReq_59_20 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h14;
  wire          compressDataVec_hitReq_60_20 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h14;
  wire          compressDataVec_hitReq_61_20 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h14;
  wire          compressDataVec_hitReq_62_20 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h14;
  wire          compressDataVec_hitReq_63_20 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h14;
  wire [7:0]    compressDataVec_selectReqData_20 =
    (compressDataVec_hitReq_0_20 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_20 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_20 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_20 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_20 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_20 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_20 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_20 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_20 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_20 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_20 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_20 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_20 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_20 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_20 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_20 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_20 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_20 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_20 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_20 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_20 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_20 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_20 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_20 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_20 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_20 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_20 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_20 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_20 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_20 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_20 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_20 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_20 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_20 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_20 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_20 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_20 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_20 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_20 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_20 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_20 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_20 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_20 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_20 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_20 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_20 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_20 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_20 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_20 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_20 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_20 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_20 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_20 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_20 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_20 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_20 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_20 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_20 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_20 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_20 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_20 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_20 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_20 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_20 ? source2Pipe[511:504] : 8'h0);
  wire          _GEN_687 = tailCount > 6'h14;
  wire          compressDataVec_useTail_20;
  assign compressDataVec_useTail_20 = _GEN_687;
  wire          compressDataVec_useTail_84;
  assign compressDataVec_useTail_84 = _GEN_687;
  wire          _GEN_688 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h15;
  wire          compressDataVec_hitReq_0_21;
  assign compressDataVec_hitReq_0_21 = _GEN_688;
  wire          compressDataVec_hitReq_0_149;
  assign compressDataVec_hitReq_0_149 = _GEN_688;
  wire          compressDataVec_hitReq_0_213;
  assign compressDataVec_hitReq_0_213 = _GEN_688;
  wire          _GEN_689 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h15;
  wire          compressDataVec_hitReq_1_21;
  assign compressDataVec_hitReq_1_21 = _GEN_689;
  wire          compressDataVec_hitReq_1_149;
  assign compressDataVec_hitReq_1_149 = _GEN_689;
  wire          compressDataVec_hitReq_1_213;
  assign compressDataVec_hitReq_1_213 = _GEN_689;
  wire          _GEN_690 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h15;
  wire          compressDataVec_hitReq_2_21;
  assign compressDataVec_hitReq_2_21 = _GEN_690;
  wire          compressDataVec_hitReq_2_149;
  assign compressDataVec_hitReq_2_149 = _GEN_690;
  wire          compressDataVec_hitReq_2_213;
  assign compressDataVec_hitReq_2_213 = _GEN_690;
  wire          _GEN_691 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h15;
  wire          compressDataVec_hitReq_3_21;
  assign compressDataVec_hitReq_3_21 = _GEN_691;
  wire          compressDataVec_hitReq_3_149;
  assign compressDataVec_hitReq_3_149 = _GEN_691;
  wire          compressDataVec_hitReq_3_213;
  assign compressDataVec_hitReq_3_213 = _GEN_691;
  wire          _GEN_692 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h15;
  wire          compressDataVec_hitReq_4_21;
  assign compressDataVec_hitReq_4_21 = _GEN_692;
  wire          compressDataVec_hitReq_4_149;
  assign compressDataVec_hitReq_4_149 = _GEN_692;
  wire          compressDataVec_hitReq_4_213;
  assign compressDataVec_hitReq_4_213 = _GEN_692;
  wire          _GEN_693 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h15;
  wire          compressDataVec_hitReq_5_21;
  assign compressDataVec_hitReq_5_21 = _GEN_693;
  wire          compressDataVec_hitReq_5_149;
  assign compressDataVec_hitReq_5_149 = _GEN_693;
  wire          compressDataVec_hitReq_5_213;
  assign compressDataVec_hitReq_5_213 = _GEN_693;
  wire          _GEN_694 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h15;
  wire          compressDataVec_hitReq_6_21;
  assign compressDataVec_hitReq_6_21 = _GEN_694;
  wire          compressDataVec_hitReq_6_149;
  assign compressDataVec_hitReq_6_149 = _GEN_694;
  wire          compressDataVec_hitReq_6_213;
  assign compressDataVec_hitReq_6_213 = _GEN_694;
  wire          _GEN_695 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h15;
  wire          compressDataVec_hitReq_7_21;
  assign compressDataVec_hitReq_7_21 = _GEN_695;
  wire          compressDataVec_hitReq_7_149;
  assign compressDataVec_hitReq_7_149 = _GEN_695;
  wire          compressDataVec_hitReq_7_213;
  assign compressDataVec_hitReq_7_213 = _GEN_695;
  wire          _GEN_696 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h15;
  wire          compressDataVec_hitReq_8_21;
  assign compressDataVec_hitReq_8_21 = _GEN_696;
  wire          compressDataVec_hitReq_8_149;
  assign compressDataVec_hitReq_8_149 = _GEN_696;
  wire          compressDataVec_hitReq_8_213;
  assign compressDataVec_hitReq_8_213 = _GEN_696;
  wire          _GEN_697 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h15;
  wire          compressDataVec_hitReq_9_21;
  assign compressDataVec_hitReq_9_21 = _GEN_697;
  wire          compressDataVec_hitReq_9_149;
  assign compressDataVec_hitReq_9_149 = _GEN_697;
  wire          compressDataVec_hitReq_9_213;
  assign compressDataVec_hitReq_9_213 = _GEN_697;
  wire          _GEN_698 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h15;
  wire          compressDataVec_hitReq_10_21;
  assign compressDataVec_hitReq_10_21 = _GEN_698;
  wire          compressDataVec_hitReq_10_149;
  assign compressDataVec_hitReq_10_149 = _GEN_698;
  wire          compressDataVec_hitReq_10_213;
  assign compressDataVec_hitReq_10_213 = _GEN_698;
  wire          _GEN_699 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h15;
  wire          compressDataVec_hitReq_11_21;
  assign compressDataVec_hitReq_11_21 = _GEN_699;
  wire          compressDataVec_hitReq_11_149;
  assign compressDataVec_hitReq_11_149 = _GEN_699;
  wire          compressDataVec_hitReq_11_213;
  assign compressDataVec_hitReq_11_213 = _GEN_699;
  wire          _GEN_700 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h15;
  wire          compressDataVec_hitReq_12_21;
  assign compressDataVec_hitReq_12_21 = _GEN_700;
  wire          compressDataVec_hitReq_12_149;
  assign compressDataVec_hitReq_12_149 = _GEN_700;
  wire          compressDataVec_hitReq_12_213;
  assign compressDataVec_hitReq_12_213 = _GEN_700;
  wire          _GEN_701 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h15;
  wire          compressDataVec_hitReq_13_21;
  assign compressDataVec_hitReq_13_21 = _GEN_701;
  wire          compressDataVec_hitReq_13_149;
  assign compressDataVec_hitReq_13_149 = _GEN_701;
  wire          compressDataVec_hitReq_13_213;
  assign compressDataVec_hitReq_13_213 = _GEN_701;
  wire          _GEN_702 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h15;
  wire          compressDataVec_hitReq_14_21;
  assign compressDataVec_hitReq_14_21 = _GEN_702;
  wire          compressDataVec_hitReq_14_149;
  assign compressDataVec_hitReq_14_149 = _GEN_702;
  wire          compressDataVec_hitReq_14_213;
  assign compressDataVec_hitReq_14_213 = _GEN_702;
  wire          _GEN_703 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h15;
  wire          compressDataVec_hitReq_15_21;
  assign compressDataVec_hitReq_15_21 = _GEN_703;
  wire          compressDataVec_hitReq_15_149;
  assign compressDataVec_hitReq_15_149 = _GEN_703;
  wire          compressDataVec_hitReq_15_213;
  assign compressDataVec_hitReq_15_213 = _GEN_703;
  wire          _GEN_704 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h15;
  wire          compressDataVec_hitReq_16_21;
  assign compressDataVec_hitReq_16_21 = _GEN_704;
  wire          compressDataVec_hitReq_16_149;
  assign compressDataVec_hitReq_16_149 = _GEN_704;
  wire          _GEN_705 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h15;
  wire          compressDataVec_hitReq_17_21;
  assign compressDataVec_hitReq_17_21 = _GEN_705;
  wire          compressDataVec_hitReq_17_149;
  assign compressDataVec_hitReq_17_149 = _GEN_705;
  wire          _GEN_706 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h15;
  wire          compressDataVec_hitReq_18_21;
  assign compressDataVec_hitReq_18_21 = _GEN_706;
  wire          compressDataVec_hitReq_18_149;
  assign compressDataVec_hitReq_18_149 = _GEN_706;
  wire          _GEN_707 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h15;
  wire          compressDataVec_hitReq_19_21;
  assign compressDataVec_hitReq_19_21 = _GEN_707;
  wire          compressDataVec_hitReq_19_149;
  assign compressDataVec_hitReq_19_149 = _GEN_707;
  wire          _GEN_708 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h15;
  wire          compressDataVec_hitReq_20_21;
  assign compressDataVec_hitReq_20_21 = _GEN_708;
  wire          compressDataVec_hitReq_20_149;
  assign compressDataVec_hitReq_20_149 = _GEN_708;
  wire          _GEN_709 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h15;
  wire          compressDataVec_hitReq_21_21;
  assign compressDataVec_hitReq_21_21 = _GEN_709;
  wire          compressDataVec_hitReq_21_149;
  assign compressDataVec_hitReq_21_149 = _GEN_709;
  wire          _GEN_710 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h15;
  wire          compressDataVec_hitReq_22_21;
  assign compressDataVec_hitReq_22_21 = _GEN_710;
  wire          compressDataVec_hitReq_22_149;
  assign compressDataVec_hitReq_22_149 = _GEN_710;
  wire          _GEN_711 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h15;
  wire          compressDataVec_hitReq_23_21;
  assign compressDataVec_hitReq_23_21 = _GEN_711;
  wire          compressDataVec_hitReq_23_149;
  assign compressDataVec_hitReq_23_149 = _GEN_711;
  wire          _GEN_712 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h15;
  wire          compressDataVec_hitReq_24_21;
  assign compressDataVec_hitReq_24_21 = _GEN_712;
  wire          compressDataVec_hitReq_24_149;
  assign compressDataVec_hitReq_24_149 = _GEN_712;
  wire          _GEN_713 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h15;
  wire          compressDataVec_hitReq_25_21;
  assign compressDataVec_hitReq_25_21 = _GEN_713;
  wire          compressDataVec_hitReq_25_149;
  assign compressDataVec_hitReq_25_149 = _GEN_713;
  wire          _GEN_714 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h15;
  wire          compressDataVec_hitReq_26_21;
  assign compressDataVec_hitReq_26_21 = _GEN_714;
  wire          compressDataVec_hitReq_26_149;
  assign compressDataVec_hitReq_26_149 = _GEN_714;
  wire          _GEN_715 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h15;
  wire          compressDataVec_hitReq_27_21;
  assign compressDataVec_hitReq_27_21 = _GEN_715;
  wire          compressDataVec_hitReq_27_149;
  assign compressDataVec_hitReq_27_149 = _GEN_715;
  wire          _GEN_716 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h15;
  wire          compressDataVec_hitReq_28_21;
  assign compressDataVec_hitReq_28_21 = _GEN_716;
  wire          compressDataVec_hitReq_28_149;
  assign compressDataVec_hitReq_28_149 = _GEN_716;
  wire          _GEN_717 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h15;
  wire          compressDataVec_hitReq_29_21;
  assign compressDataVec_hitReq_29_21 = _GEN_717;
  wire          compressDataVec_hitReq_29_149;
  assign compressDataVec_hitReq_29_149 = _GEN_717;
  wire          _GEN_718 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h15;
  wire          compressDataVec_hitReq_30_21;
  assign compressDataVec_hitReq_30_21 = _GEN_718;
  wire          compressDataVec_hitReq_30_149;
  assign compressDataVec_hitReq_30_149 = _GEN_718;
  wire          _GEN_719 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h15;
  wire          compressDataVec_hitReq_31_21;
  assign compressDataVec_hitReq_31_21 = _GEN_719;
  wire          compressDataVec_hitReq_31_149;
  assign compressDataVec_hitReq_31_149 = _GEN_719;
  wire          compressDataVec_hitReq_32_21 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h15;
  wire          compressDataVec_hitReq_33_21 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h15;
  wire          compressDataVec_hitReq_34_21 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h15;
  wire          compressDataVec_hitReq_35_21 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h15;
  wire          compressDataVec_hitReq_36_21 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h15;
  wire          compressDataVec_hitReq_37_21 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h15;
  wire          compressDataVec_hitReq_38_21 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h15;
  wire          compressDataVec_hitReq_39_21 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h15;
  wire          compressDataVec_hitReq_40_21 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h15;
  wire          compressDataVec_hitReq_41_21 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h15;
  wire          compressDataVec_hitReq_42_21 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h15;
  wire          compressDataVec_hitReq_43_21 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h15;
  wire          compressDataVec_hitReq_44_21 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h15;
  wire          compressDataVec_hitReq_45_21 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h15;
  wire          compressDataVec_hitReq_46_21 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h15;
  wire          compressDataVec_hitReq_47_21 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h15;
  wire          compressDataVec_hitReq_48_21 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h15;
  wire          compressDataVec_hitReq_49_21 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h15;
  wire          compressDataVec_hitReq_50_21 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h15;
  wire          compressDataVec_hitReq_51_21 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h15;
  wire          compressDataVec_hitReq_52_21 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h15;
  wire          compressDataVec_hitReq_53_21 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h15;
  wire          compressDataVec_hitReq_54_21 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h15;
  wire          compressDataVec_hitReq_55_21 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h15;
  wire          compressDataVec_hitReq_56_21 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h15;
  wire          compressDataVec_hitReq_57_21 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h15;
  wire          compressDataVec_hitReq_58_21 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h15;
  wire          compressDataVec_hitReq_59_21 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h15;
  wire          compressDataVec_hitReq_60_21 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h15;
  wire          compressDataVec_hitReq_61_21 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h15;
  wire          compressDataVec_hitReq_62_21 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h15;
  wire          compressDataVec_hitReq_63_21 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h15;
  wire [7:0]    compressDataVec_selectReqData_21 =
    (compressDataVec_hitReq_0_21 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_21 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_21 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_21 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_21 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_21 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_21 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_21 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_21 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_21 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_21 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_21 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_21 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_21 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_21 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_21 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_21 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_21 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_21 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_21 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_21 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_21 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_21 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_21 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_21 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_21 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_21 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_21 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_21 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_21 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_21 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_21 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_21 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_21 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_21 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_21 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_21 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_21 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_21 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_21 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_21 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_21 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_21 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_21 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_21 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_21 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_21 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_21 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_21 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_21 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_21 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_21 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_21 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_21 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_21 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_21 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_21 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_21 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_21 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_21 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_21 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_21 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_21 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_21 ? source2Pipe[511:504] : 8'h0);
  wire          _GEN_720 = tailCount > 6'h15;
  wire          compressDataVec_useTail_21;
  assign compressDataVec_useTail_21 = _GEN_720;
  wire          compressDataVec_useTail_85;
  assign compressDataVec_useTail_85 = _GEN_720;
  wire          _GEN_721 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h16;
  wire          compressDataVec_hitReq_0_22;
  assign compressDataVec_hitReq_0_22 = _GEN_721;
  wire          compressDataVec_hitReq_0_150;
  assign compressDataVec_hitReq_0_150 = _GEN_721;
  wire          compressDataVec_hitReq_0_214;
  assign compressDataVec_hitReq_0_214 = _GEN_721;
  wire          _GEN_722 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h16;
  wire          compressDataVec_hitReq_1_22;
  assign compressDataVec_hitReq_1_22 = _GEN_722;
  wire          compressDataVec_hitReq_1_150;
  assign compressDataVec_hitReq_1_150 = _GEN_722;
  wire          compressDataVec_hitReq_1_214;
  assign compressDataVec_hitReq_1_214 = _GEN_722;
  wire          _GEN_723 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h16;
  wire          compressDataVec_hitReq_2_22;
  assign compressDataVec_hitReq_2_22 = _GEN_723;
  wire          compressDataVec_hitReq_2_150;
  assign compressDataVec_hitReq_2_150 = _GEN_723;
  wire          compressDataVec_hitReq_2_214;
  assign compressDataVec_hitReq_2_214 = _GEN_723;
  wire          _GEN_724 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h16;
  wire          compressDataVec_hitReq_3_22;
  assign compressDataVec_hitReq_3_22 = _GEN_724;
  wire          compressDataVec_hitReq_3_150;
  assign compressDataVec_hitReq_3_150 = _GEN_724;
  wire          compressDataVec_hitReq_3_214;
  assign compressDataVec_hitReq_3_214 = _GEN_724;
  wire          _GEN_725 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h16;
  wire          compressDataVec_hitReq_4_22;
  assign compressDataVec_hitReq_4_22 = _GEN_725;
  wire          compressDataVec_hitReq_4_150;
  assign compressDataVec_hitReq_4_150 = _GEN_725;
  wire          compressDataVec_hitReq_4_214;
  assign compressDataVec_hitReq_4_214 = _GEN_725;
  wire          _GEN_726 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h16;
  wire          compressDataVec_hitReq_5_22;
  assign compressDataVec_hitReq_5_22 = _GEN_726;
  wire          compressDataVec_hitReq_5_150;
  assign compressDataVec_hitReq_5_150 = _GEN_726;
  wire          compressDataVec_hitReq_5_214;
  assign compressDataVec_hitReq_5_214 = _GEN_726;
  wire          _GEN_727 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h16;
  wire          compressDataVec_hitReq_6_22;
  assign compressDataVec_hitReq_6_22 = _GEN_727;
  wire          compressDataVec_hitReq_6_150;
  assign compressDataVec_hitReq_6_150 = _GEN_727;
  wire          compressDataVec_hitReq_6_214;
  assign compressDataVec_hitReq_6_214 = _GEN_727;
  wire          _GEN_728 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h16;
  wire          compressDataVec_hitReq_7_22;
  assign compressDataVec_hitReq_7_22 = _GEN_728;
  wire          compressDataVec_hitReq_7_150;
  assign compressDataVec_hitReq_7_150 = _GEN_728;
  wire          compressDataVec_hitReq_7_214;
  assign compressDataVec_hitReq_7_214 = _GEN_728;
  wire          _GEN_729 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h16;
  wire          compressDataVec_hitReq_8_22;
  assign compressDataVec_hitReq_8_22 = _GEN_729;
  wire          compressDataVec_hitReq_8_150;
  assign compressDataVec_hitReq_8_150 = _GEN_729;
  wire          compressDataVec_hitReq_8_214;
  assign compressDataVec_hitReq_8_214 = _GEN_729;
  wire          _GEN_730 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h16;
  wire          compressDataVec_hitReq_9_22;
  assign compressDataVec_hitReq_9_22 = _GEN_730;
  wire          compressDataVec_hitReq_9_150;
  assign compressDataVec_hitReq_9_150 = _GEN_730;
  wire          compressDataVec_hitReq_9_214;
  assign compressDataVec_hitReq_9_214 = _GEN_730;
  wire          _GEN_731 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h16;
  wire          compressDataVec_hitReq_10_22;
  assign compressDataVec_hitReq_10_22 = _GEN_731;
  wire          compressDataVec_hitReq_10_150;
  assign compressDataVec_hitReq_10_150 = _GEN_731;
  wire          compressDataVec_hitReq_10_214;
  assign compressDataVec_hitReq_10_214 = _GEN_731;
  wire          _GEN_732 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h16;
  wire          compressDataVec_hitReq_11_22;
  assign compressDataVec_hitReq_11_22 = _GEN_732;
  wire          compressDataVec_hitReq_11_150;
  assign compressDataVec_hitReq_11_150 = _GEN_732;
  wire          compressDataVec_hitReq_11_214;
  assign compressDataVec_hitReq_11_214 = _GEN_732;
  wire          _GEN_733 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h16;
  wire          compressDataVec_hitReq_12_22;
  assign compressDataVec_hitReq_12_22 = _GEN_733;
  wire          compressDataVec_hitReq_12_150;
  assign compressDataVec_hitReq_12_150 = _GEN_733;
  wire          compressDataVec_hitReq_12_214;
  assign compressDataVec_hitReq_12_214 = _GEN_733;
  wire          _GEN_734 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h16;
  wire          compressDataVec_hitReq_13_22;
  assign compressDataVec_hitReq_13_22 = _GEN_734;
  wire          compressDataVec_hitReq_13_150;
  assign compressDataVec_hitReq_13_150 = _GEN_734;
  wire          compressDataVec_hitReq_13_214;
  assign compressDataVec_hitReq_13_214 = _GEN_734;
  wire          _GEN_735 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h16;
  wire          compressDataVec_hitReq_14_22;
  assign compressDataVec_hitReq_14_22 = _GEN_735;
  wire          compressDataVec_hitReq_14_150;
  assign compressDataVec_hitReq_14_150 = _GEN_735;
  wire          compressDataVec_hitReq_14_214;
  assign compressDataVec_hitReq_14_214 = _GEN_735;
  wire          _GEN_736 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h16;
  wire          compressDataVec_hitReq_15_22;
  assign compressDataVec_hitReq_15_22 = _GEN_736;
  wire          compressDataVec_hitReq_15_150;
  assign compressDataVec_hitReq_15_150 = _GEN_736;
  wire          compressDataVec_hitReq_15_214;
  assign compressDataVec_hitReq_15_214 = _GEN_736;
  wire          _GEN_737 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h16;
  wire          compressDataVec_hitReq_16_22;
  assign compressDataVec_hitReq_16_22 = _GEN_737;
  wire          compressDataVec_hitReq_16_150;
  assign compressDataVec_hitReq_16_150 = _GEN_737;
  wire          _GEN_738 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h16;
  wire          compressDataVec_hitReq_17_22;
  assign compressDataVec_hitReq_17_22 = _GEN_738;
  wire          compressDataVec_hitReq_17_150;
  assign compressDataVec_hitReq_17_150 = _GEN_738;
  wire          _GEN_739 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h16;
  wire          compressDataVec_hitReq_18_22;
  assign compressDataVec_hitReq_18_22 = _GEN_739;
  wire          compressDataVec_hitReq_18_150;
  assign compressDataVec_hitReq_18_150 = _GEN_739;
  wire          _GEN_740 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h16;
  wire          compressDataVec_hitReq_19_22;
  assign compressDataVec_hitReq_19_22 = _GEN_740;
  wire          compressDataVec_hitReq_19_150;
  assign compressDataVec_hitReq_19_150 = _GEN_740;
  wire          _GEN_741 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h16;
  wire          compressDataVec_hitReq_20_22;
  assign compressDataVec_hitReq_20_22 = _GEN_741;
  wire          compressDataVec_hitReq_20_150;
  assign compressDataVec_hitReq_20_150 = _GEN_741;
  wire          _GEN_742 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h16;
  wire          compressDataVec_hitReq_21_22;
  assign compressDataVec_hitReq_21_22 = _GEN_742;
  wire          compressDataVec_hitReq_21_150;
  assign compressDataVec_hitReq_21_150 = _GEN_742;
  wire          _GEN_743 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h16;
  wire          compressDataVec_hitReq_22_22;
  assign compressDataVec_hitReq_22_22 = _GEN_743;
  wire          compressDataVec_hitReq_22_150;
  assign compressDataVec_hitReq_22_150 = _GEN_743;
  wire          _GEN_744 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h16;
  wire          compressDataVec_hitReq_23_22;
  assign compressDataVec_hitReq_23_22 = _GEN_744;
  wire          compressDataVec_hitReq_23_150;
  assign compressDataVec_hitReq_23_150 = _GEN_744;
  wire          _GEN_745 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h16;
  wire          compressDataVec_hitReq_24_22;
  assign compressDataVec_hitReq_24_22 = _GEN_745;
  wire          compressDataVec_hitReq_24_150;
  assign compressDataVec_hitReq_24_150 = _GEN_745;
  wire          _GEN_746 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h16;
  wire          compressDataVec_hitReq_25_22;
  assign compressDataVec_hitReq_25_22 = _GEN_746;
  wire          compressDataVec_hitReq_25_150;
  assign compressDataVec_hitReq_25_150 = _GEN_746;
  wire          _GEN_747 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h16;
  wire          compressDataVec_hitReq_26_22;
  assign compressDataVec_hitReq_26_22 = _GEN_747;
  wire          compressDataVec_hitReq_26_150;
  assign compressDataVec_hitReq_26_150 = _GEN_747;
  wire          _GEN_748 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h16;
  wire          compressDataVec_hitReq_27_22;
  assign compressDataVec_hitReq_27_22 = _GEN_748;
  wire          compressDataVec_hitReq_27_150;
  assign compressDataVec_hitReq_27_150 = _GEN_748;
  wire          _GEN_749 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h16;
  wire          compressDataVec_hitReq_28_22;
  assign compressDataVec_hitReq_28_22 = _GEN_749;
  wire          compressDataVec_hitReq_28_150;
  assign compressDataVec_hitReq_28_150 = _GEN_749;
  wire          _GEN_750 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h16;
  wire          compressDataVec_hitReq_29_22;
  assign compressDataVec_hitReq_29_22 = _GEN_750;
  wire          compressDataVec_hitReq_29_150;
  assign compressDataVec_hitReq_29_150 = _GEN_750;
  wire          _GEN_751 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h16;
  wire          compressDataVec_hitReq_30_22;
  assign compressDataVec_hitReq_30_22 = _GEN_751;
  wire          compressDataVec_hitReq_30_150;
  assign compressDataVec_hitReq_30_150 = _GEN_751;
  wire          _GEN_752 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h16;
  wire          compressDataVec_hitReq_31_22;
  assign compressDataVec_hitReq_31_22 = _GEN_752;
  wire          compressDataVec_hitReq_31_150;
  assign compressDataVec_hitReq_31_150 = _GEN_752;
  wire          compressDataVec_hitReq_32_22 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h16;
  wire          compressDataVec_hitReq_33_22 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h16;
  wire          compressDataVec_hitReq_34_22 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h16;
  wire          compressDataVec_hitReq_35_22 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h16;
  wire          compressDataVec_hitReq_36_22 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h16;
  wire          compressDataVec_hitReq_37_22 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h16;
  wire          compressDataVec_hitReq_38_22 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h16;
  wire          compressDataVec_hitReq_39_22 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h16;
  wire          compressDataVec_hitReq_40_22 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h16;
  wire          compressDataVec_hitReq_41_22 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h16;
  wire          compressDataVec_hitReq_42_22 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h16;
  wire          compressDataVec_hitReq_43_22 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h16;
  wire          compressDataVec_hitReq_44_22 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h16;
  wire          compressDataVec_hitReq_45_22 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h16;
  wire          compressDataVec_hitReq_46_22 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h16;
  wire          compressDataVec_hitReq_47_22 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h16;
  wire          compressDataVec_hitReq_48_22 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h16;
  wire          compressDataVec_hitReq_49_22 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h16;
  wire          compressDataVec_hitReq_50_22 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h16;
  wire          compressDataVec_hitReq_51_22 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h16;
  wire          compressDataVec_hitReq_52_22 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h16;
  wire          compressDataVec_hitReq_53_22 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h16;
  wire          compressDataVec_hitReq_54_22 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h16;
  wire          compressDataVec_hitReq_55_22 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h16;
  wire          compressDataVec_hitReq_56_22 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h16;
  wire          compressDataVec_hitReq_57_22 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h16;
  wire          compressDataVec_hitReq_58_22 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h16;
  wire          compressDataVec_hitReq_59_22 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h16;
  wire          compressDataVec_hitReq_60_22 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h16;
  wire          compressDataVec_hitReq_61_22 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h16;
  wire          compressDataVec_hitReq_62_22 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h16;
  wire          compressDataVec_hitReq_63_22 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h16;
  wire [7:0]    compressDataVec_selectReqData_22 =
    (compressDataVec_hitReq_0_22 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_22 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_22 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_22 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_22 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_22 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_22 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_22 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_22 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_22 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_22 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_22 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_22 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_22 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_22 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_22 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_22 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_22 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_22 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_22 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_22 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_22 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_22 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_22 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_22 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_22 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_22 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_22 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_22 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_22 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_22 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_22 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_22 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_22 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_22 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_22 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_22 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_22 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_22 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_22 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_22 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_22 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_22 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_22 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_22 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_22 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_22 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_22 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_22 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_22 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_22 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_22 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_22 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_22 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_22 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_22 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_22 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_22 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_22 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_22 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_22 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_22 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_22 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_22 ? source2Pipe[511:504] : 8'h0);
  wire          _GEN_753 = tailCount > 6'h16;
  wire          compressDataVec_useTail_22;
  assign compressDataVec_useTail_22 = _GEN_753;
  wire          compressDataVec_useTail_86;
  assign compressDataVec_useTail_86 = _GEN_753;
  wire          _GEN_754 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h17;
  wire          compressDataVec_hitReq_0_23;
  assign compressDataVec_hitReq_0_23 = _GEN_754;
  wire          compressDataVec_hitReq_0_151;
  assign compressDataVec_hitReq_0_151 = _GEN_754;
  wire          compressDataVec_hitReq_0_215;
  assign compressDataVec_hitReq_0_215 = _GEN_754;
  wire          _GEN_755 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h17;
  wire          compressDataVec_hitReq_1_23;
  assign compressDataVec_hitReq_1_23 = _GEN_755;
  wire          compressDataVec_hitReq_1_151;
  assign compressDataVec_hitReq_1_151 = _GEN_755;
  wire          compressDataVec_hitReq_1_215;
  assign compressDataVec_hitReq_1_215 = _GEN_755;
  wire          _GEN_756 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h17;
  wire          compressDataVec_hitReq_2_23;
  assign compressDataVec_hitReq_2_23 = _GEN_756;
  wire          compressDataVec_hitReq_2_151;
  assign compressDataVec_hitReq_2_151 = _GEN_756;
  wire          compressDataVec_hitReq_2_215;
  assign compressDataVec_hitReq_2_215 = _GEN_756;
  wire          _GEN_757 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h17;
  wire          compressDataVec_hitReq_3_23;
  assign compressDataVec_hitReq_3_23 = _GEN_757;
  wire          compressDataVec_hitReq_3_151;
  assign compressDataVec_hitReq_3_151 = _GEN_757;
  wire          compressDataVec_hitReq_3_215;
  assign compressDataVec_hitReq_3_215 = _GEN_757;
  wire          _GEN_758 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h17;
  wire          compressDataVec_hitReq_4_23;
  assign compressDataVec_hitReq_4_23 = _GEN_758;
  wire          compressDataVec_hitReq_4_151;
  assign compressDataVec_hitReq_4_151 = _GEN_758;
  wire          compressDataVec_hitReq_4_215;
  assign compressDataVec_hitReq_4_215 = _GEN_758;
  wire          _GEN_759 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h17;
  wire          compressDataVec_hitReq_5_23;
  assign compressDataVec_hitReq_5_23 = _GEN_759;
  wire          compressDataVec_hitReq_5_151;
  assign compressDataVec_hitReq_5_151 = _GEN_759;
  wire          compressDataVec_hitReq_5_215;
  assign compressDataVec_hitReq_5_215 = _GEN_759;
  wire          _GEN_760 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h17;
  wire          compressDataVec_hitReq_6_23;
  assign compressDataVec_hitReq_6_23 = _GEN_760;
  wire          compressDataVec_hitReq_6_151;
  assign compressDataVec_hitReq_6_151 = _GEN_760;
  wire          compressDataVec_hitReq_6_215;
  assign compressDataVec_hitReq_6_215 = _GEN_760;
  wire          _GEN_761 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h17;
  wire          compressDataVec_hitReq_7_23;
  assign compressDataVec_hitReq_7_23 = _GEN_761;
  wire          compressDataVec_hitReq_7_151;
  assign compressDataVec_hitReq_7_151 = _GEN_761;
  wire          compressDataVec_hitReq_7_215;
  assign compressDataVec_hitReq_7_215 = _GEN_761;
  wire          _GEN_762 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h17;
  wire          compressDataVec_hitReq_8_23;
  assign compressDataVec_hitReq_8_23 = _GEN_762;
  wire          compressDataVec_hitReq_8_151;
  assign compressDataVec_hitReq_8_151 = _GEN_762;
  wire          compressDataVec_hitReq_8_215;
  assign compressDataVec_hitReq_8_215 = _GEN_762;
  wire          _GEN_763 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h17;
  wire          compressDataVec_hitReq_9_23;
  assign compressDataVec_hitReq_9_23 = _GEN_763;
  wire          compressDataVec_hitReq_9_151;
  assign compressDataVec_hitReq_9_151 = _GEN_763;
  wire          compressDataVec_hitReq_9_215;
  assign compressDataVec_hitReq_9_215 = _GEN_763;
  wire          _GEN_764 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h17;
  wire          compressDataVec_hitReq_10_23;
  assign compressDataVec_hitReq_10_23 = _GEN_764;
  wire          compressDataVec_hitReq_10_151;
  assign compressDataVec_hitReq_10_151 = _GEN_764;
  wire          compressDataVec_hitReq_10_215;
  assign compressDataVec_hitReq_10_215 = _GEN_764;
  wire          _GEN_765 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h17;
  wire          compressDataVec_hitReq_11_23;
  assign compressDataVec_hitReq_11_23 = _GEN_765;
  wire          compressDataVec_hitReq_11_151;
  assign compressDataVec_hitReq_11_151 = _GEN_765;
  wire          compressDataVec_hitReq_11_215;
  assign compressDataVec_hitReq_11_215 = _GEN_765;
  wire          _GEN_766 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h17;
  wire          compressDataVec_hitReq_12_23;
  assign compressDataVec_hitReq_12_23 = _GEN_766;
  wire          compressDataVec_hitReq_12_151;
  assign compressDataVec_hitReq_12_151 = _GEN_766;
  wire          compressDataVec_hitReq_12_215;
  assign compressDataVec_hitReq_12_215 = _GEN_766;
  wire          _GEN_767 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h17;
  wire          compressDataVec_hitReq_13_23;
  assign compressDataVec_hitReq_13_23 = _GEN_767;
  wire          compressDataVec_hitReq_13_151;
  assign compressDataVec_hitReq_13_151 = _GEN_767;
  wire          compressDataVec_hitReq_13_215;
  assign compressDataVec_hitReq_13_215 = _GEN_767;
  wire          _GEN_768 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h17;
  wire          compressDataVec_hitReq_14_23;
  assign compressDataVec_hitReq_14_23 = _GEN_768;
  wire          compressDataVec_hitReq_14_151;
  assign compressDataVec_hitReq_14_151 = _GEN_768;
  wire          compressDataVec_hitReq_14_215;
  assign compressDataVec_hitReq_14_215 = _GEN_768;
  wire          _GEN_769 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h17;
  wire          compressDataVec_hitReq_15_23;
  assign compressDataVec_hitReq_15_23 = _GEN_769;
  wire          compressDataVec_hitReq_15_151;
  assign compressDataVec_hitReq_15_151 = _GEN_769;
  wire          compressDataVec_hitReq_15_215;
  assign compressDataVec_hitReq_15_215 = _GEN_769;
  wire          _GEN_770 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h17;
  wire          compressDataVec_hitReq_16_23;
  assign compressDataVec_hitReq_16_23 = _GEN_770;
  wire          compressDataVec_hitReq_16_151;
  assign compressDataVec_hitReq_16_151 = _GEN_770;
  wire          _GEN_771 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h17;
  wire          compressDataVec_hitReq_17_23;
  assign compressDataVec_hitReq_17_23 = _GEN_771;
  wire          compressDataVec_hitReq_17_151;
  assign compressDataVec_hitReq_17_151 = _GEN_771;
  wire          _GEN_772 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h17;
  wire          compressDataVec_hitReq_18_23;
  assign compressDataVec_hitReq_18_23 = _GEN_772;
  wire          compressDataVec_hitReq_18_151;
  assign compressDataVec_hitReq_18_151 = _GEN_772;
  wire          _GEN_773 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h17;
  wire          compressDataVec_hitReq_19_23;
  assign compressDataVec_hitReq_19_23 = _GEN_773;
  wire          compressDataVec_hitReq_19_151;
  assign compressDataVec_hitReq_19_151 = _GEN_773;
  wire          _GEN_774 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h17;
  wire          compressDataVec_hitReq_20_23;
  assign compressDataVec_hitReq_20_23 = _GEN_774;
  wire          compressDataVec_hitReq_20_151;
  assign compressDataVec_hitReq_20_151 = _GEN_774;
  wire          _GEN_775 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h17;
  wire          compressDataVec_hitReq_21_23;
  assign compressDataVec_hitReq_21_23 = _GEN_775;
  wire          compressDataVec_hitReq_21_151;
  assign compressDataVec_hitReq_21_151 = _GEN_775;
  wire          _GEN_776 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h17;
  wire          compressDataVec_hitReq_22_23;
  assign compressDataVec_hitReq_22_23 = _GEN_776;
  wire          compressDataVec_hitReq_22_151;
  assign compressDataVec_hitReq_22_151 = _GEN_776;
  wire          _GEN_777 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h17;
  wire          compressDataVec_hitReq_23_23;
  assign compressDataVec_hitReq_23_23 = _GEN_777;
  wire          compressDataVec_hitReq_23_151;
  assign compressDataVec_hitReq_23_151 = _GEN_777;
  wire          _GEN_778 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h17;
  wire          compressDataVec_hitReq_24_23;
  assign compressDataVec_hitReq_24_23 = _GEN_778;
  wire          compressDataVec_hitReq_24_151;
  assign compressDataVec_hitReq_24_151 = _GEN_778;
  wire          _GEN_779 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h17;
  wire          compressDataVec_hitReq_25_23;
  assign compressDataVec_hitReq_25_23 = _GEN_779;
  wire          compressDataVec_hitReq_25_151;
  assign compressDataVec_hitReq_25_151 = _GEN_779;
  wire          _GEN_780 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h17;
  wire          compressDataVec_hitReq_26_23;
  assign compressDataVec_hitReq_26_23 = _GEN_780;
  wire          compressDataVec_hitReq_26_151;
  assign compressDataVec_hitReq_26_151 = _GEN_780;
  wire          _GEN_781 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h17;
  wire          compressDataVec_hitReq_27_23;
  assign compressDataVec_hitReq_27_23 = _GEN_781;
  wire          compressDataVec_hitReq_27_151;
  assign compressDataVec_hitReq_27_151 = _GEN_781;
  wire          _GEN_782 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h17;
  wire          compressDataVec_hitReq_28_23;
  assign compressDataVec_hitReq_28_23 = _GEN_782;
  wire          compressDataVec_hitReq_28_151;
  assign compressDataVec_hitReq_28_151 = _GEN_782;
  wire          _GEN_783 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h17;
  wire          compressDataVec_hitReq_29_23;
  assign compressDataVec_hitReq_29_23 = _GEN_783;
  wire          compressDataVec_hitReq_29_151;
  assign compressDataVec_hitReq_29_151 = _GEN_783;
  wire          _GEN_784 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h17;
  wire          compressDataVec_hitReq_30_23;
  assign compressDataVec_hitReq_30_23 = _GEN_784;
  wire          compressDataVec_hitReq_30_151;
  assign compressDataVec_hitReq_30_151 = _GEN_784;
  wire          _GEN_785 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h17;
  wire          compressDataVec_hitReq_31_23;
  assign compressDataVec_hitReq_31_23 = _GEN_785;
  wire          compressDataVec_hitReq_31_151;
  assign compressDataVec_hitReq_31_151 = _GEN_785;
  wire          compressDataVec_hitReq_32_23 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h17;
  wire          compressDataVec_hitReq_33_23 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h17;
  wire          compressDataVec_hitReq_34_23 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h17;
  wire          compressDataVec_hitReq_35_23 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h17;
  wire          compressDataVec_hitReq_36_23 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h17;
  wire          compressDataVec_hitReq_37_23 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h17;
  wire          compressDataVec_hitReq_38_23 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h17;
  wire          compressDataVec_hitReq_39_23 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h17;
  wire          compressDataVec_hitReq_40_23 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h17;
  wire          compressDataVec_hitReq_41_23 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h17;
  wire          compressDataVec_hitReq_42_23 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h17;
  wire          compressDataVec_hitReq_43_23 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h17;
  wire          compressDataVec_hitReq_44_23 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h17;
  wire          compressDataVec_hitReq_45_23 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h17;
  wire          compressDataVec_hitReq_46_23 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h17;
  wire          compressDataVec_hitReq_47_23 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h17;
  wire          compressDataVec_hitReq_48_23 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h17;
  wire          compressDataVec_hitReq_49_23 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h17;
  wire          compressDataVec_hitReq_50_23 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h17;
  wire          compressDataVec_hitReq_51_23 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h17;
  wire          compressDataVec_hitReq_52_23 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h17;
  wire          compressDataVec_hitReq_53_23 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h17;
  wire          compressDataVec_hitReq_54_23 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h17;
  wire          compressDataVec_hitReq_55_23 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h17;
  wire          compressDataVec_hitReq_56_23 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h17;
  wire          compressDataVec_hitReq_57_23 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h17;
  wire          compressDataVec_hitReq_58_23 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h17;
  wire          compressDataVec_hitReq_59_23 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h17;
  wire          compressDataVec_hitReq_60_23 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h17;
  wire          compressDataVec_hitReq_61_23 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h17;
  wire          compressDataVec_hitReq_62_23 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h17;
  wire          compressDataVec_hitReq_63_23 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h17;
  wire [7:0]    compressDataVec_selectReqData_23 =
    (compressDataVec_hitReq_0_23 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_23 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_23 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_23 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_23 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_23 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_23 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_23 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_23 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_23 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_23 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_23 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_23 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_23 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_23 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_23 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_23 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_23 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_23 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_23 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_23 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_23 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_23 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_23 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_23 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_23 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_23 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_23 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_23 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_23 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_23 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_23 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_23 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_23 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_23 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_23 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_23 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_23 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_23 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_23 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_23 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_23 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_23 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_23 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_23 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_23 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_23 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_23 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_23 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_23 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_23 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_23 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_23 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_23 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_23 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_23 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_23 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_23 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_23 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_23 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_23 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_23 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_23 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_23 ? source2Pipe[511:504] : 8'h0);
  wire          _GEN_786 = tailCount > 6'h17;
  wire          compressDataVec_useTail_23;
  assign compressDataVec_useTail_23 = _GEN_786;
  wire          compressDataVec_useTail_87;
  assign compressDataVec_useTail_87 = _GEN_786;
  wire          _GEN_787 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h18;
  wire          compressDataVec_hitReq_0_24;
  assign compressDataVec_hitReq_0_24 = _GEN_787;
  wire          compressDataVec_hitReq_0_152;
  assign compressDataVec_hitReq_0_152 = _GEN_787;
  wire          compressDataVec_hitReq_0_216;
  assign compressDataVec_hitReq_0_216 = _GEN_787;
  wire          _GEN_788 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h18;
  wire          compressDataVec_hitReq_1_24;
  assign compressDataVec_hitReq_1_24 = _GEN_788;
  wire          compressDataVec_hitReq_1_152;
  assign compressDataVec_hitReq_1_152 = _GEN_788;
  wire          compressDataVec_hitReq_1_216;
  assign compressDataVec_hitReq_1_216 = _GEN_788;
  wire          _GEN_789 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h18;
  wire          compressDataVec_hitReq_2_24;
  assign compressDataVec_hitReq_2_24 = _GEN_789;
  wire          compressDataVec_hitReq_2_152;
  assign compressDataVec_hitReq_2_152 = _GEN_789;
  wire          compressDataVec_hitReq_2_216;
  assign compressDataVec_hitReq_2_216 = _GEN_789;
  wire          _GEN_790 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h18;
  wire          compressDataVec_hitReq_3_24;
  assign compressDataVec_hitReq_3_24 = _GEN_790;
  wire          compressDataVec_hitReq_3_152;
  assign compressDataVec_hitReq_3_152 = _GEN_790;
  wire          compressDataVec_hitReq_3_216;
  assign compressDataVec_hitReq_3_216 = _GEN_790;
  wire          _GEN_791 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h18;
  wire          compressDataVec_hitReq_4_24;
  assign compressDataVec_hitReq_4_24 = _GEN_791;
  wire          compressDataVec_hitReq_4_152;
  assign compressDataVec_hitReq_4_152 = _GEN_791;
  wire          compressDataVec_hitReq_4_216;
  assign compressDataVec_hitReq_4_216 = _GEN_791;
  wire          _GEN_792 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h18;
  wire          compressDataVec_hitReq_5_24;
  assign compressDataVec_hitReq_5_24 = _GEN_792;
  wire          compressDataVec_hitReq_5_152;
  assign compressDataVec_hitReq_5_152 = _GEN_792;
  wire          compressDataVec_hitReq_5_216;
  assign compressDataVec_hitReq_5_216 = _GEN_792;
  wire          _GEN_793 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h18;
  wire          compressDataVec_hitReq_6_24;
  assign compressDataVec_hitReq_6_24 = _GEN_793;
  wire          compressDataVec_hitReq_6_152;
  assign compressDataVec_hitReq_6_152 = _GEN_793;
  wire          compressDataVec_hitReq_6_216;
  assign compressDataVec_hitReq_6_216 = _GEN_793;
  wire          _GEN_794 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h18;
  wire          compressDataVec_hitReq_7_24;
  assign compressDataVec_hitReq_7_24 = _GEN_794;
  wire          compressDataVec_hitReq_7_152;
  assign compressDataVec_hitReq_7_152 = _GEN_794;
  wire          compressDataVec_hitReq_7_216;
  assign compressDataVec_hitReq_7_216 = _GEN_794;
  wire          _GEN_795 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h18;
  wire          compressDataVec_hitReq_8_24;
  assign compressDataVec_hitReq_8_24 = _GEN_795;
  wire          compressDataVec_hitReq_8_152;
  assign compressDataVec_hitReq_8_152 = _GEN_795;
  wire          compressDataVec_hitReq_8_216;
  assign compressDataVec_hitReq_8_216 = _GEN_795;
  wire          _GEN_796 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h18;
  wire          compressDataVec_hitReq_9_24;
  assign compressDataVec_hitReq_9_24 = _GEN_796;
  wire          compressDataVec_hitReq_9_152;
  assign compressDataVec_hitReq_9_152 = _GEN_796;
  wire          compressDataVec_hitReq_9_216;
  assign compressDataVec_hitReq_9_216 = _GEN_796;
  wire          _GEN_797 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h18;
  wire          compressDataVec_hitReq_10_24;
  assign compressDataVec_hitReq_10_24 = _GEN_797;
  wire          compressDataVec_hitReq_10_152;
  assign compressDataVec_hitReq_10_152 = _GEN_797;
  wire          compressDataVec_hitReq_10_216;
  assign compressDataVec_hitReq_10_216 = _GEN_797;
  wire          _GEN_798 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h18;
  wire          compressDataVec_hitReq_11_24;
  assign compressDataVec_hitReq_11_24 = _GEN_798;
  wire          compressDataVec_hitReq_11_152;
  assign compressDataVec_hitReq_11_152 = _GEN_798;
  wire          compressDataVec_hitReq_11_216;
  assign compressDataVec_hitReq_11_216 = _GEN_798;
  wire          _GEN_799 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h18;
  wire          compressDataVec_hitReq_12_24;
  assign compressDataVec_hitReq_12_24 = _GEN_799;
  wire          compressDataVec_hitReq_12_152;
  assign compressDataVec_hitReq_12_152 = _GEN_799;
  wire          compressDataVec_hitReq_12_216;
  assign compressDataVec_hitReq_12_216 = _GEN_799;
  wire          _GEN_800 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h18;
  wire          compressDataVec_hitReq_13_24;
  assign compressDataVec_hitReq_13_24 = _GEN_800;
  wire          compressDataVec_hitReq_13_152;
  assign compressDataVec_hitReq_13_152 = _GEN_800;
  wire          compressDataVec_hitReq_13_216;
  assign compressDataVec_hitReq_13_216 = _GEN_800;
  wire          _GEN_801 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h18;
  wire          compressDataVec_hitReq_14_24;
  assign compressDataVec_hitReq_14_24 = _GEN_801;
  wire          compressDataVec_hitReq_14_152;
  assign compressDataVec_hitReq_14_152 = _GEN_801;
  wire          compressDataVec_hitReq_14_216;
  assign compressDataVec_hitReq_14_216 = _GEN_801;
  wire          _GEN_802 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h18;
  wire          compressDataVec_hitReq_15_24;
  assign compressDataVec_hitReq_15_24 = _GEN_802;
  wire          compressDataVec_hitReq_15_152;
  assign compressDataVec_hitReq_15_152 = _GEN_802;
  wire          compressDataVec_hitReq_15_216;
  assign compressDataVec_hitReq_15_216 = _GEN_802;
  wire          _GEN_803 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h18;
  wire          compressDataVec_hitReq_16_24;
  assign compressDataVec_hitReq_16_24 = _GEN_803;
  wire          compressDataVec_hitReq_16_152;
  assign compressDataVec_hitReq_16_152 = _GEN_803;
  wire          _GEN_804 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h18;
  wire          compressDataVec_hitReq_17_24;
  assign compressDataVec_hitReq_17_24 = _GEN_804;
  wire          compressDataVec_hitReq_17_152;
  assign compressDataVec_hitReq_17_152 = _GEN_804;
  wire          _GEN_805 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h18;
  wire          compressDataVec_hitReq_18_24;
  assign compressDataVec_hitReq_18_24 = _GEN_805;
  wire          compressDataVec_hitReq_18_152;
  assign compressDataVec_hitReq_18_152 = _GEN_805;
  wire          _GEN_806 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h18;
  wire          compressDataVec_hitReq_19_24;
  assign compressDataVec_hitReq_19_24 = _GEN_806;
  wire          compressDataVec_hitReq_19_152;
  assign compressDataVec_hitReq_19_152 = _GEN_806;
  wire          _GEN_807 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h18;
  wire          compressDataVec_hitReq_20_24;
  assign compressDataVec_hitReq_20_24 = _GEN_807;
  wire          compressDataVec_hitReq_20_152;
  assign compressDataVec_hitReq_20_152 = _GEN_807;
  wire          _GEN_808 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h18;
  wire          compressDataVec_hitReq_21_24;
  assign compressDataVec_hitReq_21_24 = _GEN_808;
  wire          compressDataVec_hitReq_21_152;
  assign compressDataVec_hitReq_21_152 = _GEN_808;
  wire          _GEN_809 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h18;
  wire          compressDataVec_hitReq_22_24;
  assign compressDataVec_hitReq_22_24 = _GEN_809;
  wire          compressDataVec_hitReq_22_152;
  assign compressDataVec_hitReq_22_152 = _GEN_809;
  wire          _GEN_810 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h18;
  wire          compressDataVec_hitReq_23_24;
  assign compressDataVec_hitReq_23_24 = _GEN_810;
  wire          compressDataVec_hitReq_23_152;
  assign compressDataVec_hitReq_23_152 = _GEN_810;
  wire          _GEN_811 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h18;
  wire          compressDataVec_hitReq_24_24;
  assign compressDataVec_hitReq_24_24 = _GEN_811;
  wire          compressDataVec_hitReq_24_152;
  assign compressDataVec_hitReq_24_152 = _GEN_811;
  wire          _GEN_812 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h18;
  wire          compressDataVec_hitReq_25_24;
  assign compressDataVec_hitReq_25_24 = _GEN_812;
  wire          compressDataVec_hitReq_25_152;
  assign compressDataVec_hitReq_25_152 = _GEN_812;
  wire          _GEN_813 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h18;
  wire          compressDataVec_hitReq_26_24;
  assign compressDataVec_hitReq_26_24 = _GEN_813;
  wire          compressDataVec_hitReq_26_152;
  assign compressDataVec_hitReq_26_152 = _GEN_813;
  wire          _GEN_814 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h18;
  wire          compressDataVec_hitReq_27_24;
  assign compressDataVec_hitReq_27_24 = _GEN_814;
  wire          compressDataVec_hitReq_27_152;
  assign compressDataVec_hitReq_27_152 = _GEN_814;
  wire          _GEN_815 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h18;
  wire          compressDataVec_hitReq_28_24;
  assign compressDataVec_hitReq_28_24 = _GEN_815;
  wire          compressDataVec_hitReq_28_152;
  assign compressDataVec_hitReq_28_152 = _GEN_815;
  wire          _GEN_816 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h18;
  wire          compressDataVec_hitReq_29_24;
  assign compressDataVec_hitReq_29_24 = _GEN_816;
  wire          compressDataVec_hitReq_29_152;
  assign compressDataVec_hitReq_29_152 = _GEN_816;
  wire          _GEN_817 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h18;
  wire          compressDataVec_hitReq_30_24;
  assign compressDataVec_hitReq_30_24 = _GEN_817;
  wire          compressDataVec_hitReq_30_152;
  assign compressDataVec_hitReq_30_152 = _GEN_817;
  wire          _GEN_818 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h18;
  wire          compressDataVec_hitReq_31_24;
  assign compressDataVec_hitReq_31_24 = _GEN_818;
  wire          compressDataVec_hitReq_31_152;
  assign compressDataVec_hitReq_31_152 = _GEN_818;
  wire          compressDataVec_hitReq_32_24 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h18;
  wire          compressDataVec_hitReq_33_24 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h18;
  wire          compressDataVec_hitReq_34_24 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h18;
  wire          compressDataVec_hitReq_35_24 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h18;
  wire          compressDataVec_hitReq_36_24 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h18;
  wire          compressDataVec_hitReq_37_24 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h18;
  wire          compressDataVec_hitReq_38_24 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h18;
  wire          compressDataVec_hitReq_39_24 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h18;
  wire          compressDataVec_hitReq_40_24 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h18;
  wire          compressDataVec_hitReq_41_24 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h18;
  wire          compressDataVec_hitReq_42_24 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h18;
  wire          compressDataVec_hitReq_43_24 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h18;
  wire          compressDataVec_hitReq_44_24 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h18;
  wire          compressDataVec_hitReq_45_24 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h18;
  wire          compressDataVec_hitReq_46_24 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h18;
  wire          compressDataVec_hitReq_47_24 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h18;
  wire          compressDataVec_hitReq_48_24 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h18;
  wire          compressDataVec_hitReq_49_24 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h18;
  wire          compressDataVec_hitReq_50_24 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h18;
  wire          compressDataVec_hitReq_51_24 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h18;
  wire          compressDataVec_hitReq_52_24 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h18;
  wire          compressDataVec_hitReq_53_24 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h18;
  wire          compressDataVec_hitReq_54_24 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h18;
  wire          compressDataVec_hitReq_55_24 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h18;
  wire          compressDataVec_hitReq_56_24 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h18;
  wire          compressDataVec_hitReq_57_24 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h18;
  wire          compressDataVec_hitReq_58_24 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h18;
  wire          compressDataVec_hitReq_59_24 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h18;
  wire          compressDataVec_hitReq_60_24 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h18;
  wire          compressDataVec_hitReq_61_24 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h18;
  wire          compressDataVec_hitReq_62_24 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h18;
  wire          compressDataVec_hitReq_63_24 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h18;
  wire [7:0]    compressDataVec_selectReqData_24 =
    (compressDataVec_hitReq_0_24 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_24 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_24 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_24 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_24 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_24 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_24 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_24 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_24 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_24 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_24 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_24 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_24 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_24 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_24 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_24 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_24 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_24 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_24 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_24 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_24 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_24 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_24 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_24 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_24 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_24 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_24 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_24 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_24 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_24 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_24 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_24 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_24 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_24 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_24 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_24 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_24 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_24 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_24 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_24 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_24 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_24 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_24 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_24 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_24 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_24 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_24 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_24 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_24 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_24 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_24 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_24 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_24 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_24 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_24 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_24 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_24 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_24 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_24 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_24 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_24 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_24 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_24 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_24 ? source2Pipe[511:504] : 8'h0);
  wire          _GEN_819 = tailCount > 6'h18;
  wire          compressDataVec_useTail_24;
  assign compressDataVec_useTail_24 = _GEN_819;
  wire          compressDataVec_useTail_88;
  assign compressDataVec_useTail_88 = _GEN_819;
  wire          _GEN_820 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h19;
  wire          compressDataVec_hitReq_0_25;
  assign compressDataVec_hitReq_0_25 = _GEN_820;
  wire          compressDataVec_hitReq_0_153;
  assign compressDataVec_hitReq_0_153 = _GEN_820;
  wire          compressDataVec_hitReq_0_217;
  assign compressDataVec_hitReq_0_217 = _GEN_820;
  wire          _GEN_821 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h19;
  wire          compressDataVec_hitReq_1_25;
  assign compressDataVec_hitReq_1_25 = _GEN_821;
  wire          compressDataVec_hitReq_1_153;
  assign compressDataVec_hitReq_1_153 = _GEN_821;
  wire          compressDataVec_hitReq_1_217;
  assign compressDataVec_hitReq_1_217 = _GEN_821;
  wire          _GEN_822 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h19;
  wire          compressDataVec_hitReq_2_25;
  assign compressDataVec_hitReq_2_25 = _GEN_822;
  wire          compressDataVec_hitReq_2_153;
  assign compressDataVec_hitReq_2_153 = _GEN_822;
  wire          compressDataVec_hitReq_2_217;
  assign compressDataVec_hitReq_2_217 = _GEN_822;
  wire          _GEN_823 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h19;
  wire          compressDataVec_hitReq_3_25;
  assign compressDataVec_hitReq_3_25 = _GEN_823;
  wire          compressDataVec_hitReq_3_153;
  assign compressDataVec_hitReq_3_153 = _GEN_823;
  wire          compressDataVec_hitReq_3_217;
  assign compressDataVec_hitReq_3_217 = _GEN_823;
  wire          _GEN_824 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h19;
  wire          compressDataVec_hitReq_4_25;
  assign compressDataVec_hitReq_4_25 = _GEN_824;
  wire          compressDataVec_hitReq_4_153;
  assign compressDataVec_hitReq_4_153 = _GEN_824;
  wire          compressDataVec_hitReq_4_217;
  assign compressDataVec_hitReq_4_217 = _GEN_824;
  wire          _GEN_825 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h19;
  wire          compressDataVec_hitReq_5_25;
  assign compressDataVec_hitReq_5_25 = _GEN_825;
  wire          compressDataVec_hitReq_5_153;
  assign compressDataVec_hitReq_5_153 = _GEN_825;
  wire          compressDataVec_hitReq_5_217;
  assign compressDataVec_hitReq_5_217 = _GEN_825;
  wire          _GEN_826 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h19;
  wire          compressDataVec_hitReq_6_25;
  assign compressDataVec_hitReq_6_25 = _GEN_826;
  wire          compressDataVec_hitReq_6_153;
  assign compressDataVec_hitReq_6_153 = _GEN_826;
  wire          compressDataVec_hitReq_6_217;
  assign compressDataVec_hitReq_6_217 = _GEN_826;
  wire          _GEN_827 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h19;
  wire          compressDataVec_hitReq_7_25;
  assign compressDataVec_hitReq_7_25 = _GEN_827;
  wire          compressDataVec_hitReq_7_153;
  assign compressDataVec_hitReq_7_153 = _GEN_827;
  wire          compressDataVec_hitReq_7_217;
  assign compressDataVec_hitReq_7_217 = _GEN_827;
  wire          _GEN_828 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h19;
  wire          compressDataVec_hitReq_8_25;
  assign compressDataVec_hitReq_8_25 = _GEN_828;
  wire          compressDataVec_hitReq_8_153;
  assign compressDataVec_hitReq_8_153 = _GEN_828;
  wire          compressDataVec_hitReq_8_217;
  assign compressDataVec_hitReq_8_217 = _GEN_828;
  wire          _GEN_829 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h19;
  wire          compressDataVec_hitReq_9_25;
  assign compressDataVec_hitReq_9_25 = _GEN_829;
  wire          compressDataVec_hitReq_9_153;
  assign compressDataVec_hitReq_9_153 = _GEN_829;
  wire          compressDataVec_hitReq_9_217;
  assign compressDataVec_hitReq_9_217 = _GEN_829;
  wire          _GEN_830 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h19;
  wire          compressDataVec_hitReq_10_25;
  assign compressDataVec_hitReq_10_25 = _GEN_830;
  wire          compressDataVec_hitReq_10_153;
  assign compressDataVec_hitReq_10_153 = _GEN_830;
  wire          compressDataVec_hitReq_10_217;
  assign compressDataVec_hitReq_10_217 = _GEN_830;
  wire          _GEN_831 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h19;
  wire          compressDataVec_hitReq_11_25;
  assign compressDataVec_hitReq_11_25 = _GEN_831;
  wire          compressDataVec_hitReq_11_153;
  assign compressDataVec_hitReq_11_153 = _GEN_831;
  wire          compressDataVec_hitReq_11_217;
  assign compressDataVec_hitReq_11_217 = _GEN_831;
  wire          _GEN_832 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h19;
  wire          compressDataVec_hitReq_12_25;
  assign compressDataVec_hitReq_12_25 = _GEN_832;
  wire          compressDataVec_hitReq_12_153;
  assign compressDataVec_hitReq_12_153 = _GEN_832;
  wire          compressDataVec_hitReq_12_217;
  assign compressDataVec_hitReq_12_217 = _GEN_832;
  wire          _GEN_833 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h19;
  wire          compressDataVec_hitReq_13_25;
  assign compressDataVec_hitReq_13_25 = _GEN_833;
  wire          compressDataVec_hitReq_13_153;
  assign compressDataVec_hitReq_13_153 = _GEN_833;
  wire          compressDataVec_hitReq_13_217;
  assign compressDataVec_hitReq_13_217 = _GEN_833;
  wire          _GEN_834 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h19;
  wire          compressDataVec_hitReq_14_25;
  assign compressDataVec_hitReq_14_25 = _GEN_834;
  wire          compressDataVec_hitReq_14_153;
  assign compressDataVec_hitReq_14_153 = _GEN_834;
  wire          compressDataVec_hitReq_14_217;
  assign compressDataVec_hitReq_14_217 = _GEN_834;
  wire          _GEN_835 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h19;
  wire          compressDataVec_hitReq_15_25;
  assign compressDataVec_hitReq_15_25 = _GEN_835;
  wire          compressDataVec_hitReq_15_153;
  assign compressDataVec_hitReq_15_153 = _GEN_835;
  wire          compressDataVec_hitReq_15_217;
  assign compressDataVec_hitReq_15_217 = _GEN_835;
  wire          _GEN_836 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h19;
  wire          compressDataVec_hitReq_16_25;
  assign compressDataVec_hitReq_16_25 = _GEN_836;
  wire          compressDataVec_hitReq_16_153;
  assign compressDataVec_hitReq_16_153 = _GEN_836;
  wire          _GEN_837 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h19;
  wire          compressDataVec_hitReq_17_25;
  assign compressDataVec_hitReq_17_25 = _GEN_837;
  wire          compressDataVec_hitReq_17_153;
  assign compressDataVec_hitReq_17_153 = _GEN_837;
  wire          _GEN_838 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h19;
  wire          compressDataVec_hitReq_18_25;
  assign compressDataVec_hitReq_18_25 = _GEN_838;
  wire          compressDataVec_hitReq_18_153;
  assign compressDataVec_hitReq_18_153 = _GEN_838;
  wire          _GEN_839 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h19;
  wire          compressDataVec_hitReq_19_25;
  assign compressDataVec_hitReq_19_25 = _GEN_839;
  wire          compressDataVec_hitReq_19_153;
  assign compressDataVec_hitReq_19_153 = _GEN_839;
  wire          _GEN_840 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h19;
  wire          compressDataVec_hitReq_20_25;
  assign compressDataVec_hitReq_20_25 = _GEN_840;
  wire          compressDataVec_hitReq_20_153;
  assign compressDataVec_hitReq_20_153 = _GEN_840;
  wire          _GEN_841 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h19;
  wire          compressDataVec_hitReq_21_25;
  assign compressDataVec_hitReq_21_25 = _GEN_841;
  wire          compressDataVec_hitReq_21_153;
  assign compressDataVec_hitReq_21_153 = _GEN_841;
  wire          _GEN_842 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h19;
  wire          compressDataVec_hitReq_22_25;
  assign compressDataVec_hitReq_22_25 = _GEN_842;
  wire          compressDataVec_hitReq_22_153;
  assign compressDataVec_hitReq_22_153 = _GEN_842;
  wire          _GEN_843 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h19;
  wire          compressDataVec_hitReq_23_25;
  assign compressDataVec_hitReq_23_25 = _GEN_843;
  wire          compressDataVec_hitReq_23_153;
  assign compressDataVec_hitReq_23_153 = _GEN_843;
  wire          _GEN_844 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h19;
  wire          compressDataVec_hitReq_24_25;
  assign compressDataVec_hitReq_24_25 = _GEN_844;
  wire          compressDataVec_hitReq_24_153;
  assign compressDataVec_hitReq_24_153 = _GEN_844;
  wire          _GEN_845 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h19;
  wire          compressDataVec_hitReq_25_25;
  assign compressDataVec_hitReq_25_25 = _GEN_845;
  wire          compressDataVec_hitReq_25_153;
  assign compressDataVec_hitReq_25_153 = _GEN_845;
  wire          _GEN_846 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h19;
  wire          compressDataVec_hitReq_26_25;
  assign compressDataVec_hitReq_26_25 = _GEN_846;
  wire          compressDataVec_hitReq_26_153;
  assign compressDataVec_hitReq_26_153 = _GEN_846;
  wire          _GEN_847 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h19;
  wire          compressDataVec_hitReq_27_25;
  assign compressDataVec_hitReq_27_25 = _GEN_847;
  wire          compressDataVec_hitReq_27_153;
  assign compressDataVec_hitReq_27_153 = _GEN_847;
  wire          _GEN_848 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h19;
  wire          compressDataVec_hitReq_28_25;
  assign compressDataVec_hitReq_28_25 = _GEN_848;
  wire          compressDataVec_hitReq_28_153;
  assign compressDataVec_hitReq_28_153 = _GEN_848;
  wire          _GEN_849 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h19;
  wire          compressDataVec_hitReq_29_25;
  assign compressDataVec_hitReq_29_25 = _GEN_849;
  wire          compressDataVec_hitReq_29_153;
  assign compressDataVec_hitReq_29_153 = _GEN_849;
  wire          _GEN_850 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h19;
  wire          compressDataVec_hitReq_30_25;
  assign compressDataVec_hitReq_30_25 = _GEN_850;
  wire          compressDataVec_hitReq_30_153;
  assign compressDataVec_hitReq_30_153 = _GEN_850;
  wire          _GEN_851 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h19;
  wire          compressDataVec_hitReq_31_25;
  assign compressDataVec_hitReq_31_25 = _GEN_851;
  wire          compressDataVec_hitReq_31_153;
  assign compressDataVec_hitReq_31_153 = _GEN_851;
  wire          compressDataVec_hitReq_32_25 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h19;
  wire          compressDataVec_hitReq_33_25 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h19;
  wire          compressDataVec_hitReq_34_25 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h19;
  wire          compressDataVec_hitReq_35_25 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h19;
  wire          compressDataVec_hitReq_36_25 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h19;
  wire          compressDataVec_hitReq_37_25 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h19;
  wire          compressDataVec_hitReq_38_25 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h19;
  wire          compressDataVec_hitReq_39_25 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h19;
  wire          compressDataVec_hitReq_40_25 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h19;
  wire          compressDataVec_hitReq_41_25 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h19;
  wire          compressDataVec_hitReq_42_25 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h19;
  wire          compressDataVec_hitReq_43_25 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h19;
  wire          compressDataVec_hitReq_44_25 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h19;
  wire          compressDataVec_hitReq_45_25 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h19;
  wire          compressDataVec_hitReq_46_25 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h19;
  wire          compressDataVec_hitReq_47_25 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h19;
  wire          compressDataVec_hitReq_48_25 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h19;
  wire          compressDataVec_hitReq_49_25 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h19;
  wire          compressDataVec_hitReq_50_25 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h19;
  wire          compressDataVec_hitReq_51_25 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h19;
  wire          compressDataVec_hitReq_52_25 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h19;
  wire          compressDataVec_hitReq_53_25 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h19;
  wire          compressDataVec_hitReq_54_25 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h19;
  wire          compressDataVec_hitReq_55_25 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h19;
  wire          compressDataVec_hitReq_56_25 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h19;
  wire          compressDataVec_hitReq_57_25 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h19;
  wire          compressDataVec_hitReq_58_25 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h19;
  wire          compressDataVec_hitReq_59_25 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h19;
  wire          compressDataVec_hitReq_60_25 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h19;
  wire          compressDataVec_hitReq_61_25 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h19;
  wire          compressDataVec_hitReq_62_25 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h19;
  wire          compressDataVec_hitReq_63_25 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h19;
  wire [7:0]    compressDataVec_selectReqData_25 =
    (compressDataVec_hitReq_0_25 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_25 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_25 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_25 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_25 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_25 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_25 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_25 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_25 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_25 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_25 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_25 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_25 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_25 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_25 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_25 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_25 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_25 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_25 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_25 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_25 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_25 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_25 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_25 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_25 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_25 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_25 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_25 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_25 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_25 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_25 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_25 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_25 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_25 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_25 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_25 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_25 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_25 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_25 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_25 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_25 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_25 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_25 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_25 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_25 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_25 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_25 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_25 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_25 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_25 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_25 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_25 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_25 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_25 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_25 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_25 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_25 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_25 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_25 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_25 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_25 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_25 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_25 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_25 ? source2Pipe[511:504] : 8'h0);
  wire          _GEN_852 = tailCount > 6'h19;
  wire          compressDataVec_useTail_25;
  assign compressDataVec_useTail_25 = _GEN_852;
  wire          compressDataVec_useTail_89;
  assign compressDataVec_useTail_89 = _GEN_852;
  wire          _GEN_853 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h1A;
  wire          compressDataVec_hitReq_0_26;
  assign compressDataVec_hitReq_0_26 = _GEN_853;
  wire          compressDataVec_hitReq_0_154;
  assign compressDataVec_hitReq_0_154 = _GEN_853;
  wire          compressDataVec_hitReq_0_218;
  assign compressDataVec_hitReq_0_218 = _GEN_853;
  wire          _GEN_854 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h1A;
  wire          compressDataVec_hitReq_1_26;
  assign compressDataVec_hitReq_1_26 = _GEN_854;
  wire          compressDataVec_hitReq_1_154;
  assign compressDataVec_hitReq_1_154 = _GEN_854;
  wire          compressDataVec_hitReq_1_218;
  assign compressDataVec_hitReq_1_218 = _GEN_854;
  wire          _GEN_855 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h1A;
  wire          compressDataVec_hitReq_2_26;
  assign compressDataVec_hitReq_2_26 = _GEN_855;
  wire          compressDataVec_hitReq_2_154;
  assign compressDataVec_hitReq_2_154 = _GEN_855;
  wire          compressDataVec_hitReq_2_218;
  assign compressDataVec_hitReq_2_218 = _GEN_855;
  wire          _GEN_856 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h1A;
  wire          compressDataVec_hitReq_3_26;
  assign compressDataVec_hitReq_3_26 = _GEN_856;
  wire          compressDataVec_hitReq_3_154;
  assign compressDataVec_hitReq_3_154 = _GEN_856;
  wire          compressDataVec_hitReq_3_218;
  assign compressDataVec_hitReq_3_218 = _GEN_856;
  wire          _GEN_857 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h1A;
  wire          compressDataVec_hitReq_4_26;
  assign compressDataVec_hitReq_4_26 = _GEN_857;
  wire          compressDataVec_hitReq_4_154;
  assign compressDataVec_hitReq_4_154 = _GEN_857;
  wire          compressDataVec_hitReq_4_218;
  assign compressDataVec_hitReq_4_218 = _GEN_857;
  wire          _GEN_858 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h1A;
  wire          compressDataVec_hitReq_5_26;
  assign compressDataVec_hitReq_5_26 = _GEN_858;
  wire          compressDataVec_hitReq_5_154;
  assign compressDataVec_hitReq_5_154 = _GEN_858;
  wire          compressDataVec_hitReq_5_218;
  assign compressDataVec_hitReq_5_218 = _GEN_858;
  wire          _GEN_859 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h1A;
  wire          compressDataVec_hitReq_6_26;
  assign compressDataVec_hitReq_6_26 = _GEN_859;
  wire          compressDataVec_hitReq_6_154;
  assign compressDataVec_hitReq_6_154 = _GEN_859;
  wire          compressDataVec_hitReq_6_218;
  assign compressDataVec_hitReq_6_218 = _GEN_859;
  wire          _GEN_860 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h1A;
  wire          compressDataVec_hitReq_7_26;
  assign compressDataVec_hitReq_7_26 = _GEN_860;
  wire          compressDataVec_hitReq_7_154;
  assign compressDataVec_hitReq_7_154 = _GEN_860;
  wire          compressDataVec_hitReq_7_218;
  assign compressDataVec_hitReq_7_218 = _GEN_860;
  wire          _GEN_861 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h1A;
  wire          compressDataVec_hitReq_8_26;
  assign compressDataVec_hitReq_8_26 = _GEN_861;
  wire          compressDataVec_hitReq_8_154;
  assign compressDataVec_hitReq_8_154 = _GEN_861;
  wire          compressDataVec_hitReq_8_218;
  assign compressDataVec_hitReq_8_218 = _GEN_861;
  wire          _GEN_862 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h1A;
  wire          compressDataVec_hitReq_9_26;
  assign compressDataVec_hitReq_9_26 = _GEN_862;
  wire          compressDataVec_hitReq_9_154;
  assign compressDataVec_hitReq_9_154 = _GEN_862;
  wire          compressDataVec_hitReq_9_218;
  assign compressDataVec_hitReq_9_218 = _GEN_862;
  wire          _GEN_863 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h1A;
  wire          compressDataVec_hitReq_10_26;
  assign compressDataVec_hitReq_10_26 = _GEN_863;
  wire          compressDataVec_hitReq_10_154;
  assign compressDataVec_hitReq_10_154 = _GEN_863;
  wire          compressDataVec_hitReq_10_218;
  assign compressDataVec_hitReq_10_218 = _GEN_863;
  wire          _GEN_864 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h1A;
  wire          compressDataVec_hitReq_11_26;
  assign compressDataVec_hitReq_11_26 = _GEN_864;
  wire          compressDataVec_hitReq_11_154;
  assign compressDataVec_hitReq_11_154 = _GEN_864;
  wire          compressDataVec_hitReq_11_218;
  assign compressDataVec_hitReq_11_218 = _GEN_864;
  wire          _GEN_865 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h1A;
  wire          compressDataVec_hitReq_12_26;
  assign compressDataVec_hitReq_12_26 = _GEN_865;
  wire          compressDataVec_hitReq_12_154;
  assign compressDataVec_hitReq_12_154 = _GEN_865;
  wire          compressDataVec_hitReq_12_218;
  assign compressDataVec_hitReq_12_218 = _GEN_865;
  wire          _GEN_866 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h1A;
  wire          compressDataVec_hitReq_13_26;
  assign compressDataVec_hitReq_13_26 = _GEN_866;
  wire          compressDataVec_hitReq_13_154;
  assign compressDataVec_hitReq_13_154 = _GEN_866;
  wire          compressDataVec_hitReq_13_218;
  assign compressDataVec_hitReq_13_218 = _GEN_866;
  wire          _GEN_867 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h1A;
  wire          compressDataVec_hitReq_14_26;
  assign compressDataVec_hitReq_14_26 = _GEN_867;
  wire          compressDataVec_hitReq_14_154;
  assign compressDataVec_hitReq_14_154 = _GEN_867;
  wire          compressDataVec_hitReq_14_218;
  assign compressDataVec_hitReq_14_218 = _GEN_867;
  wire          _GEN_868 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h1A;
  wire          compressDataVec_hitReq_15_26;
  assign compressDataVec_hitReq_15_26 = _GEN_868;
  wire          compressDataVec_hitReq_15_154;
  assign compressDataVec_hitReq_15_154 = _GEN_868;
  wire          compressDataVec_hitReq_15_218;
  assign compressDataVec_hitReq_15_218 = _GEN_868;
  wire          _GEN_869 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h1A;
  wire          compressDataVec_hitReq_16_26;
  assign compressDataVec_hitReq_16_26 = _GEN_869;
  wire          compressDataVec_hitReq_16_154;
  assign compressDataVec_hitReq_16_154 = _GEN_869;
  wire          _GEN_870 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h1A;
  wire          compressDataVec_hitReq_17_26;
  assign compressDataVec_hitReq_17_26 = _GEN_870;
  wire          compressDataVec_hitReq_17_154;
  assign compressDataVec_hitReq_17_154 = _GEN_870;
  wire          _GEN_871 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h1A;
  wire          compressDataVec_hitReq_18_26;
  assign compressDataVec_hitReq_18_26 = _GEN_871;
  wire          compressDataVec_hitReq_18_154;
  assign compressDataVec_hitReq_18_154 = _GEN_871;
  wire          _GEN_872 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h1A;
  wire          compressDataVec_hitReq_19_26;
  assign compressDataVec_hitReq_19_26 = _GEN_872;
  wire          compressDataVec_hitReq_19_154;
  assign compressDataVec_hitReq_19_154 = _GEN_872;
  wire          _GEN_873 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h1A;
  wire          compressDataVec_hitReq_20_26;
  assign compressDataVec_hitReq_20_26 = _GEN_873;
  wire          compressDataVec_hitReq_20_154;
  assign compressDataVec_hitReq_20_154 = _GEN_873;
  wire          _GEN_874 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h1A;
  wire          compressDataVec_hitReq_21_26;
  assign compressDataVec_hitReq_21_26 = _GEN_874;
  wire          compressDataVec_hitReq_21_154;
  assign compressDataVec_hitReq_21_154 = _GEN_874;
  wire          _GEN_875 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h1A;
  wire          compressDataVec_hitReq_22_26;
  assign compressDataVec_hitReq_22_26 = _GEN_875;
  wire          compressDataVec_hitReq_22_154;
  assign compressDataVec_hitReq_22_154 = _GEN_875;
  wire          _GEN_876 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h1A;
  wire          compressDataVec_hitReq_23_26;
  assign compressDataVec_hitReq_23_26 = _GEN_876;
  wire          compressDataVec_hitReq_23_154;
  assign compressDataVec_hitReq_23_154 = _GEN_876;
  wire          _GEN_877 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h1A;
  wire          compressDataVec_hitReq_24_26;
  assign compressDataVec_hitReq_24_26 = _GEN_877;
  wire          compressDataVec_hitReq_24_154;
  assign compressDataVec_hitReq_24_154 = _GEN_877;
  wire          _GEN_878 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h1A;
  wire          compressDataVec_hitReq_25_26;
  assign compressDataVec_hitReq_25_26 = _GEN_878;
  wire          compressDataVec_hitReq_25_154;
  assign compressDataVec_hitReq_25_154 = _GEN_878;
  wire          _GEN_879 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h1A;
  wire          compressDataVec_hitReq_26_26;
  assign compressDataVec_hitReq_26_26 = _GEN_879;
  wire          compressDataVec_hitReq_26_154;
  assign compressDataVec_hitReq_26_154 = _GEN_879;
  wire          _GEN_880 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h1A;
  wire          compressDataVec_hitReq_27_26;
  assign compressDataVec_hitReq_27_26 = _GEN_880;
  wire          compressDataVec_hitReq_27_154;
  assign compressDataVec_hitReq_27_154 = _GEN_880;
  wire          _GEN_881 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h1A;
  wire          compressDataVec_hitReq_28_26;
  assign compressDataVec_hitReq_28_26 = _GEN_881;
  wire          compressDataVec_hitReq_28_154;
  assign compressDataVec_hitReq_28_154 = _GEN_881;
  wire          _GEN_882 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h1A;
  wire          compressDataVec_hitReq_29_26;
  assign compressDataVec_hitReq_29_26 = _GEN_882;
  wire          compressDataVec_hitReq_29_154;
  assign compressDataVec_hitReq_29_154 = _GEN_882;
  wire          _GEN_883 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h1A;
  wire          compressDataVec_hitReq_30_26;
  assign compressDataVec_hitReq_30_26 = _GEN_883;
  wire          compressDataVec_hitReq_30_154;
  assign compressDataVec_hitReq_30_154 = _GEN_883;
  wire          _GEN_884 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h1A;
  wire          compressDataVec_hitReq_31_26;
  assign compressDataVec_hitReq_31_26 = _GEN_884;
  wire          compressDataVec_hitReq_31_154;
  assign compressDataVec_hitReq_31_154 = _GEN_884;
  wire          compressDataVec_hitReq_32_26 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h1A;
  wire          compressDataVec_hitReq_33_26 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h1A;
  wire          compressDataVec_hitReq_34_26 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h1A;
  wire          compressDataVec_hitReq_35_26 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h1A;
  wire          compressDataVec_hitReq_36_26 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h1A;
  wire          compressDataVec_hitReq_37_26 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h1A;
  wire          compressDataVec_hitReq_38_26 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h1A;
  wire          compressDataVec_hitReq_39_26 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h1A;
  wire          compressDataVec_hitReq_40_26 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h1A;
  wire          compressDataVec_hitReq_41_26 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h1A;
  wire          compressDataVec_hitReq_42_26 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h1A;
  wire          compressDataVec_hitReq_43_26 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h1A;
  wire          compressDataVec_hitReq_44_26 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h1A;
  wire          compressDataVec_hitReq_45_26 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h1A;
  wire          compressDataVec_hitReq_46_26 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h1A;
  wire          compressDataVec_hitReq_47_26 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h1A;
  wire          compressDataVec_hitReq_48_26 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h1A;
  wire          compressDataVec_hitReq_49_26 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h1A;
  wire          compressDataVec_hitReq_50_26 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h1A;
  wire          compressDataVec_hitReq_51_26 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h1A;
  wire          compressDataVec_hitReq_52_26 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h1A;
  wire          compressDataVec_hitReq_53_26 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h1A;
  wire          compressDataVec_hitReq_54_26 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h1A;
  wire          compressDataVec_hitReq_55_26 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h1A;
  wire          compressDataVec_hitReq_56_26 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h1A;
  wire          compressDataVec_hitReq_57_26 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h1A;
  wire          compressDataVec_hitReq_58_26 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h1A;
  wire          compressDataVec_hitReq_59_26 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h1A;
  wire          compressDataVec_hitReq_60_26 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h1A;
  wire          compressDataVec_hitReq_61_26 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h1A;
  wire          compressDataVec_hitReq_62_26 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h1A;
  wire          compressDataVec_hitReq_63_26 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h1A;
  wire [7:0]    compressDataVec_selectReqData_26 =
    (compressDataVec_hitReq_0_26 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_26 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_26 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_26 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_26 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_26 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_26 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_26 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_26 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_26 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_26 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_26 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_26 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_26 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_26 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_26 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_26 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_26 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_26 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_26 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_26 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_26 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_26 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_26 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_26 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_26 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_26 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_26 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_26 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_26 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_26 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_26 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_26 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_26 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_26 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_26 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_26 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_26 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_26 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_26 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_26 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_26 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_26 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_26 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_26 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_26 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_26 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_26 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_26 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_26 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_26 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_26 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_26 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_26 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_26 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_26 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_26 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_26 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_26 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_26 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_26 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_26 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_26 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_26 ? source2Pipe[511:504] : 8'h0);
  wire          _GEN_885 = tailCount > 6'h1A;
  wire          compressDataVec_useTail_26;
  assign compressDataVec_useTail_26 = _GEN_885;
  wire          compressDataVec_useTail_90;
  assign compressDataVec_useTail_90 = _GEN_885;
  wire          _GEN_886 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h1B;
  wire          compressDataVec_hitReq_0_27;
  assign compressDataVec_hitReq_0_27 = _GEN_886;
  wire          compressDataVec_hitReq_0_155;
  assign compressDataVec_hitReq_0_155 = _GEN_886;
  wire          compressDataVec_hitReq_0_219;
  assign compressDataVec_hitReq_0_219 = _GEN_886;
  wire          _GEN_887 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h1B;
  wire          compressDataVec_hitReq_1_27;
  assign compressDataVec_hitReq_1_27 = _GEN_887;
  wire          compressDataVec_hitReq_1_155;
  assign compressDataVec_hitReq_1_155 = _GEN_887;
  wire          compressDataVec_hitReq_1_219;
  assign compressDataVec_hitReq_1_219 = _GEN_887;
  wire          _GEN_888 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h1B;
  wire          compressDataVec_hitReq_2_27;
  assign compressDataVec_hitReq_2_27 = _GEN_888;
  wire          compressDataVec_hitReq_2_155;
  assign compressDataVec_hitReq_2_155 = _GEN_888;
  wire          compressDataVec_hitReq_2_219;
  assign compressDataVec_hitReq_2_219 = _GEN_888;
  wire          _GEN_889 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h1B;
  wire          compressDataVec_hitReq_3_27;
  assign compressDataVec_hitReq_3_27 = _GEN_889;
  wire          compressDataVec_hitReq_3_155;
  assign compressDataVec_hitReq_3_155 = _GEN_889;
  wire          compressDataVec_hitReq_3_219;
  assign compressDataVec_hitReq_3_219 = _GEN_889;
  wire          _GEN_890 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h1B;
  wire          compressDataVec_hitReq_4_27;
  assign compressDataVec_hitReq_4_27 = _GEN_890;
  wire          compressDataVec_hitReq_4_155;
  assign compressDataVec_hitReq_4_155 = _GEN_890;
  wire          compressDataVec_hitReq_4_219;
  assign compressDataVec_hitReq_4_219 = _GEN_890;
  wire          _GEN_891 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h1B;
  wire          compressDataVec_hitReq_5_27;
  assign compressDataVec_hitReq_5_27 = _GEN_891;
  wire          compressDataVec_hitReq_5_155;
  assign compressDataVec_hitReq_5_155 = _GEN_891;
  wire          compressDataVec_hitReq_5_219;
  assign compressDataVec_hitReq_5_219 = _GEN_891;
  wire          _GEN_892 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h1B;
  wire          compressDataVec_hitReq_6_27;
  assign compressDataVec_hitReq_6_27 = _GEN_892;
  wire          compressDataVec_hitReq_6_155;
  assign compressDataVec_hitReq_6_155 = _GEN_892;
  wire          compressDataVec_hitReq_6_219;
  assign compressDataVec_hitReq_6_219 = _GEN_892;
  wire          _GEN_893 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h1B;
  wire          compressDataVec_hitReq_7_27;
  assign compressDataVec_hitReq_7_27 = _GEN_893;
  wire          compressDataVec_hitReq_7_155;
  assign compressDataVec_hitReq_7_155 = _GEN_893;
  wire          compressDataVec_hitReq_7_219;
  assign compressDataVec_hitReq_7_219 = _GEN_893;
  wire          _GEN_894 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h1B;
  wire          compressDataVec_hitReq_8_27;
  assign compressDataVec_hitReq_8_27 = _GEN_894;
  wire          compressDataVec_hitReq_8_155;
  assign compressDataVec_hitReq_8_155 = _GEN_894;
  wire          compressDataVec_hitReq_8_219;
  assign compressDataVec_hitReq_8_219 = _GEN_894;
  wire          _GEN_895 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h1B;
  wire          compressDataVec_hitReq_9_27;
  assign compressDataVec_hitReq_9_27 = _GEN_895;
  wire          compressDataVec_hitReq_9_155;
  assign compressDataVec_hitReq_9_155 = _GEN_895;
  wire          compressDataVec_hitReq_9_219;
  assign compressDataVec_hitReq_9_219 = _GEN_895;
  wire          _GEN_896 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h1B;
  wire          compressDataVec_hitReq_10_27;
  assign compressDataVec_hitReq_10_27 = _GEN_896;
  wire          compressDataVec_hitReq_10_155;
  assign compressDataVec_hitReq_10_155 = _GEN_896;
  wire          compressDataVec_hitReq_10_219;
  assign compressDataVec_hitReq_10_219 = _GEN_896;
  wire          _GEN_897 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h1B;
  wire          compressDataVec_hitReq_11_27;
  assign compressDataVec_hitReq_11_27 = _GEN_897;
  wire          compressDataVec_hitReq_11_155;
  assign compressDataVec_hitReq_11_155 = _GEN_897;
  wire          compressDataVec_hitReq_11_219;
  assign compressDataVec_hitReq_11_219 = _GEN_897;
  wire          _GEN_898 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h1B;
  wire          compressDataVec_hitReq_12_27;
  assign compressDataVec_hitReq_12_27 = _GEN_898;
  wire          compressDataVec_hitReq_12_155;
  assign compressDataVec_hitReq_12_155 = _GEN_898;
  wire          compressDataVec_hitReq_12_219;
  assign compressDataVec_hitReq_12_219 = _GEN_898;
  wire          _GEN_899 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h1B;
  wire          compressDataVec_hitReq_13_27;
  assign compressDataVec_hitReq_13_27 = _GEN_899;
  wire          compressDataVec_hitReq_13_155;
  assign compressDataVec_hitReq_13_155 = _GEN_899;
  wire          compressDataVec_hitReq_13_219;
  assign compressDataVec_hitReq_13_219 = _GEN_899;
  wire          _GEN_900 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h1B;
  wire          compressDataVec_hitReq_14_27;
  assign compressDataVec_hitReq_14_27 = _GEN_900;
  wire          compressDataVec_hitReq_14_155;
  assign compressDataVec_hitReq_14_155 = _GEN_900;
  wire          compressDataVec_hitReq_14_219;
  assign compressDataVec_hitReq_14_219 = _GEN_900;
  wire          _GEN_901 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h1B;
  wire          compressDataVec_hitReq_15_27;
  assign compressDataVec_hitReq_15_27 = _GEN_901;
  wire          compressDataVec_hitReq_15_155;
  assign compressDataVec_hitReq_15_155 = _GEN_901;
  wire          compressDataVec_hitReq_15_219;
  assign compressDataVec_hitReq_15_219 = _GEN_901;
  wire          _GEN_902 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h1B;
  wire          compressDataVec_hitReq_16_27;
  assign compressDataVec_hitReq_16_27 = _GEN_902;
  wire          compressDataVec_hitReq_16_155;
  assign compressDataVec_hitReq_16_155 = _GEN_902;
  wire          _GEN_903 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h1B;
  wire          compressDataVec_hitReq_17_27;
  assign compressDataVec_hitReq_17_27 = _GEN_903;
  wire          compressDataVec_hitReq_17_155;
  assign compressDataVec_hitReq_17_155 = _GEN_903;
  wire          _GEN_904 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h1B;
  wire          compressDataVec_hitReq_18_27;
  assign compressDataVec_hitReq_18_27 = _GEN_904;
  wire          compressDataVec_hitReq_18_155;
  assign compressDataVec_hitReq_18_155 = _GEN_904;
  wire          _GEN_905 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h1B;
  wire          compressDataVec_hitReq_19_27;
  assign compressDataVec_hitReq_19_27 = _GEN_905;
  wire          compressDataVec_hitReq_19_155;
  assign compressDataVec_hitReq_19_155 = _GEN_905;
  wire          _GEN_906 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h1B;
  wire          compressDataVec_hitReq_20_27;
  assign compressDataVec_hitReq_20_27 = _GEN_906;
  wire          compressDataVec_hitReq_20_155;
  assign compressDataVec_hitReq_20_155 = _GEN_906;
  wire          _GEN_907 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h1B;
  wire          compressDataVec_hitReq_21_27;
  assign compressDataVec_hitReq_21_27 = _GEN_907;
  wire          compressDataVec_hitReq_21_155;
  assign compressDataVec_hitReq_21_155 = _GEN_907;
  wire          _GEN_908 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h1B;
  wire          compressDataVec_hitReq_22_27;
  assign compressDataVec_hitReq_22_27 = _GEN_908;
  wire          compressDataVec_hitReq_22_155;
  assign compressDataVec_hitReq_22_155 = _GEN_908;
  wire          _GEN_909 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h1B;
  wire          compressDataVec_hitReq_23_27;
  assign compressDataVec_hitReq_23_27 = _GEN_909;
  wire          compressDataVec_hitReq_23_155;
  assign compressDataVec_hitReq_23_155 = _GEN_909;
  wire          _GEN_910 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h1B;
  wire          compressDataVec_hitReq_24_27;
  assign compressDataVec_hitReq_24_27 = _GEN_910;
  wire          compressDataVec_hitReq_24_155;
  assign compressDataVec_hitReq_24_155 = _GEN_910;
  wire          _GEN_911 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h1B;
  wire          compressDataVec_hitReq_25_27;
  assign compressDataVec_hitReq_25_27 = _GEN_911;
  wire          compressDataVec_hitReq_25_155;
  assign compressDataVec_hitReq_25_155 = _GEN_911;
  wire          _GEN_912 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h1B;
  wire          compressDataVec_hitReq_26_27;
  assign compressDataVec_hitReq_26_27 = _GEN_912;
  wire          compressDataVec_hitReq_26_155;
  assign compressDataVec_hitReq_26_155 = _GEN_912;
  wire          _GEN_913 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h1B;
  wire          compressDataVec_hitReq_27_27;
  assign compressDataVec_hitReq_27_27 = _GEN_913;
  wire          compressDataVec_hitReq_27_155;
  assign compressDataVec_hitReq_27_155 = _GEN_913;
  wire          _GEN_914 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h1B;
  wire          compressDataVec_hitReq_28_27;
  assign compressDataVec_hitReq_28_27 = _GEN_914;
  wire          compressDataVec_hitReq_28_155;
  assign compressDataVec_hitReq_28_155 = _GEN_914;
  wire          _GEN_915 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h1B;
  wire          compressDataVec_hitReq_29_27;
  assign compressDataVec_hitReq_29_27 = _GEN_915;
  wire          compressDataVec_hitReq_29_155;
  assign compressDataVec_hitReq_29_155 = _GEN_915;
  wire          _GEN_916 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h1B;
  wire          compressDataVec_hitReq_30_27;
  assign compressDataVec_hitReq_30_27 = _GEN_916;
  wire          compressDataVec_hitReq_30_155;
  assign compressDataVec_hitReq_30_155 = _GEN_916;
  wire          _GEN_917 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h1B;
  wire          compressDataVec_hitReq_31_27;
  assign compressDataVec_hitReq_31_27 = _GEN_917;
  wire          compressDataVec_hitReq_31_155;
  assign compressDataVec_hitReq_31_155 = _GEN_917;
  wire          compressDataVec_hitReq_32_27 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h1B;
  wire          compressDataVec_hitReq_33_27 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h1B;
  wire          compressDataVec_hitReq_34_27 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h1B;
  wire          compressDataVec_hitReq_35_27 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h1B;
  wire          compressDataVec_hitReq_36_27 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h1B;
  wire          compressDataVec_hitReq_37_27 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h1B;
  wire          compressDataVec_hitReq_38_27 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h1B;
  wire          compressDataVec_hitReq_39_27 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h1B;
  wire          compressDataVec_hitReq_40_27 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h1B;
  wire          compressDataVec_hitReq_41_27 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h1B;
  wire          compressDataVec_hitReq_42_27 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h1B;
  wire          compressDataVec_hitReq_43_27 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h1B;
  wire          compressDataVec_hitReq_44_27 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h1B;
  wire          compressDataVec_hitReq_45_27 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h1B;
  wire          compressDataVec_hitReq_46_27 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h1B;
  wire          compressDataVec_hitReq_47_27 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h1B;
  wire          compressDataVec_hitReq_48_27 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h1B;
  wire          compressDataVec_hitReq_49_27 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h1B;
  wire          compressDataVec_hitReq_50_27 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h1B;
  wire          compressDataVec_hitReq_51_27 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h1B;
  wire          compressDataVec_hitReq_52_27 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h1B;
  wire          compressDataVec_hitReq_53_27 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h1B;
  wire          compressDataVec_hitReq_54_27 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h1B;
  wire          compressDataVec_hitReq_55_27 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h1B;
  wire          compressDataVec_hitReq_56_27 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h1B;
  wire          compressDataVec_hitReq_57_27 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h1B;
  wire          compressDataVec_hitReq_58_27 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h1B;
  wire          compressDataVec_hitReq_59_27 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h1B;
  wire          compressDataVec_hitReq_60_27 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h1B;
  wire          compressDataVec_hitReq_61_27 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h1B;
  wire          compressDataVec_hitReq_62_27 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h1B;
  wire          compressDataVec_hitReq_63_27 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h1B;
  wire [7:0]    compressDataVec_selectReqData_27 =
    (compressDataVec_hitReq_0_27 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_27 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_27 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_27 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_27 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_27 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_27 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_27 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_27 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_27 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_27 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_27 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_27 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_27 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_27 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_27 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_27 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_27 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_27 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_27 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_27 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_27 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_27 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_27 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_27 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_27 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_27 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_27 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_27 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_27 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_27 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_27 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_27 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_27 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_27 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_27 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_27 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_27 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_27 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_27 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_27 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_27 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_27 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_27 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_27 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_27 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_27 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_27 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_27 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_27 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_27 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_27 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_27 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_27 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_27 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_27 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_27 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_27 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_27 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_27 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_27 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_27 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_27 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_27 ? source2Pipe[511:504] : 8'h0);
  wire          _GEN_918 = tailCount > 6'h1B;
  wire          compressDataVec_useTail_27;
  assign compressDataVec_useTail_27 = _GEN_918;
  wire          compressDataVec_useTail_91;
  assign compressDataVec_useTail_91 = _GEN_918;
  wire          _GEN_919 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h1C;
  wire          compressDataVec_hitReq_0_28;
  assign compressDataVec_hitReq_0_28 = _GEN_919;
  wire          compressDataVec_hitReq_0_156;
  assign compressDataVec_hitReq_0_156 = _GEN_919;
  wire          compressDataVec_hitReq_0_220;
  assign compressDataVec_hitReq_0_220 = _GEN_919;
  wire          _GEN_920 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h1C;
  wire          compressDataVec_hitReq_1_28;
  assign compressDataVec_hitReq_1_28 = _GEN_920;
  wire          compressDataVec_hitReq_1_156;
  assign compressDataVec_hitReq_1_156 = _GEN_920;
  wire          compressDataVec_hitReq_1_220;
  assign compressDataVec_hitReq_1_220 = _GEN_920;
  wire          _GEN_921 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h1C;
  wire          compressDataVec_hitReq_2_28;
  assign compressDataVec_hitReq_2_28 = _GEN_921;
  wire          compressDataVec_hitReq_2_156;
  assign compressDataVec_hitReq_2_156 = _GEN_921;
  wire          compressDataVec_hitReq_2_220;
  assign compressDataVec_hitReq_2_220 = _GEN_921;
  wire          _GEN_922 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h1C;
  wire          compressDataVec_hitReq_3_28;
  assign compressDataVec_hitReq_3_28 = _GEN_922;
  wire          compressDataVec_hitReq_3_156;
  assign compressDataVec_hitReq_3_156 = _GEN_922;
  wire          compressDataVec_hitReq_3_220;
  assign compressDataVec_hitReq_3_220 = _GEN_922;
  wire          _GEN_923 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h1C;
  wire          compressDataVec_hitReq_4_28;
  assign compressDataVec_hitReq_4_28 = _GEN_923;
  wire          compressDataVec_hitReq_4_156;
  assign compressDataVec_hitReq_4_156 = _GEN_923;
  wire          compressDataVec_hitReq_4_220;
  assign compressDataVec_hitReq_4_220 = _GEN_923;
  wire          _GEN_924 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h1C;
  wire          compressDataVec_hitReq_5_28;
  assign compressDataVec_hitReq_5_28 = _GEN_924;
  wire          compressDataVec_hitReq_5_156;
  assign compressDataVec_hitReq_5_156 = _GEN_924;
  wire          compressDataVec_hitReq_5_220;
  assign compressDataVec_hitReq_5_220 = _GEN_924;
  wire          _GEN_925 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h1C;
  wire          compressDataVec_hitReq_6_28;
  assign compressDataVec_hitReq_6_28 = _GEN_925;
  wire          compressDataVec_hitReq_6_156;
  assign compressDataVec_hitReq_6_156 = _GEN_925;
  wire          compressDataVec_hitReq_6_220;
  assign compressDataVec_hitReq_6_220 = _GEN_925;
  wire          _GEN_926 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h1C;
  wire          compressDataVec_hitReq_7_28;
  assign compressDataVec_hitReq_7_28 = _GEN_926;
  wire          compressDataVec_hitReq_7_156;
  assign compressDataVec_hitReq_7_156 = _GEN_926;
  wire          compressDataVec_hitReq_7_220;
  assign compressDataVec_hitReq_7_220 = _GEN_926;
  wire          _GEN_927 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h1C;
  wire          compressDataVec_hitReq_8_28;
  assign compressDataVec_hitReq_8_28 = _GEN_927;
  wire          compressDataVec_hitReq_8_156;
  assign compressDataVec_hitReq_8_156 = _GEN_927;
  wire          compressDataVec_hitReq_8_220;
  assign compressDataVec_hitReq_8_220 = _GEN_927;
  wire          _GEN_928 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h1C;
  wire          compressDataVec_hitReq_9_28;
  assign compressDataVec_hitReq_9_28 = _GEN_928;
  wire          compressDataVec_hitReq_9_156;
  assign compressDataVec_hitReq_9_156 = _GEN_928;
  wire          compressDataVec_hitReq_9_220;
  assign compressDataVec_hitReq_9_220 = _GEN_928;
  wire          _GEN_929 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h1C;
  wire          compressDataVec_hitReq_10_28;
  assign compressDataVec_hitReq_10_28 = _GEN_929;
  wire          compressDataVec_hitReq_10_156;
  assign compressDataVec_hitReq_10_156 = _GEN_929;
  wire          compressDataVec_hitReq_10_220;
  assign compressDataVec_hitReq_10_220 = _GEN_929;
  wire          _GEN_930 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h1C;
  wire          compressDataVec_hitReq_11_28;
  assign compressDataVec_hitReq_11_28 = _GEN_930;
  wire          compressDataVec_hitReq_11_156;
  assign compressDataVec_hitReq_11_156 = _GEN_930;
  wire          compressDataVec_hitReq_11_220;
  assign compressDataVec_hitReq_11_220 = _GEN_930;
  wire          _GEN_931 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h1C;
  wire          compressDataVec_hitReq_12_28;
  assign compressDataVec_hitReq_12_28 = _GEN_931;
  wire          compressDataVec_hitReq_12_156;
  assign compressDataVec_hitReq_12_156 = _GEN_931;
  wire          compressDataVec_hitReq_12_220;
  assign compressDataVec_hitReq_12_220 = _GEN_931;
  wire          _GEN_932 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h1C;
  wire          compressDataVec_hitReq_13_28;
  assign compressDataVec_hitReq_13_28 = _GEN_932;
  wire          compressDataVec_hitReq_13_156;
  assign compressDataVec_hitReq_13_156 = _GEN_932;
  wire          compressDataVec_hitReq_13_220;
  assign compressDataVec_hitReq_13_220 = _GEN_932;
  wire          _GEN_933 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h1C;
  wire          compressDataVec_hitReq_14_28;
  assign compressDataVec_hitReq_14_28 = _GEN_933;
  wire          compressDataVec_hitReq_14_156;
  assign compressDataVec_hitReq_14_156 = _GEN_933;
  wire          compressDataVec_hitReq_14_220;
  assign compressDataVec_hitReq_14_220 = _GEN_933;
  wire          _GEN_934 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h1C;
  wire          compressDataVec_hitReq_15_28;
  assign compressDataVec_hitReq_15_28 = _GEN_934;
  wire          compressDataVec_hitReq_15_156;
  assign compressDataVec_hitReq_15_156 = _GEN_934;
  wire          compressDataVec_hitReq_15_220;
  assign compressDataVec_hitReq_15_220 = _GEN_934;
  wire          _GEN_935 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h1C;
  wire          compressDataVec_hitReq_16_28;
  assign compressDataVec_hitReq_16_28 = _GEN_935;
  wire          compressDataVec_hitReq_16_156;
  assign compressDataVec_hitReq_16_156 = _GEN_935;
  wire          _GEN_936 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h1C;
  wire          compressDataVec_hitReq_17_28;
  assign compressDataVec_hitReq_17_28 = _GEN_936;
  wire          compressDataVec_hitReq_17_156;
  assign compressDataVec_hitReq_17_156 = _GEN_936;
  wire          _GEN_937 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h1C;
  wire          compressDataVec_hitReq_18_28;
  assign compressDataVec_hitReq_18_28 = _GEN_937;
  wire          compressDataVec_hitReq_18_156;
  assign compressDataVec_hitReq_18_156 = _GEN_937;
  wire          _GEN_938 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h1C;
  wire          compressDataVec_hitReq_19_28;
  assign compressDataVec_hitReq_19_28 = _GEN_938;
  wire          compressDataVec_hitReq_19_156;
  assign compressDataVec_hitReq_19_156 = _GEN_938;
  wire          _GEN_939 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h1C;
  wire          compressDataVec_hitReq_20_28;
  assign compressDataVec_hitReq_20_28 = _GEN_939;
  wire          compressDataVec_hitReq_20_156;
  assign compressDataVec_hitReq_20_156 = _GEN_939;
  wire          _GEN_940 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h1C;
  wire          compressDataVec_hitReq_21_28;
  assign compressDataVec_hitReq_21_28 = _GEN_940;
  wire          compressDataVec_hitReq_21_156;
  assign compressDataVec_hitReq_21_156 = _GEN_940;
  wire          _GEN_941 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h1C;
  wire          compressDataVec_hitReq_22_28;
  assign compressDataVec_hitReq_22_28 = _GEN_941;
  wire          compressDataVec_hitReq_22_156;
  assign compressDataVec_hitReq_22_156 = _GEN_941;
  wire          _GEN_942 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h1C;
  wire          compressDataVec_hitReq_23_28;
  assign compressDataVec_hitReq_23_28 = _GEN_942;
  wire          compressDataVec_hitReq_23_156;
  assign compressDataVec_hitReq_23_156 = _GEN_942;
  wire          _GEN_943 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h1C;
  wire          compressDataVec_hitReq_24_28;
  assign compressDataVec_hitReq_24_28 = _GEN_943;
  wire          compressDataVec_hitReq_24_156;
  assign compressDataVec_hitReq_24_156 = _GEN_943;
  wire          _GEN_944 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h1C;
  wire          compressDataVec_hitReq_25_28;
  assign compressDataVec_hitReq_25_28 = _GEN_944;
  wire          compressDataVec_hitReq_25_156;
  assign compressDataVec_hitReq_25_156 = _GEN_944;
  wire          _GEN_945 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h1C;
  wire          compressDataVec_hitReq_26_28;
  assign compressDataVec_hitReq_26_28 = _GEN_945;
  wire          compressDataVec_hitReq_26_156;
  assign compressDataVec_hitReq_26_156 = _GEN_945;
  wire          _GEN_946 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h1C;
  wire          compressDataVec_hitReq_27_28;
  assign compressDataVec_hitReq_27_28 = _GEN_946;
  wire          compressDataVec_hitReq_27_156;
  assign compressDataVec_hitReq_27_156 = _GEN_946;
  wire          _GEN_947 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h1C;
  wire          compressDataVec_hitReq_28_28;
  assign compressDataVec_hitReq_28_28 = _GEN_947;
  wire          compressDataVec_hitReq_28_156;
  assign compressDataVec_hitReq_28_156 = _GEN_947;
  wire          _GEN_948 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h1C;
  wire          compressDataVec_hitReq_29_28;
  assign compressDataVec_hitReq_29_28 = _GEN_948;
  wire          compressDataVec_hitReq_29_156;
  assign compressDataVec_hitReq_29_156 = _GEN_948;
  wire          _GEN_949 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h1C;
  wire          compressDataVec_hitReq_30_28;
  assign compressDataVec_hitReq_30_28 = _GEN_949;
  wire          compressDataVec_hitReq_30_156;
  assign compressDataVec_hitReq_30_156 = _GEN_949;
  wire          _GEN_950 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h1C;
  wire          compressDataVec_hitReq_31_28;
  assign compressDataVec_hitReq_31_28 = _GEN_950;
  wire          compressDataVec_hitReq_31_156;
  assign compressDataVec_hitReq_31_156 = _GEN_950;
  wire          compressDataVec_hitReq_32_28 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h1C;
  wire          compressDataVec_hitReq_33_28 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h1C;
  wire          compressDataVec_hitReq_34_28 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h1C;
  wire          compressDataVec_hitReq_35_28 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h1C;
  wire          compressDataVec_hitReq_36_28 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h1C;
  wire          compressDataVec_hitReq_37_28 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h1C;
  wire          compressDataVec_hitReq_38_28 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h1C;
  wire          compressDataVec_hitReq_39_28 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h1C;
  wire          compressDataVec_hitReq_40_28 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h1C;
  wire          compressDataVec_hitReq_41_28 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h1C;
  wire          compressDataVec_hitReq_42_28 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h1C;
  wire          compressDataVec_hitReq_43_28 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h1C;
  wire          compressDataVec_hitReq_44_28 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h1C;
  wire          compressDataVec_hitReq_45_28 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h1C;
  wire          compressDataVec_hitReq_46_28 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h1C;
  wire          compressDataVec_hitReq_47_28 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h1C;
  wire          compressDataVec_hitReq_48_28 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h1C;
  wire          compressDataVec_hitReq_49_28 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h1C;
  wire          compressDataVec_hitReq_50_28 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h1C;
  wire          compressDataVec_hitReq_51_28 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h1C;
  wire          compressDataVec_hitReq_52_28 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h1C;
  wire          compressDataVec_hitReq_53_28 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h1C;
  wire          compressDataVec_hitReq_54_28 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h1C;
  wire          compressDataVec_hitReq_55_28 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h1C;
  wire          compressDataVec_hitReq_56_28 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h1C;
  wire          compressDataVec_hitReq_57_28 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h1C;
  wire          compressDataVec_hitReq_58_28 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h1C;
  wire          compressDataVec_hitReq_59_28 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h1C;
  wire          compressDataVec_hitReq_60_28 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h1C;
  wire          compressDataVec_hitReq_61_28 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h1C;
  wire          compressDataVec_hitReq_62_28 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h1C;
  wire          compressDataVec_hitReq_63_28 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h1C;
  wire [7:0]    compressDataVec_selectReqData_28 =
    (compressDataVec_hitReq_0_28 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_28 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_28 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_28 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_28 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_28 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_28 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_28 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_28 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_28 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_28 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_28 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_28 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_28 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_28 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_28 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_28 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_28 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_28 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_28 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_28 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_28 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_28 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_28 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_28 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_28 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_28 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_28 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_28 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_28 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_28 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_28 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_28 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_28 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_28 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_28 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_28 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_28 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_28 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_28 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_28 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_28 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_28 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_28 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_28 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_28 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_28 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_28 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_28 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_28 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_28 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_28 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_28 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_28 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_28 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_28 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_28 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_28 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_28 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_28 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_28 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_28 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_28 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_28 ? source2Pipe[511:504] : 8'h0);
  wire          _GEN_951 = tailCount > 6'h1C;
  wire          compressDataVec_useTail_28;
  assign compressDataVec_useTail_28 = _GEN_951;
  wire          compressDataVec_useTail_92;
  assign compressDataVec_useTail_92 = _GEN_951;
  wire          _GEN_952 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h1D;
  wire          compressDataVec_hitReq_0_29;
  assign compressDataVec_hitReq_0_29 = _GEN_952;
  wire          compressDataVec_hitReq_0_157;
  assign compressDataVec_hitReq_0_157 = _GEN_952;
  wire          compressDataVec_hitReq_0_221;
  assign compressDataVec_hitReq_0_221 = _GEN_952;
  wire          _GEN_953 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h1D;
  wire          compressDataVec_hitReq_1_29;
  assign compressDataVec_hitReq_1_29 = _GEN_953;
  wire          compressDataVec_hitReq_1_157;
  assign compressDataVec_hitReq_1_157 = _GEN_953;
  wire          compressDataVec_hitReq_1_221;
  assign compressDataVec_hitReq_1_221 = _GEN_953;
  wire          _GEN_954 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h1D;
  wire          compressDataVec_hitReq_2_29;
  assign compressDataVec_hitReq_2_29 = _GEN_954;
  wire          compressDataVec_hitReq_2_157;
  assign compressDataVec_hitReq_2_157 = _GEN_954;
  wire          compressDataVec_hitReq_2_221;
  assign compressDataVec_hitReq_2_221 = _GEN_954;
  wire          _GEN_955 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h1D;
  wire          compressDataVec_hitReq_3_29;
  assign compressDataVec_hitReq_3_29 = _GEN_955;
  wire          compressDataVec_hitReq_3_157;
  assign compressDataVec_hitReq_3_157 = _GEN_955;
  wire          compressDataVec_hitReq_3_221;
  assign compressDataVec_hitReq_3_221 = _GEN_955;
  wire          _GEN_956 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h1D;
  wire          compressDataVec_hitReq_4_29;
  assign compressDataVec_hitReq_4_29 = _GEN_956;
  wire          compressDataVec_hitReq_4_157;
  assign compressDataVec_hitReq_4_157 = _GEN_956;
  wire          compressDataVec_hitReq_4_221;
  assign compressDataVec_hitReq_4_221 = _GEN_956;
  wire          _GEN_957 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h1D;
  wire          compressDataVec_hitReq_5_29;
  assign compressDataVec_hitReq_5_29 = _GEN_957;
  wire          compressDataVec_hitReq_5_157;
  assign compressDataVec_hitReq_5_157 = _GEN_957;
  wire          compressDataVec_hitReq_5_221;
  assign compressDataVec_hitReq_5_221 = _GEN_957;
  wire          _GEN_958 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h1D;
  wire          compressDataVec_hitReq_6_29;
  assign compressDataVec_hitReq_6_29 = _GEN_958;
  wire          compressDataVec_hitReq_6_157;
  assign compressDataVec_hitReq_6_157 = _GEN_958;
  wire          compressDataVec_hitReq_6_221;
  assign compressDataVec_hitReq_6_221 = _GEN_958;
  wire          _GEN_959 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h1D;
  wire          compressDataVec_hitReq_7_29;
  assign compressDataVec_hitReq_7_29 = _GEN_959;
  wire          compressDataVec_hitReq_7_157;
  assign compressDataVec_hitReq_7_157 = _GEN_959;
  wire          compressDataVec_hitReq_7_221;
  assign compressDataVec_hitReq_7_221 = _GEN_959;
  wire          _GEN_960 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h1D;
  wire          compressDataVec_hitReq_8_29;
  assign compressDataVec_hitReq_8_29 = _GEN_960;
  wire          compressDataVec_hitReq_8_157;
  assign compressDataVec_hitReq_8_157 = _GEN_960;
  wire          compressDataVec_hitReq_8_221;
  assign compressDataVec_hitReq_8_221 = _GEN_960;
  wire          _GEN_961 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h1D;
  wire          compressDataVec_hitReq_9_29;
  assign compressDataVec_hitReq_9_29 = _GEN_961;
  wire          compressDataVec_hitReq_9_157;
  assign compressDataVec_hitReq_9_157 = _GEN_961;
  wire          compressDataVec_hitReq_9_221;
  assign compressDataVec_hitReq_9_221 = _GEN_961;
  wire          _GEN_962 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h1D;
  wire          compressDataVec_hitReq_10_29;
  assign compressDataVec_hitReq_10_29 = _GEN_962;
  wire          compressDataVec_hitReq_10_157;
  assign compressDataVec_hitReq_10_157 = _GEN_962;
  wire          compressDataVec_hitReq_10_221;
  assign compressDataVec_hitReq_10_221 = _GEN_962;
  wire          _GEN_963 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h1D;
  wire          compressDataVec_hitReq_11_29;
  assign compressDataVec_hitReq_11_29 = _GEN_963;
  wire          compressDataVec_hitReq_11_157;
  assign compressDataVec_hitReq_11_157 = _GEN_963;
  wire          compressDataVec_hitReq_11_221;
  assign compressDataVec_hitReq_11_221 = _GEN_963;
  wire          _GEN_964 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h1D;
  wire          compressDataVec_hitReq_12_29;
  assign compressDataVec_hitReq_12_29 = _GEN_964;
  wire          compressDataVec_hitReq_12_157;
  assign compressDataVec_hitReq_12_157 = _GEN_964;
  wire          compressDataVec_hitReq_12_221;
  assign compressDataVec_hitReq_12_221 = _GEN_964;
  wire          _GEN_965 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h1D;
  wire          compressDataVec_hitReq_13_29;
  assign compressDataVec_hitReq_13_29 = _GEN_965;
  wire          compressDataVec_hitReq_13_157;
  assign compressDataVec_hitReq_13_157 = _GEN_965;
  wire          compressDataVec_hitReq_13_221;
  assign compressDataVec_hitReq_13_221 = _GEN_965;
  wire          _GEN_966 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h1D;
  wire          compressDataVec_hitReq_14_29;
  assign compressDataVec_hitReq_14_29 = _GEN_966;
  wire          compressDataVec_hitReq_14_157;
  assign compressDataVec_hitReq_14_157 = _GEN_966;
  wire          compressDataVec_hitReq_14_221;
  assign compressDataVec_hitReq_14_221 = _GEN_966;
  wire          _GEN_967 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h1D;
  wire          compressDataVec_hitReq_15_29;
  assign compressDataVec_hitReq_15_29 = _GEN_967;
  wire          compressDataVec_hitReq_15_157;
  assign compressDataVec_hitReq_15_157 = _GEN_967;
  wire          compressDataVec_hitReq_15_221;
  assign compressDataVec_hitReq_15_221 = _GEN_967;
  wire          _GEN_968 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h1D;
  wire          compressDataVec_hitReq_16_29;
  assign compressDataVec_hitReq_16_29 = _GEN_968;
  wire          compressDataVec_hitReq_16_157;
  assign compressDataVec_hitReq_16_157 = _GEN_968;
  wire          _GEN_969 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h1D;
  wire          compressDataVec_hitReq_17_29;
  assign compressDataVec_hitReq_17_29 = _GEN_969;
  wire          compressDataVec_hitReq_17_157;
  assign compressDataVec_hitReq_17_157 = _GEN_969;
  wire          _GEN_970 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h1D;
  wire          compressDataVec_hitReq_18_29;
  assign compressDataVec_hitReq_18_29 = _GEN_970;
  wire          compressDataVec_hitReq_18_157;
  assign compressDataVec_hitReq_18_157 = _GEN_970;
  wire          _GEN_971 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h1D;
  wire          compressDataVec_hitReq_19_29;
  assign compressDataVec_hitReq_19_29 = _GEN_971;
  wire          compressDataVec_hitReq_19_157;
  assign compressDataVec_hitReq_19_157 = _GEN_971;
  wire          _GEN_972 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h1D;
  wire          compressDataVec_hitReq_20_29;
  assign compressDataVec_hitReq_20_29 = _GEN_972;
  wire          compressDataVec_hitReq_20_157;
  assign compressDataVec_hitReq_20_157 = _GEN_972;
  wire          _GEN_973 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h1D;
  wire          compressDataVec_hitReq_21_29;
  assign compressDataVec_hitReq_21_29 = _GEN_973;
  wire          compressDataVec_hitReq_21_157;
  assign compressDataVec_hitReq_21_157 = _GEN_973;
  wire          _GEN_974 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h1D;
  wire          compressDataVec_hitReq_22_29;
  assign compressDataVec_hitReq_22_29 = _GEN_974;
  wire          compressDataVec_hitReq_22_157;
  assign compressDataVec_hitReq_22_157 = _GEN_974;
  wire          _GEN_975 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h1D;
  wire          compressDataVec_hitReq_23_29;
  assign compressDataVec_hitReq_23_29 = _GEN_975;
  wire          compressDataVec_hitReq_23_157;
  assign compressDataVec_hitReq_23_157 = _GEN_975;
  wire          _GEN_976 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h1D;
  wire          compressDataVec_hitReq_24_29;
  assign compressDataVec_hitReq_24_29 = _GEN_976;
  wire          compressDataVec_hitReq_24_157;
  assign compressDataVec_hitReq_24_157 = _GEN_976;
  wire          _GEN_977 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h1D;
  wire          compressDataVec_hitReq_25_29;
  assign compressDataVec_hitReq_25_29 = _GEN_977;
  wire          compressDataVec_hitReq_25_157;
  assign compressDataVec_hitReq_25_157 = _GEN_977;
  wire          _GEN_978 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h1D;
  wire          compressDataVec_hitReq_26_29;
  assign compressDataVec_hitReq_26_29 = _GEN_978;
  wire          compressDataVec_hitReq_26_157;
  assign compressDataVec_hitReq_26_157 = _GEN_978;
  wire          _GEN_979 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h1D;
  wire          compressDataVec_hitReq_27_29;
  assign compressDataVec_hitReq_27_29 = _GEN_979;
  wire          compressDataVec_hitReq_27_157;
  assign compressDataVec_hitReq_27_157 = _GEN_979;
  wire          _GEN_980 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h1D;
  wire          compressDataVec_hitReq_28_29;
  assign compressDataVec_hitReq_28_29 = _GEN_980;
  wire          compressDataVec_hitReq_28_157;
  assign compressDataVec_hitReq_28_157 = _GEN_980;
  wire          _GEN_981 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h1D;
  wire          compressDataVec_hitReq_29_29;
  assign compressDataVec_hitReq_29_29 = _GEN_981;
  wire          compressDataVec_hitReq_29_157;
  assign compressDataVec_hitReq_29_157 = _GEN_981;
  wire          _GEN_982 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h1D;
  wire          compressDataVec_hitReq_30_29;
  assign compressDataVec_hitReq_30_29 = _GEN_982;
  wire          compressDataVec_hitReq_30_157;
  assign compressDataVec_hitReq_30_157 = _GEN_982;
  wire          _GEN_983 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h1D;
  wire          compressDataVec_hitReq_31_29;
  assign compressDataVec_hitReq_31_29 = _GEN_983;
  wire          compressDataVec_hitReq_31_157;
  assign compressDataVec_hitReq_31_157 = _GEN_983;
  wire          compressDataVec_hitReq_32_29 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h1D;
  wire          compressDataVec_hitReq_33_29 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h1D;
  wire          compressDataVec_hitReq_34_29 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h1D;
  wire          compressDataVec_hitReq_35_29 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h1D;
  wire          compressDataVec_hitReq_36_29 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h1D;
  wire          compressDataVec_hitReq_37_29 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h1D;
  wire          compressDataVec_hitReq_38_29 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h1D;
  wire          compressDataVec_hitReq_39_29 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h1D;
  wire          compressDataVec_hitReq_40_29 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h1D;
  wire          compressDataVec_hitReq_41_29 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h1D;
  wire          compressDataVec_hitReq_42_29 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h1D;
  wire          compressDataVec_hitReq_43_29 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h1D;
  wire          compressDataVec_hitReq_44_29 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h1D;
  wire          compressDataVec_hitReq_45_29 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h1D;
  wire          compressDataVec_hitReq_46_29 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h1D;
  wire          compressDataVec_hitReq_47_29 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h1D;
  wire          compressDataVec_hitReq_48_29 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h1D;
  wire          compressDataVec_hitReq_49_29 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h1D;
  wire          compressDataVec_hitReq_50_29 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h1D;
  wire          compressDataVec_hitReq_51_29 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h1D;
  wire          compressDataVec_hitReq_52_29 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h1D;
  wire          compressDataVec_hitReq_53_29 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h1D;
  wire          compressDataVec_hitReq_54_29 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h1D;
  wire          compressDataVec_hitReq_55_29 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h1D;
  wire          compressDataVec_hitReq_56_29 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h1D;
  wire          compressDataVec_hitReq_57_29 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h1D;
  wire          compressDataVec_hitReq_58_29 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h1D;
  wire          compressDataVec_hitReq_59_29 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h1D;
  wire          compressDataVec_hitReq_60_29 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h1D;
  wire          compressDataVec_hitReq_61_29 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h1D;
  wire          compressDataVec_hitReq_62_29 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h1D;
  wire          compressDataVec_hitReq_63_29 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h1D;
  wire [7:0]    compressDataVec_selectReqData_29 =
    (compressDataVec_hitReq_0_29 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_29 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_29 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_29 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_29 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_29 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_29 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_29 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_29 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_29 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_29 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_29 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_29 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_29 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_29 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_29 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_29 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_29 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_29 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_29 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_29 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_29 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_29 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_29 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_29 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_29 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_29 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_29 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_29 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_29 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_29 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_29 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_29 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_29 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_29 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_29 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_29 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_29 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_29 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_29 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_29 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_29 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_29 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_29 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_29 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_29 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_29 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_29 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_29 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_29 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_29 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_29 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_29 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_29 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_29 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_29 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_29 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_29 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_29 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_29 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_29 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_29 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_29 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_29 ? source2Pipe[511:504] : 8'h0);
  wire          _GEN_984 = tailCount > 6'h1D;
  wire          compressDataVec_useTail_29;
  assign compressDataVec_useTail_29 = _GEN_984;
  wire          compressDataVec_useTail_93;
  assign compressDataVec_useTail_93 = _GEN_984;
  wire          _GEN_985 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h1E;
  wire          compressDataVec_hitReq_0_30;
  assign compressDataVec_hitReq_0_30 = _GEN_985;
  wire          compressDataVec_hitReq_0_158;
  assign compressDataVec_hitReq_0_158 = _GEN_985;
  wire          compressDataVec_hitReq_0_222;
  assign compressDataVec_hitReq_0_222 = _GEN_985;
  wire          _GEN_986 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h1E;
  wire          compressDataVec_hitReq_1_30;
  assign compressDataVec_hitReq_1_30 = _GEN_986;
  wire          compressDataVec_hitReq_1_158;
  assign compressDataVec_hitReq_1_158 = _GEN_986;
  wire          compressDataVec_hitReq_1_222;
  assign compressDataVec_hitReq_1_222 = _GEN_986;
  wire          _GEN_987 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h1E;
  wire          compressDataVec_hitReq_2_30;
  assign compressDataVec_hitReq_2_30 = _GEN_987;
  wire          compressDataVec_hitReq_2_158;
  assign compressDataVec_hitReq_2_158 = _GEN_987;
  wire          compressDataVec_hitReq_2_222;
  assign compressDataVec_hitReq_2_222 = _GEN_987;
  wire          _GEN_988 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h1E;
  wire          compressDataVec_hitReq_3_30;
  assign compressDataVec_hitReq_3_30 = _GEN_988;
  wire          compressDataVec_hitReq_3_158;
  assign compressDataVec_hitReq_3_158 = _GEN_988;
  wire          compressDataVec_hitReq_3_222;
  assign compressDataVec_hitReq_3_222 = _GEN_988;
  wire          _GEN_989 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h1E;
  wire          compressDataVec_hitReq_4_30;
  assign compressDataVec_hitReq_4_30 = _GEN_989;
  wire          compressDataVec_hitReq_4_158;
  assign compressDataVec_hitReq_4_158 = _GEN_989;
  wire          compressDataVec_hitReq_4_222;
  assign compressDataVec_hitReq_4_222 = _GEN_989;
  wire          _GEN_990 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h1E;
  wire          compressDataVec_hitReq_5_30;
  assign compressDataVec_hitReq_5_30 = _GEN_990;
  wire          compressDataVec_hitReq_5_158;
  assign compressDataVec_hitReq_5_158 = _GEN_990;
  wire          compressDataVec_hitReq_5_222;
  assign compressDataVec_hitReq_5_222 = _GEN_990;
  wire          _GEN_991 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h1E;
  wire          compressDataVec_hitReq_6_30;
  assign compressDataVec_hitReq_6_30 = _GEN_991;
  wire          compressDataVec_hitReq_6_158;
  assign compressDataVec_hitReq_6_158 = _GEN_991;
  wire          compressDataVec_hitReq_6_222;
  assign compressDataVec_hitReq_6_222 = _GEN_991;
  wire          _GEN_992 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h1E;
  wire          compressDataVec_hitReq_7_30;
  assign compressDataVec_hitReq_7_30 = _GEN_992;
  wire          compressDataVec_hitReq_7_158;
  assign compressDataVec_hitReq_7_158 = _GEN_992;
  wire          compressDataVec_hitReq_7_222;
  assign compressDataVec_hitReq_7_222 = _GEN_992;
  wire          _GEN_993 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h1E;
  wire          compressDataVec_hitReq_8_30;
  assign compressDataVec_hitReq_8_30 = _GEN_993;
  wire          compressDataVec_hitReq_8_158;
  assign compressDataVec_hitReq_8_158 = _GEN_993;
  wire          compressDataVec_hitReq_8_222;
  assign compressDataVec_hitReq_8_222 = _GEN_993;
  wire          _GEN_994 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h1E;
  wire          compressDataVec_hitReq_9_30;
  assign compressDataVec_hitReq_9_30 = _GEN_994;
  wire          compressDataVec_hitReq_9_158;
  assign compressDataVec_hitReq_9_158 = _GEN_994;
  wire          compressDataVec_hitReq_9_222;
  assign compressDataVec_hitReq_9_222 = _GEN_994;
  wire          _GEN_995 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h1E;
  wire          compressDataVec_hitReq_10_30;
  assign compressDataVec_hitReq_10_30 = _GEN_995;
  wire          compressDataVec_hitReq_10_158;
  assign compressDataVec_hitReq_10_158 = _GEN_995;
  wire          compressDataVec_hitReq_10_222;
  assign compressDataVec_hitReq_10_222 = _GEN_995;
  wire          _GEN_996 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h1E;
  wire          compressDataVec_hitReq_11_30;
  assign compressDataVec_hitReq_11_30 = _GEN_996;
  wire          compressDataVec_hitReq_11_158;
  assign compressDataVec_hitReq_11_158 = _GEN_996;
  wire          compressDataVec_hitReq_11_222;
  assign compressDataVec_hitReq_11_222 = _GEN_996;
  wire          _GEN_997 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h1E;
  wire          compressDataVec_hitReq_12_30;
  assign compressDataVec_hitReq_12_30 = _GEN_997;
  wire          compressDataVec_hitReq_12_158;
  assign compressDataVec_hitReq_12_158 = _GEN_997;
  wire          compressDataVec_hitReq_12_222;
  assign compressDataVec_hitReq_12_222 = _GEN_997;
  wire          _GEN_998 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h1E;
  wire          compressDataVec_hitReq_13_30;
  assign compressDataVec_hitReq_13_30 = _GEN_998;
  wire          compressDataVec_hitReq_13_158;
  assign compressDataVec_hitReq_13_158 = _GEN_998;
  wire          compressDataVec_hitReq_13_222;
  assign compressDataVec_hitReq_13_222 = _GEN_998;
  wire          _GEN_999 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h1E;
  wire          compressDataVec_hitReq_14_30;
  assign compressDataVec_hitReq_14_30 = _GEN_999;
  wire          compressDataVec_hitReq_14_158;
  assign compressDataVec_hitReq_14_158 = _GEN_999;
  wire          compressDataVec_hitReq_14_222;
  assign compressDataVec_hitReq_14_222 = _GEN_999;
  wire          _GEN_1000 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h1E;
  wire          compressDataVec_hitReq_15_30;
  assign compressDataVec_hitReq_15_30 = _GEN_1000;
  wire          compressDataVec_hitReq_15_158;
  assign compressDataVec_hitReq_15_158 = _GEN_1000;
  wire          compressDataVec_hitReq_15_222;
  assign compressDataVec_hitReq_15_222 = _GEN_1000;
  wire          _GEN_1001 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h1E;
  wire          compressDataVec_hitReq_16_30;
  assign compressDataVec_hitReq_16_30 = _GEN_1001;
  wire          compressDataVec_hitReq_16_158;
  assign compressDataVec_hitReq_16_158 = _GEN_1001;
  wire          _GEN_1002 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h1E;
  wire          compressDataVec_hitReq_17_30;
  assign compressDataVec_hitReq_17_30 = _GEN_1002;
  wire          compressDataVec_hitReq_17_158;
  assign compressDataVec_hitReq_17_158 = _GEN_1002;
  wire          _GEN_1003 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h1E;
  wire          compressDataVec_hitReq_18_30;
  assign compressDataVec_hitReq_18_30 = _GEN_1003;
  wire          compressDataVec_hitReq_18_158;
  assign compressDataVec_hitReq_18_158 = _GEN_1003;
  wire          _GEN_1004 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h1E;
  wire          compressDataVec_hitReq_19_30;
  assign compressDataVec_hitReq_19_30 = _GEN_1004;
  wire          compressDataVec_hitReq_19_158;
  assign compressDataVec_hitReq_19_158 = _GEN_1004;
  wire          _GEN_1005 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h1E;
  wire          compressDataVec_hitReq_20_30;
  assign compressDataVec_hitReq_20_30 = _GEN_1005;
  wire          compressDataVec_hitReq_20_158;
  assign compressDataVec_hitReq_20_158 = _GEN_1005;
  wire          _GEN_1006 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h1E;
  wire          compressDataVec_hitReq_21_30;
  assign compressDataVec_hitReq_21_30 = _GEN_1006;
  wire          compressDataVec_hitReq_21_158;
  assign compressDataVec_hitReq_21_158 = _GEN_1006;
  wire          _GEN_1007 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h1E;
  wire          compressDataVec_hitReq_22_30;
  assign compressDataVec_hitReq_22_30 = _GEN_1007;
  wire          compressDataVec_hitReq_22_158;
  assign compressDataVec_hitReq_22_158 = _GEN_1007;
  wire          _GEN_1008 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h1E;
  wire          compressDataVec_hitReq_23_30;
  assign compressDataVec_hitReq_23_30 = _GEN_1008;
  wire          compressDataVec_hitReq_23_158;
  assign compressDataVec_hitReq_23_158 = _GEN_1008;
  wire          _GEN_1009 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h1E;
  wire          compressDataVec_hitReq_24_30;
  assign compressDataVec_hitReq_24_30 = _GEN_1009;
  wire          compressDataVec_hitReq_24_158;
  assign compressDataVec_hitReq_24_158 = _GEN_1009;
  wire          _GEN_1010 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h1E;
  wire          compressDataVec_hitReq_25_30;
  assign compressDataVec_hitReq_25_30 = _GEN_1010;
  wire          compressDataVec_hitReq_25_158;
  assign compressDataVec_hitReq_25_158 = _GEN_1010;
  wire          _GEN_1011 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h1E;
  wire          compressDataVec_hitReq_26_30;
  assign compressDataVec_hitReq_26_30 = _GEN_1011;
  wire          compressDataVec_hitReq_26_158;
  assign compressDataVec_hitReq_26_158 = _GEN_1011;
  wire          _GEN_1012 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h1E;
  wire          compressDataVec_hitReq_27_30;
  assign compressDataVec_hitReq_27_30 = _GEN_1012;
  wire          compressDataVec_hitReq_27_158;
  assign compressDataVec_hitReq_27_158 = _GEN_1012;
  wire          _GEN_1013 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h1E;
  wire          compressDataVec_hitReq_28_30;
  assign compressDataVec_hitReq_28_30 = _GEN_1013;
  wire          compressDataVec_hitReq_28_158;
  assign compressDataVec_hitReq_28_158 = _GEN_1013;
  wire          _GEN_1014 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h1E;
  wire          compressDataVec_hitReq_29_30;
  assign compressDataVec_hitReq_29_30 = _GEN_1014;
  wire          compressDataVec_hitReq_29_158;
  assign compressDataVec_hitReq_29_158 = _GEN_1014;
  wire          _GEN_1015 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h1E;
  wire          compressDataVec_hitReq_30_30;
  assign compressDataVec_hitReq_30_30 = _GEN_1015;
  wire          compressDataVec_hitReq_30_158;
  assign compressDataVec_hitReq_30_158 = _GEN_1015;
  wire          _GEN_1016 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h1E;
  wire          compressDataVec_hitReq_31_30;
  assign compressDataVec_hitReq_31_30 = _GEN_1016;
  wire          compressDataVec_hitReq_31_158;
  assign compressDataVec_hitReq_31_158 = _GEN_1016;
  wire          compressDataVec_hitReq_32_30 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h1E;
  wire          compressDataVec_hitReq_33_30 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h1E;
  wire          compressDataVec_hitReq_34_30 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h1E;
  wire          compressDataVec_hitReq_35_30 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h1E;
  wire          compressDataVec_hitReq_36_30 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h1E;
  wire          compressDataVec_hitReq_37_30 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h1E;
  wire          compressDataVec_hitReq_38_30 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h1E;
  wire          compressDataVec_hitReq_39_30 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h1E;
  wire          compressDataVec_hitReq_40_30 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h1E;
  wire          compressDataVec_hitReq_41_30 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h1E;
  wire          compressDataVec_hitReq_42_30 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h1E;
  wire          compressDataVec_hitReq_43_30 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h1E;
  wire          compressDataVec_hitReq_44_30 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h1E;
  wire          compressDataVec_hitReq_45_30 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h1E;
  wire          compressDataVec_hitReq_46_30 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h1E;
  wire          compressDataVec_hitReq_47_30 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h1E;
  wire          compressDataVec_hitReq_48_30 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h1E;
  wire          compressDataVec_hitReq_49_30 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h1E;
  wire          compressDataVec_hitReq_50_30 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h1E;
  wire          compressDataVec_hitReq_51_30 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h1E;
  wire          compressDataVec_hitReq_52_30 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h1E;
  wire          compressDataVec_hitReq_53_30 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h1E;
  wire          compressDataVec_hitReq_54_30 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h1E;
  wire          compressDataVec_hitReq_55_30 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h1E;
  wire          compressDataVec_hitReq_56_30 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h1E;
  wire          compressDataVec_hitReq_57_30 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h1E;
  wire          compressDataVec_hitReq_58_30 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h1E;
  wire          compressDataVec_hitReq_59_30 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h1E;
  wire          compressDataVec_hitReq_60_30 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h1E;
  wire          compressDataVec_hitReq_61_30 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h1E;
  wire          compressDataVec_hitReq_62_30 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h1E;
  wire          compressDataVec_hitReq_63_30 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h1E;
  wire [7:0]    compressDataVec_selectReqData_30 =
    (compressDataVec_hitReq_0_30 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_30 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_30 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_30 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_30 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_30 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_30 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_30 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_30 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_30 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_30 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_30 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_30 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_30 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_30 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_30 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_30 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_30 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_30 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_30 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_30 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_30 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_30 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_30 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_30 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_30 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_30 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_30 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_30 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_30 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_30 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_30 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_30 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_30 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_30 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_30 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_30 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_30 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_30 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_30 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_30 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_30 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_30 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_30 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_30 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_30 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_30 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_30 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_30 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_30 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_30 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_30 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_30 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_30 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_30 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_30 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_30 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_30 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_30 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_30 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_30 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_30 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_30 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_30 ? source2Pipe[511:504] : 8'h0);
  wire          _GEN_1017 = tailCount > 6'h1E;
  wire          compressDataVec_useTail_30;
  assign compressDataVec_useTail_30 = _GEN_1017;
  wire          compressDataVec_useTail_94;
  assign compressDataVec_useTail_94 = _GEN_1017;
  wire          _GEN_1018 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h1F;
  wire          compressDataVec_hitReq_0_31;
  assign compressDataVec_hitReq_0_31 = _GEN_1018;
  wire          compressDataVec_hitReq_0_159;
  assign compressDataVec_hitReq_0_159 = _GEN_1018;
  wire          compressDataVec_hitReq_0_223;
  assign compressDataVec_hitReq_0_223 = _GEN_1018;
  wire          _GEN_1019 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h1F;
  wire          compressDataVec_hitReq_1_31;
  assign compressDataVec_hitReq_1_31 = _GEN_1019;
  wire          compressDataVec_hitReq_1_159;
  assign compressDataVec_hitReq_1_159 = _GEN_1019;
  wire          compressDataVec_hitReq_1_223;
  assign compressDataVec_hitReq_1_223 = _GEN_1019;
  wire          _GEN_1020 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h1F;
  wire          compressDataVec_hitReq_2_31;
  assign compressDataVec_hitReq_2_31 = _GEN_1020;
  wire          compressDataVec_hitReq_2_159;
  assign compressDataVec_hitReq_2_159 = _GEN_1020;
  wire          compressDataVec_hitReq_2_223;
  assign compressDataVec_hitReq_2_223 = _GEN_1020;
  wire          _GEN_1021 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h1F;
  wire          compressDataVec_hitReq_3_31;
  assign compressDataVec_hitReq_3_31 = _GEN_1021;
  wire          compressDataVec_hitReq_3_159;
  assign compressDataVec_hitReq_3_159 = _GEN_1021;
  wire          compressDataVec_hitReq_3_223;
  assign compressDataVec_hitReq_3_223 = _GEN_1021;
  wire          _GEN_1022 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h1F;
  wire          compressDataVec_hitReq_4_31;
  assign compressDataVec_hitReq_4_31 = _GEN_1022;
  wire          compressDataVec_hitReq_4_159;
  assign compressDataVec_hitReq_4_159 = _GEN_1022;
  wire          compressDataVec_hitReq_4_223;
  assign compressDataVec_hitReq_4_223 = _GEN_1022;
  wire          _GEN_1023 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h1F;
  wire          compressDataVec_hitReq_5_31;
  assign compressDataVec_hitReq_5_31 = _GEN_1023;
  wire          compressDataVec_hitReq_5_159;
  assign compressDataVec_hitReq_5_159 = _GEN_1023;
  wire          compressDataVec_hitReq_5_223;
  assign compressDataVec_hitReq_5_223 = _GEN_1023;
  wire          _GEN_1024 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h1F;
  wire          compressDataVec_hitReq_6_31;
  assign compressDataVec_hitReq_6_31 = _GEN_1024;
  wire          compressDataVec_hitReq_6_159;
  assign compressDataVec_hitReq_6_159 = _GEN_1024;
  wire          compressDataVec_hitReq_6_223;
  assign compressDataVec_hitReq_6_223 = _GEN_1024;
  wire          _GEN_1025 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h1F;
  wire          compressDataVec_hitReq_7_31;
  assign compressDataVec_hitReq_7_31 = _GEN_1025;
  wire          compressDataVec_hitReq_7_159;
  assign compressDataVec_hitReq_7_159 = _GEN_1025;
  wire          compressDataVec_hitReq_7_223;
  assign compressDataVec_hitReq_7_223 = _GEN_1025;
  wire          _GEN_1026 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h1F;
  wire          compressDataVec_hitReq_8_31;
  assign compressDataVec_hitReq_8_31 = _GEN_1026;
  wire          compressDataVec_hitReq_8_159;
  assign compressDataVec_hitReq_8_159 = _GEN_1026;
  wire          compressDataVec_hitReq_8_223;
  assign compressDataVec_hitReq_8_223 = _GEN_1026;
  wire          _GEN_1027 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h1F;
  wire          compressDataVec_hitReq_9_31;
  assign compressDataVec_hitReq_9_31 = _GEN_1027;
  wire          compressDataVec_hitReq_9_159;
  assign compressDataVec_hitReq_9_159 = _GEN_1027;
  wire          compressDataVec_hitReq_9_223;
  assign compressDataVec_hitReq_9_223 = _GEN_1027;
  wire          _GEN_1028 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h1F;
  wire          compressDataVec_hitReq_10_31;
  assign compressDataVec_hitReq_10_31 = _GEN_1028;
  wire          compressDataVec_hitReq_10_159;
  assign compressDataVec_hitReq_10_159 = _GEN_1028;
  wire          compressDataVec_hitReq_10_223;
  assign compressDataVec_hitReq_10_223 = _GEN_1028;
  wire          _GEN_1029 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h1F;
  wire          compressDataVec_hitReq_11_31;
  assign compressDataVec_hitReq_11_31 = _GEN_1029;
  wire          compressDataVec_hitReq_11_159;
  assign compressDataVec_hitReq_11_159 = _GEN_1029;
  wire          compressDataVec_hitReq_11_223;
  assign compressDataVec_hitReq_11_223 = _GEN_1029;
  wire          _GEN_1030 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h1F;
  wire          compressDataVec_hitReq_12_31;
  assign compressDataVec_hitReq_12_31 = _GEN_1030;
  wire          compressDataVec_hitReq_12_159;
  assign compressDataVec_hitReq_12_159 = _GEN_1030;
  wire          compressDataVec_hitReq_12_223;
  assign compressDataVec_hitReq_12_223 = _GEN_1030;
  wire          _GEN_1031 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h1F;
  wire          compressDataVec_hitReq_13_31;
  assign compressDataVec_hitReq_13_31 = _GEN_1031;
  wire          compressDataVec_hitReq_13_159;
  assign compressDataVec_hitReq_13_159 = _GEN_1031;
  wire          compressDataVec_hitReq_13_223;
  assign compressDataVec_hitReq_13_223 = _GEN_1031;
  wire          _GEN_1032 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h1F;
  wire          compressDataVec_hitReq_14_31;
  assign compressDataVec_hitReq_14_31 = _GEN_1032;
  wire          compressDataVec_hitReq_14_159;
  assign compressDataVec_hitReq_14_159 = _GEN_1032;
  wire          compressDataVec_hitReq_14_223;
  assign compressDataVec_hitReq_14_223 = _GEN_1032;
  wire          _GEN_1033 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h1F;
  wire          compressDataVec_hitReq_15_31;
  assign compressDataVec_hitReq_15_31 = _GEN_1033;
  wire          compressDataVec_hitReq_15_159;
  assign compressDataVec_hitReq_15_159 = _GEN_1033;
  wire          compressDataVec_hitReq_15_223;
  assign compressDataVec_hitReq_15_223 = _GEN_1033;
  wire          _GEN_1034 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h1F;
  wire          compressDataVec_hitReq_16_31;
  assign compressDataVec_hitReq_16_31 = _GEN_1034;
  wire          compressDataVec_hitReq_16_159;
  assign compressDataVec_hitReq_16_159 = _GEN_1034;
  wire          _GEN_1035 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h1F;
  wire          compressDataVec_hitReq_17_31;
  assign compressDataVec_hitReq_17_31 = _GEN_1035;
  wire          compressDataVec_hitReq_17_159;
  assign compressDataVec_hitReq_17_159 = _GEN_1035;
  wire          _GEN_1036 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h1F;
  wire          compressDataVec_hitReq_18_31;
  assign compressDataVec_hitReq_18_31 = _GEN_1036;
  wire          compressDataVec_hitReq_18_159;
  assign compressDataVec_hitReq_18_159 = _GEN_1036;
  wire          _GEN_1037 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h1F;
  wire          compressDataVec_hitReq_19_31;
  assign compressDataVec_hitReq_19_31 = _GEN_1037;
  wire          compressDataVec_hitReq_19_159;
  assign compressDataVec_hitReq_19_159 = _GEN_1037;
  wire          _GEN_1038 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h1F;
  wire          compressDataVec_hitReq_20_31;
  assign compressDataVec_hitReq_20_31 = _GEN_1038;
  wire          compressDataVec_hitReq_20_159;
  assign compressDataVec_hitReq_20_159 = _GEN_1038;
  wire          _GEN_1039 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h1F;
  wire          compressDataVec_hitReq_21_31;
  assign compressDataVec_hitReq_21_31 = _GEN_1039;
  wire          compressDataVec_hitReq_21_159;
  assign compressDataVec_hitReq_21_159 = _GEN_1039;
  wire          _GEN_1040 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h1F;
  wire          compressDataVec_hitReq_22_31;
  assign compressDataVec_hitReq_22_31 = _GEN_1040;
  wire          compressDataVec_hitReq_22_159;
  assign compressDataVec_hitReq_22_159 = _GEN_1040;
  wire          _GEN_1041 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h1F;
  wire          compressDataVec_hitReq_23_31;
  assign compressDataVec_hitReq_23_31 = _GEN_1041;
  wire          compressDataVec_hitReq_23_159;
  assign compressDataVec_hitReq_23_159 = _GEN_1041;
  wire          _GEN_1042 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h1F;
  wire          compressDataVec_hitReq_24_31;
  assign compressDataVec_hitReq_24_31 = _GEN_1042;
  wire          compressDataVec_hitReq_24_159;
  assign compressDataVec_hitReq_24_159 = _GEN_1042;
  wire          _GEN_1043 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h1F;
  wire          compressDataVec_hitReq_25_31;
  assign compressDataVec_hitReq_25_31 = _GEN_1043;
  wire          compressDataVec_hitReq_25_159;
  assign compressDataVec_hitReq_25_159 = _GEN_1043;
  wire          _GEN_1044 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h1F;
  wire          compressDataVec_hitReq_26_31;
  assign compressDataVec_hitReq_26_31 = _GEN_1044;
  wire          compressDataVec_hitReq_26_159;
  assign compressDataVec_hitReq_26_159 = _GEN_1044;
  wire          _GEN_1045 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h1F;
  wire          compressDataVec_hitReq_27_31;
  assign compressDataVec_hitReq_27_31 = _GEN_1045;
  wire          compressDataVec_hitReq_27_159;
  assign compressDataVec_hitReq_27_159 = _GEN_1045;
  wire          _GEN_1046 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h1F;
  wire          compressDataVec_hitReq_28_31;
  assign compressDataVec_hitReq_28_31 = _GEN_1046;
  wire          compressDataVec_hitReq_28_159;
  assign compressDataVec_hitReq_28_159 = _GEN_1046;
  wire          _GEN_1047 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h1F;
  wire          compressDataVec_hitReq_29_31;
  assign compressDataVec_hitReq_29_31 = _GEN_1047;
  wire          compressDataVec_hitReq_29_159;
  assign compressDataVec_hitReq_29_159 = _GEN_1047;
  wire          _GEN_1048 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h1F;
  wire          compressDataVec_hitReq_30_31;
  assign compressDataVec_hitReq_30_31 = _GEN_1048;
  wire          compressDataVec_hitReq_30_159;
  assign compressDataVec_hitReq_30_159 = _GEN_1048;
  wire          _GEN_1049 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h1F;
  wire          compressDataVec_hitReq_31_31;
  assign compressDataVec_hitReq_31_31 = _GEN_1049;
  wire          compressDataVec_hitReq_31_159;
  assign compressDataVec_hitReq_31_159 = _GEN_1049;
  wire          compressDataVec_hitReq_32_31 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h1F;
  wire          compressDataVec_hitReq_33_31 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h1F;
  wire          compressDataVec_hitReq_34_31 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h1F;
  wire          compressDataVec_hitReq_35_31 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h1F;
  wire          compressDataVec_hitReq_36_31 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h1F;
  wire          compressDataVec_hitReq_37_31 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h1F;
  wire          compressDataVec_hitReq_38_31 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h1F;
  wire          compressDataVec_hitReq_39_31 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h1F;
  wire          compressDataVec_hitReq_40_31 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h1F;
  wire          compressDataVec_hitReq_41_31 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h1F;
  wire          compressDataVec_hitReq_42_31 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h1F;
  wire          compressDataVec_hitReq_43_31 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h1F;
  wire          compressDataVec_hitReq_44_31 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h1F;
  wire          compressDataVec_hitReq_45_31 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h1F;
  wire          compressDataVec_hitReq_46_31 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h1F;
  wire          compressDataVec_hitReq_47_31 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h1F;
  wire          compressDataVec_hitReq_48_31 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h1F;
  wire          compressDataVec_hitReq_49_31 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h1F;
  wire          compressDataVec_hitReq_50_31 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h1F;
  wire          compressDataVec_hitReq_51_31 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h1F;
  wire          compressDataVec_hitReq_52_31 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h1F;
  wire          compressDataVec_hitReq_53_31 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h1F;
  wire          compressDataVec_hitReq_54_31 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h1F;
  wire          compressDataVec_hitReq_55_31 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h1F;
  wire          compressDataVec_hitReq_56_31 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h1F;
  wire          compressDataVec_hitReq_57_31 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h1F;
  wire          compressDataVec_hitReq_58_31 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h1F;
  wire          compressDataVec_hitReq_59_31 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h1F;
  wire          compressDataVec_hitReq_60_31 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h1F;
  wire          compressDataVec_hitReq_61_31 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h1F;
  wire          compressDataVec_hitReq_62_31 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h1F;
  wire          compressDataVec_hitReq_63_31 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h1F;
  wire [7:0]    compressDataVec_selectReqData_31 =
    (compressDataVec_hitReq_0_31 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_31 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_31 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_31 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_31 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_31 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_31 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_31 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_31 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_31 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_31 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_31 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_31 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_31 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_31 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_31 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_31 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_31 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_31 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_31 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_31 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_31 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_31 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_31 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_31 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_31 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_31 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_31 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_31 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_31 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_31 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_31 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_31 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_31 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_31 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_31 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_31 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_31 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_31 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_31 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_31 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_31 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_31 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_31 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_31 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_31 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_31 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_31 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_31 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_31 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_31 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_31 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_31 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_31 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_31 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_31 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_31 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_31 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_31 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_31 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_31 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_31 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_31 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_31 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_31 = tailCount[5];
  wire          compressDataVec_useTail_95 = tailCount[5];
  wire          _GEN_1050 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h20;
  wire          compressDataVec_hitReq_0_32;
  assign compressDataVec_hitReq_0_32 = _GEN_1050;
  wire          compressDataVec_hitReq_0_160;
  assign compressDataVec_hitReq_0_160 = _GEN_1050;
  wire          _GEN_1051 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h20;
  wire          compressDataVec_hitReq_1_32;
  assign compressDataVec_hitReq_1_32 = _GEN_1051;
  wire          compressDataVec_hitReq_1_160;
  assign compressDataVec_hitReq_1_160 = _GEN_1051;
  wire          _GEN_1052 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h20;
  wire          compressDataVec_hitReq_2_32;
  assign compressDataVec_hitReq_2_32 = _GEN_1052;
  wire          compressDataVec_hitReq_2_160;
  assign compressDataVec_hitReq_2_160 = _GEN_1052;
  wire          _GEN_1053 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h20;
  wire          compressDataVec_hitReq_3_32;
  assign compressDataVec_hitReq_3_32 = _GEN_1053;
  wire          compressDataVec_hitReq_3_160;
  assign compressDataVec_hitReq_3_160 = _GEN_1053;
  wire          _GEN_1054 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h20;
  wire          compressDataVec_hitReq_4_32;
  assign compressDataVec_hitReq_4_32 = _GEN_1054;
  wire          compressDataVec_hitReq_4_160;
  assign compressDataVec_hitReq_4_160 = _GEN_1054;
  wire          _GEN_1055 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h20;
  wire          compressDataVec_hitReq_5_32;
  assign compressDataVec_hitReq_5_32 = _GEN_1055;
  wire          compressDataVec_hitReq_5_160;
  assign compressDataVec_hitReq_5_160 = _GEN_1055;
  wire          _GEN_1056 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h20;
  wire          compressDataVec_hitReq_6_32;
  assign compressDataVec_hitReq_6_32 = _GEN_1056;
  wire          compressDataVec_hitReq_6_160;
  assign compressDataVec_hitReq_6_160 = _GEN_1056;
  wire          _GEN_1057 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h20;
  wire          compressDataVec_hitReq_7_32;
  assign compressDataVec_hitReq_7_32 = _GEN_1057;
  wire          compressDataVec_hitReq_7_160;
  assign compressDataVec_hitReq_7_160 = _GEN_1057;
  wire          _GEN_1058 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h20;
  wire          compressDataVec_hitReq_8_32;
  assign compressDataVec_hitReq_8_32 = _GEN_1058;
  wire          compressDataVec_hitReq_8_160;
  assign compressDataVec_hitReq_8_160 = _GEN_1058;
  wire          _GEN_1059 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h20;
  wire          compressDataVec_hitReq_9_32;
  assign compressDataVec_hitReq_9_32 = _GEN_1059;
  wire          compressDataVec_hitReq_9_160;
  assign compressDataVec_hitReq_9_160 = _GEN_1059;
  wire          _GEN_1060 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h20;
  wire          compressDataVec_hitReq_10_32;
  assign compressDataVec_hitReq_10_32 = _GEN_1060;
  wire          compressDataVec_hitReq_10_160;
  assign compressDataVec_hitReq_10_160 = _GEN_1060;
  wire          _GEN_1061 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h20;
  wire          compressDataVec_hitReq_11_32;
  assign compressDataVec_hitReq_11_32 = _GEN_1061;
  wire          compressDataVec_hitReq_11_160;
  assign compressDataVec_hitReq_11_160 = _GEN_1061;
  wire          _GEN_1062 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h20;
  wire          compressDataVec_hitReq_12_32;
  assign compressDataVec_hitReq_12_32 = _GEN_1062;
  wire          compressDataVec_hitReq_12_160;
  assign compressDataVec_hitReq_12_160 = _GEN_1062;
  wire          _GEN_1063 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h20;
  wire          compressDataVec_hitReq_13_32;
  assign compressDataVec_hitReq_13_32 = _GEN_1063;
  wire          compressDataVec_hitReq_13_160;
  assign compressDataVec_hitReq_13_160 = _GEN_1063;
  wire          _GEN_1064 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h20;
  wire          compressDataVec_hitReq_14_32;
  assign compressDataVec_hitReq_14_32 = _GEN_1064;
  wire          compressDataVec_hitReq_14_160;
  assign compressDataVec_hitReq_14_160 = _GEN_1064;
  wire          _GEN_1065 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h20;
  wire          compressDataVec_hitReq_15_32;
  assign compressDataVec_hitReq_15_32 = _GEN_1065;
  wire          compressDataVec_hitReq_15_160;
  assign compressDataVec_hitReq_15_160 = _GEN_1065;
  wire          _GEN_1066 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h20;
  wire          compressDataVec_hitReq_16_32;
  assign compressDataVec_hitReq_16_32 = _GEN_1066;
  wire          compressDataVec_hitReq_16_160;
  assign compressDataVec_hitReq_16_160 = _GEN_1066;
  wire          _GEN_1067 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h20;
  wire          compressDataVec_hitReq_17_32;
  assign compressDataVec_hitReq_17_32 = _GEN_1067;
  wire          compressDataVec_hitReq_17_160;
  assign compressDataVec_hitReq_17_160 = _GEN_1067;
  wire          _GEN_1068 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h20;
  wire          compressDataVec_hitReq_18_32;
  assign compressDataVec_hitReq_18_32 = _GEN_1068;
  wire          compressDataVec_hitReq_18_160;
  assign compressDataVec_hitReq_18_160 = _GEN_1068;
  wire          _GEN_1069 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h20;
  wire          compressDataVec_hitReq_19_32;
  assign compressDataVec_hitReq_19_32 = _GEN_1069;
  wire          compressDataVec_hitReq_19_160;
  assign compressDataVec_hitReq_19_160 = _GEN_1069;
  wire          _GEN_1070 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h20;
  wire          compressDataVec_hitReq_20_32;
  assign compressDataVec_hitReq_20_32 = _GEN_1070;
  wire          compressDataVec_hitReq_20_160;
  assign compressDataVec_hitReq_20_160 = _GEN_1070;
  wire          _GEN_1071 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h20;
  wire          compressDataVec_hitReq_21_32;
  assign compressDataVec_hitReq_21_32 = _GEN_1071;
  wire          compressDataVec_hitReq_21_160;
  assign compressDataVec_hitReq_21_160 = _GEN_1071;
  wire          _GEN_1072 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h20;
  wire          compressDataVec_hitReq_22_32;
  assign compressDataVec_hitReq_22_32 = _GEN_1072;
  wire          compressDataVec_hitReq_22_160;
  assign compressDataVec_hitReq_22_160 = _GEN_1072;
  wire          _GEN_1073 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h20;
  wire          compressDataVec_hitReq_23_32;
  assign compressDataVec_hitReq_23_32 = _GEN_1073;
  wire          compressDataVec_hitReq_23_160;
  assign compressDataVec_hitReq_23_160 = _GEN_1073;
  wire          _GEN_1074 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h20;
  wire          compressDataVec_hitReq_24_32;
  assign compressDataVec_hitReq_24_32 = _GEN_1074;
  wire          compressDataVec_hitReq_24_160;
  assign compressDataVec_hitReq_24_160 = _GEN_1074;
  wire          _GEN_1075 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h20;
  wire          compressDataVec_hitReq_25_32;
  assign compressDataVec_hitReq_25_32 = _GEN_1075;
  wire          compressDataVec_hitReq_25_160;
  assign compressDataVec_hitReq_25_160 = _GEN_1075;
  wire          _GEN_1076 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h20;
  wire          compressDataVec_hitReq_26_32;
  assign compressDataVec_hitReq_26_32 = _GEN_1076;
  wire          compressDataVec_hitReq_26_160;
  assign compressDataVec_hitReq_26_160 = _GEN_1076;
  wire          _GEN_1077 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h20;
  wire          compressDataVec_hitReq_27_32;
  assign compressDataVec_hitReq_27_32 = _GEN_1077;
  wire          compressDataVec_hitReq_27_160;
  assign compressDataVec_hitReq_27_160 = _GEN_1077;
  wire          _GEN_1078 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h20;
  wire          compressDataVec_hitReq_28_32;
  assign compressDataVec_hitReq_28_32 = _GEN_1078;
  wire          compressDataVec_hitReq_28_160;
  assign compressDataVec_hitReq_28_160 = _GEN_1078;
  wire          _GEN_1079 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h20;
  wire          compressDataVec_hitReq_29_32;
  assign compressDataVec_hitReq_29_32 = _GEN_1079;
  wire          compressDataVec_hitReq_29_160;
  assign compressDataVec_hitReq_29_160 = _GEN_1079;
  wire          _GEN_1080 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h20;
  wire          compressDataVec_hitReq_30_32;
  assign compressDataVec_hitReq_30_32 = _GEN_1080;
  wire          compressDataVec_hitReq_30_160;
  assign compressDataVec_hitReq_30_160 = _GEN_1080;
  wire          _GEN_1081 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h20;
  wire          compressDataVec_hitReq_31_32;
  assign compressDataVec_hitReq_31_32 = _GEN_1081;
  wire          compressDataVec_hitReq_31_160;
  assign compressDataVec_hitReq_31_160 = _GEN_1081;
  wire          compressDataVec_hitReq_32_32 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h20;
  wire          compressDataVec_hitReq_33_32 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h20;
  wire          compressDataVec_hitReq_34_32 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h20;
  wire          compressDataVec_hitReq_35_32 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h20;
  wire          compressDataVec_hitReq_36_32 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h20;
  wire          compressDataVec_hitReq_37_32 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h20;
  wire          compressDataVec_hitReq_38_32 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h20;
  wire          compressDataVec_hitReq_39_32 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h20;
  wire          compressDataVec_hitReq_40_32 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h20;
  wire          compressDataVec_hitReq_41_32 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h20;
  wire          compressDataVec_hitReq_42_32 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h20;
  wire          compressDataVec_hitReq_43_32 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h20;
  wire          compressDataVec_hitReq_44_32 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h20;
  wire          compressDataVec_hitReq_45_32 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h20;
  wire          compressDataVec_hitReq_46_32 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h20;
  wire          compressDataVec_hitReq_47_32 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h20;
  wire          compressDataVec_hitReq_48_32 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h20;
  wire          compressDataVec_hitReq_49_32 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h20;
  wire          compressDataVec_hitReq_50_32 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h20;
  wire          compressDataVec_hitReq_51_32 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h20;
  wire          compressDataVec_hitReq_52_32 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h20;
  wire          compressDataVec_hitReq_53_32 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h20;
  wire          compressDataVec_hitReq_54_32 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h20;
  wire          compressDataVec_hitReq_55_32 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h20;
  wire          compressDataVec_hitReq_56_32 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h20;
  wire          compressDataVec_hitReq_57_32 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h20;
  wire          compressDataVec_hitReq_58_32 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h20;
  wire          compressDataVec_hitReq_59_32 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h20;
  wire          compressDataVec_hitReq_60_32 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h20;
  wire          compressDataVec_hitReq_61_32 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h20;
  wire          compressDataVec_hitReq_62_32 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h20;
  wire          compressDataVec_hitReq_63_32 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h20;
  wire [7:0]    compressDataVec_selectReqData_32 =
    (compressDataVec_hitReq_0_32 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_32 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_32 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_32 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_32 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_32 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_32 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_32 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_32 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_32 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_32 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_32 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_32 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_32 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_32 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_32 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_32 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_32 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_32 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_32 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_32 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_32 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_32 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_32 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_32 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_32 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_32 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_32 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_32 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_32 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_32 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_32 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_32 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_32 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_32 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_32 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_32 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_32 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_32 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_32 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_32 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_32 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_32 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_32 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_32 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_32 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_32 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_32 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_32 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_32 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_32 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_32 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_32 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_32 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_32 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_32 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_32 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_32 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_32 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_32 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_32 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_32 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_32 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_32 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_32 = tailCount > 6'h20;
  wire          _GEN_1082 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h21;
  wire          compressDataVec_hitReq_0_33;
  assign compressDataVec_hitReq_0_33 = _GEN_1082;
  wire          compressDataVec_hitReq_0_161;
  assign compressDataVec_hitReq_0_161 = _GEN_1082;
  wire          _GEN_1083 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h21;
  wire          compressDataVec_hitReq_1_33;
  assign compressDataVec_hitReq_1_33 = _GEN_1083;
  wire          compressDataVec_hitReq_1_161;
  assign compressDataVec_hitReq_1_161 = _GEN_1083;
  wire          _GEN_1084 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h21;
  wire          compressDataVec_hitReq_2_33;
  assign compressDataVec_hitReq_2_33 = _GEN_1084;
  wire          compressDataVec_hitReq_2_161;
  assign compressDataVec_hitReq_2_161 = _GEN_1084;
  wire          _GEN_1085 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h21;
  wire          compressDataVec_hitReq_3_33;
  assign compressDataVec_hitReq_3_33 = _GEN_1085;
  wire          compressDataVec_hitReq_3_161;
  assign compressDataVec_hitReq_3_161 = _GEN_1085;
  wire          _GEN_1086 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h21;
  wire          compressDataVec_hitReq_4_33;
  assign compressDataVec_hitReq_4_33 = _GEN_1086;
  wire          compressDataVec_hitReq_4_161;
  assign compressDataVec_hitReq_4_161 = _GEN_1086;
  wire          _GEN_1087 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h21;
  wire          compressDataVec_hitReq_5_33;
  assign compressDataVec_hitReq_5_33 = _GEN_1087;
  wire          compressDataVec_hitReq_5_161;
  assign compressDataVec_hitReq_5_161 = _GEN_1087;
  wire          _GEN_1088 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h21;
  wire          compressDataVec_hitReq_6_33;
  assign compressDataVec_hitReq_6_33 = _GEN_1088;
  wire          compressDataVec_hitReq_6_161;
  assign compressDataVec_hitReq_6_161 = _GEN_1088;
  wire          _GEN_1089 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h21;
  wire          compressDataVec_hitReq_7_33;
  assign compressDataVec_hitReq_7_33 = _GEN_1089;
  wire          compressDataVec_hitReq_7_161;
  assign compressDataVec_hitReq_7_161 = _GEN_1089;
  wire          _GEN_1090 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h21;
  wire          compressDataVec_hitReq_8_33;
  assign compressDataVec_hitReq_8_33 = _GEN_1090;
  wire          compressDataVec_hitReq_8_161;
  assign compressDataVec_hitReq_8_161 = _GEN_1090;
  wire          _GEN_1091 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h21;
  wire          compressDataVec_hitReq_9_33;
  assign compressDataVec_hitReq_9_33 = _GEN_1091;
  wire          compressDataVec_hitReq_9_161;
  assign compressDataVec_hitReq_9_161 = _GEN_1091;
  wire          _GEN_1092 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h21;
  wire          compressDataVec_hitReq_10_33;
  assign compressDataVec_hitReq_10_33 = _GEN_1092;
  wire          compressDataVec_hitReq_10_161;
  assign compressDataVec_hitReq_10_161 = _GEN_1092;
  wire          _GEN_1093 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h21;
  wire          compressDataVec_hitReq_11_33;
  assign compressDataVec_hitReq_11_33 = _GEN_1093;
  wire          compressDataVec_hitReq_11_161;
  assign compressDataVec_hitReq_11_161 = _GEN_1093;
  wire          _GEN_1094 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h21;
  wire          compressDataVec_hitReq_12_33;
  assign compressDataVec_hitReq_12_33 = _GEN_1094;
  wire          compressDataVec_hitReq_12_161;
  assign compressDataVec_hitReq_12_161 = _GEN_1094;
  wire          _GEN_1095 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h21;
  wire          compressDataVec_hitReq_13_33;
  assign compressDataVec_hitReq_13_33 = _GEN_1095;
  wire          compressDataVec_hitReq_13_161;
  assign compressDataVec_hitReq_13_161 = _GEN_1095;
  wire          _GEN_1096 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h21;
  wire          compressDataVec_hitReq_14_33;
  assign compressDataVec_hitReq_14_33 = _GEN_1096;
  wire          compressDataVec_hitReq_14_161;
  assign compressDataVec_hitReq_14_161 = _GEN_1096;
  wire          _GEN_1097 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h21;
  wire          compressDataVec_hitReq_15_33;
  assign compressDataVec_hitReq_15_33 = _GEN_1097;
  wire          compressDataVec_hitReq_15_161;
  assign compressDataVec_hitReq_15_161 = _GEN_1097;
  wire          _GEN_1098 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h21;
  wire          compressDataVec_hitReq_16_33;
  assign compressDataVec_hitReq_16_33 = _GEN_1098;
  wire          compressDataVec_hitReq_16_161;
  assign compressDataVec_hitReq_16_161 = _GEN_1098;
  wire          _GEN_1099 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h21;
  wire          compressDataVec_hitReq_17_33;
  assign compressDataVec_hitReq_17_33 = _GEN_1099;
  wire          compressDataVec_hitReq_17_161;
  assign compressDataVec_hitReq_17_161 = _GEN_1099;
  wire          _GEN_1100 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h21;
  wire          compressDataVec_hitReq_18_33;
  assign compressDataVec_hitReq_18_33 = _GEN_1100;
  wire          compressDataVec_hitReq_18_161;
  assign compressDataVec_hitReq_18_161 = _GEN_1100;
  wire          _GEN_1101 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h21;
  wire          compressDataVec_hitReq_19_33;
  assign compressDataVec_hitReq_19_33 = _GEN_1101;
  wire          compressDataVec_hitReq_19_161;
  assign compressDataVec_hitReq_19_161 = _GEN_1101;
  wire          _GEN_1102 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h21;
  wire          compressDataVec_hitReq_20_33;
  assign compressDataVec_hitReq_20_33 = _GEN_1102;
  wire          compressDataVec_hitReq_20_161;
  assign compressDataVec_hitReq_20_161 = _GEN_1102;
  wire          _GEN_1103 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h21;
  wire          compressDataVec_hitReq_21_33;
  assign compressDataVec_hitReq_21_33 = _GEN_1103;
  wire          compressDataVec_hitReq_21_161;
  assign compressDataVec_hitReq_21_161 = _GEN_1103;
  wire          _GEN_1104 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h21;
  wire          compressDataVec_hitReq_22_33;
  assign compressDataVec_hitReq_22_33 = _GEN_1104;
  wire          compressDataVec_hitReq_22_161;
  assign compressDataVec_hitReq_22_161 = _GEN_1104;
  wire          _GEN_1105 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h21;
  wire          compressDataVec_hitReq_23_33;
  assign compressDataVec_hitReq_23_33 = _GEN_1105;
  wire          compressDataVec_hitReq_23_161;
  assign compressDataVec_hitReq_23_161 = _GEN_1105;
  wire          _GEN_1106 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h21;
  wire          compressDataVec_hitReq_24_33;
  assign compressDataVec_hitReq_24_33 = _GEN_1106;
  wire          compressDataVec_hitReq_24_161;
  assign compressDataVec_hitReq_24_161 = _GEN_1106;
  wire          _GEN_1107 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h21;
  wire          compressDataVec_hitReq_25_33;
  assign compressDataVec_hitReq_25_33 = _GEN_1107;
  wire          compressDataVec_hitReq_25_161;
  assign compressDataVec_hitReq_25_161 = _GEN_1107;
  wire          _GEN_1108 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h21;
  wire          compressDataVec_hitReq_26_33;
  assign compressDataVec_hitReq_26_33 = _GEN_1108;
  wire          compressDataVec_hitReq_26_161;
  assign compressDataVec_hitReq_26_161 = _GEN_1108;
  wire          _GEN_1109 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h21;
  wire          compressDataVec_hitReq_27_33;
  assign compressDataVec_hitReq_27_33 = _GEN_1109;
  wire          compressDataVec_hitReq_27_161;
  assign compressDataVec_hitReq_27_161 = _GEN_1109;
  wire          _GEN_1110 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h21;
  wire          compressDataVec_hitReq_28_33;
  assign compressDataVec_hitReq_28_33 = _GEN_1110;
  wire          compressDataVec_hitReq_28_161;
  assign compressDataVec_hitReq_28_161 = _GEN_1110;
  wire          _GEN_1111 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h21;
  wire          compressDataVec_hitReq_29_33;
  assign compressDataVec_hitReq_29_33 = _GEN_1111;
  wire          compressDataVec_hitReq_29_161;
  assign compressDataVec_hitReq_29_161 = _GEN_1111;
  wire          _GEN_1112 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h21;
  wire          compressDataVec_hitReq_30_33;
  assign compressDataVec_hitReq_30_33 = _GEN_1112;
  wire          compressDataVec_hitReq_30_161;
  assign compressDataVec_hitReq_30_161 = _GEN_1112;
  wire          _GEN_1113 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h21;
  wire          compressDataVec_hitReq_31_33;
  assign compressDataVec_hitReq_31_33 = _GEN_1113;
  wire          compressDataVec_hitReq_31_161;
  assign compressDataVec_hitReq_31_161 = _GEN_1113;
  wire          compressDataVec_hitReq_32_33 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h21;
  wire          compressDataVec_hitReq_33_33 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h21;
  wire          compressDataVec_hitReq_34_33 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h21;
  wire          compressDataVec_hitReq_35_33 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h21;
  wire          compressDataVec_hitReq_36_33 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h21;
  wire          compressDataVec_hitReq_37_33 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h21;
  wire          compressDataVec_hitReq_38_33 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h21;
  wire          compressDataVec_hitReq_39_33 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h21;
  wire          compressDataVec_hitReq_40_33 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h21;
  wire          compressDataVec_hitReq_41_33 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h21;
  wire          compressDataVec_hitReq_42_33 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h21;
  wire          compressDataVec_hitReq_43_33 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h21;
  wire          compressDataVec_hitReq_44_33 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h21;
  wire          compressDataVec_hitReq_45_33 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h21;
  wire          compressDataVec_hitReq_46_33 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h21;
  wire          compressDataVec_hitReq_47_33 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h21;
  wire          compressDataVec_hitReq_48_33 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h21;
  wire          compressDataVec_hitReq_49_33 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h21;
  wire          compressDataVec_hitReq_50_33 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h21;
  wire          compressDataVec_hitReq_51_33 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h21;
  wire          compressDataVec_hitReq_52_33 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h21;
  wire          compressDataVec_hitReq_53_33 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h21;
  wire          compressDataVec_hitReq_54_33 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h21;
  wire          compressDataVec_hitReq_55_33 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h21;
  wire          compressDataVec_hitReq_56_33 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h21;
  wire          compressDataVec_hitReq_57_33 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h21;
  wire          compressDataVec_hitReq_58_33 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h21;
  wire          compressDataVec_hitReq_59_33 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h21;
  wire          compressDataVec_hitReq_60_33 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h21;
  wire          compressDataVec_hitReq_61_33 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h21;
  wire          compressDataVec_hitReq_62_33 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h21;
  wire          compressDataVec_hitReq_63_33 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h21;
  wire [7:0]    compressDataVec_selectReqData_33 =
    (compressDataVec_hitReq_0_33 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_33 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_33 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_33 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_33 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_33 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_33 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_33 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_33 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_33 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_33 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_33 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_33 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_33 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_33 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_33 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_33 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_33 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_33 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_33 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_33 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_33 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_33 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_33 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_33 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_33 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_33 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_33 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_33 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_33 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_33 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_33 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_33 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_33 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_33 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_33 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_33 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_33 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_33 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_33 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_33 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_33 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_33 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_33 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_33 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_33 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_33 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_33 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_33 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_33 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_33 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_33 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_33 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_33 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_33 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_33 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_33 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_33 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_33 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_33 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_33 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_33 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_33 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_33 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_33 = tailCount > 6'h21;
  wire          _GEN_1114 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h22;
  wire          compressDataVec_hitReq_0_34;
  assign compressDataVec_hitReq_0_34 = _GEN_1114;
  wire          compressDataVec_hitReq_0_162;
  assign compressDataVec_hitReq_0_162 = _GEN_1114;
  wire          _GEN_1115 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h22;
  wire          compressDataVec_hitReq_1_34;
  assign compressDataVec_hitReq_1_34 = _GEN_1115;
  wire          compressDataVec_hitReq_1_162;
  assign compressDataVec_hitReq_1_162 = _GEN_1115;
  wire          _GEN_1116 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h22;
  wire          compressDataVec_hitReq_2_34;
  assign compressDataVec_hitReq_2_34 = _GEN_1116;
  wire          compressDataVec_hitReq_2_162;
  assign compressDataVec_hitReq_2_162 = _GEN_1116;
  wire          _GEN_1117 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h22;
  wire          compressDataVec_hitReq_3_34;
  assign compressDataVec_hitReq_3_34 = _GEN_1117;
  wire          compressDataVec_hitReq_3_162;
  assign compressDataVec_hitReq_3_162 = _GEN_1117;
  wire          _GEN_1118 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h22;
  wire          compressDataVec_hitReq_4_34;
  assign compressDataVec_hitReq_4_34 = _GEN_1118;
  wire          compressDataVec_hitReq_4_162;
  assign compressDataVec_hitReq_4_162 = _GEN_1118;
  wire          _GEN_1119 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h22;
  wire          compressDataVec_hitReq_5_34;
  assign compressDataVec_hitReq_5_34 = _GEN_1119;
  wire          compressDataVec_hitReq_5_162;
  assign compressDataVec_hitReq_5_162 = _GEN_1119;
  wire          _GEN_1120 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h22;
  wire          compressDataVec_hitReq_6_34;
  assign compressDataVec_hitReq_6_34 = _GEN_1120;
  wire          compressDataVec_hitReq_6_162;
  assign compressDataVec_hitReq_6_162 = _GEN_1120;
  wire          _GEN_1121 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h22;
  wire          compressDataVec_hitReq_7_34;
  assign compressDataVec_hitReq_7_34 = _GEN_1121;
  wire          compressDataVec_hitReq_7_162;
  assign compressDataVec_hitReq_7_162 = _GEN_1121;
  wire          _GEN_1122 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h22;
  wire          compressDataVec_hitReq_8_34;
  assign compressDataVec_hitReq_8_34 = _GEN_1122;
  wire          compressDataVec_hitReq_8_162;
  assign compressDataVec_hitReq_8_162 = _GEN_1122;
  wire          _GEN_1123 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h22;
  wire          compressDataVec_hitReq_9_34;
  assign compressDataVec_hitReq_9_34 = _GEN_1123;
  wire          compressDataVec_hitReq_9_162;
  assign compressDataVec_hitReq_9_162 = _GEN_1123;
  wire          _GEN_1124 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h22;
  wire          compressDataVec_hitReq_10_34;
  assign compressDataVec_hitReq_10_34 = _GEN_1124;
  wire          compressDataVec_hitReq_10_162;
  assign compressDataVec_hitReq_10_162 = _GEN_1124;
  wire          _GEN_1125 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h22;
  wire          compressDataVec_hitReq_11_34;
  assign compressDataVec_hitReq_11_34 = _GEN_1125;
  wire          compressDataVec_hitReq_11_162;
  assign compressDataVec_hitReq_11_162 = _GEN_1125;
  wire          _GEN_1126 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h22;
  wire          compressDataVec_hitReq_12_34;
  assign compressDataVec_hitReq_12_34 = _GEN_1126;
  wire          compressDataVec_hitReq_12_162;
  assign compressDataVec_hitReq_12_162 = _GEN_1126;
  wire          _GEN_1127 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h22;
  wire          compressDataVec_hitReq_13_34;
  assign compressDataVec_hitReq_13_34 = _GEN_1127;
  wire          compressDataVec_hitReq_13_162;
  assign compressDataVec_hitReq_13_162 = _GEN_1127;
  wire          _GEN_1128 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h22;
  wire          compressDataVec_hitReq_14_34;
  assign compressDataVec_hitReq_14_34 = _GEN_1128;
  wire          compressDataVec_hitReq_14_162;
  assign compressDataVec_hitReq_14_162 = _GEN_1128;
  wire          _GEN_1129 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h22;
  wire          compressDataVec_hitReq_15_34;
  assign compressDataVec_hitReq_15_34 = _GEN_1129;
  wire          compressDataVec_hitReq_15_162;
  assign compressDataVec_hitReq_15_162 = _GEN_1129;
  wire          _GEN_1130 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h22;
  wire          compressDataVec_hitReq_16_34;
  assign compressDataVec_hitReq_16_34 = _GEN_1130;
  wire          compressDataVec_hitReq_16_162;
  assign compressDataVec_hitReq_16_162 = _GEN_1130;
  wire          _GEN_1131 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h22;
  wire          compressDataVec_hitReq_17_34;
  assign compressDataVec_hitReq_17_34 = _GEN_1131;
  wire          compressDataVec_hitReq_17_162;
  assign compressDataVec_hitReq_17_162 = _GEN_1131;
  wire          _GEN_1132 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h22;
  wire          compressDataVec_hitReq_18_34;
  assign compressDataVec_hitReq_18_34 = _GEN_1132;
  wire          compressDataVec_hitReq_18_162;
  assign compressDataVec_hitReq_18_162 = _GEN_1132;
  wire          _GEN_1133 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h22;
  wire          compressDataVec_hitReq_19_34;
  assign compressDataVec_hitReq_19_34 = _GEN_1133;
  wire          compressDataVec_hitReq_19_162;
  assign compressDataVec_hitReq_19_162 = _GEN_1133;
  wire          _GEN_1134 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h22;
  wire          compressDataVec_hitReq_20_34;
  assign compressDataVec_hitReq_20_34 = _GEN_1134;
  wire          compressDataVec_hitReq_20_162;
  assign compressDataVec_hitReq_20_162 = _GEN_1134;
  wire          _GEN_1135 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h22;
  wire          compressDataVec_hitReq_21_34;
  assign compressDataVec_hitReq_21_34 = _GEN_1135;
  wire          compressDataVec_hitReq_21_162;
  assign compressDataVec_hitReq_21_162 = _GEN_1135;
  wire          _GEN_1136 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h22;
  wire          compressDataVec_hitReq_22_34;
  assign compressDataVec_hitReq_22_34 = _GEN_1136;
  wire          compressDataVec_hitReq_22_162;
  assign compressDataVec_hitReq_22_162 = _GEN_1136;
  wire          _GEN_1137 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h22;
  wire          compressDataVec_hitReq_23_34;
  assign compressDataVec_hitReq_23_34 = _GEN_1137;
  wire          compressDataVec_hitReq_23_162;
  assign compressDataVec_hitReq_23_162 = _GEN_1137;
  wire          _GEN_1138 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h22;
  wire          compressDataVec_hitReq_24_34;
  assign compressDataVec_hitReq_24_34 = _GEN_1138;
  wire          compressDataVec_hitReq_24_162;
  assign compressDataVec_hitReq_24_162 = _GEN_1138;
  wire          _GEN_1139 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h22;
  wire          compressDataVec_hitReq_25_34;
  assign compressDataVec_hitReq_25_34 = _GEN_1139;
  wire          compressDataVec_hitReq_25_162;
  assign compressDataVec_hitReq_25_162 = _GEN_1139;
  wire          _GEN_1140 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h22;
  wire          compressDataVec_hitReq_26_34;
  assign compressDataVec_hitReq_26_34 = _GEN_1140;
  wire          compressDataVec_hitReq_26_162;
  assign compressDataVec_hitReq_26_162 = _GEN_1140;
  wire          _GEN_1141 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h22;
  wire          compressDataVec_hitReq_27_34;
  assign compressDataVec_hitReq_27_34 = _GEN_1141;
  wire          compressDataVec_hitReq_27_162;
  assign compressDataVec_hitReq_27_162 = _GEN_1141;
  wire          _GEN_1142 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h22;
  wire          compressDataVec_hitReq_28_34;
  assign compressDataVec_hitReq_28_34 = _GEN_1142;
  wire          compressDataVec_hitReq_28_162;
  assign compressDataVec_hitReq_28_162 = _GEN_1142;
  wire          _GEN_1143 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h22;
  wire          compressDataVec_hitReq_29_34;
  assign compressDataVec_hitReq_29_34 = _GEN_1143;
  wire          compressDataVec_hitReq_29_162;
  assign compressDataVec_hitReq_29_162 = _GEN_1143;
  wire          _GEN_1144 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h22;
  wire          compressDataVec_hitReq_30_34;
  assign compressDataVec_hitReq_30_34 = _GEN_1144;
  wire          compressDataVec_hitReq_30_162;
  assign compressDataVec_hitReq_30_162 = _GEN_1144;
  wire          _GEN_1145 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h22;
  wire          compressDataVec_hitReq_31_34;
  assign compressDataVec_hitReq_31_34 = _GEN_1145;
  wire          compressDataVec_hitReq_31_162;
  assign compressDataVec_hitReq_31_162 = _GEN_1145;
  wire          compressDataVec_hitReq_32_34 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h22;
  wire          compressDataVec_hitReq_33_34 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h22;
  wire          compressDataVec_hitReq_34_34 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h22;
  wire          compressDataVec_hitReq_35_34 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h22;
  wire          compressDataVec_hitReq_36_34 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h22;
  wire          compressDataVec_hitReq_37_34 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h22;
  wire          compressDataVec_hitReq_38_34 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h22;
  wire          compressDataVec_hitReq_39_34 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h22;
  wire          compressDataVec_hitReq_40_34 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h22;
  wire          compressDataVec_hitReq_41_34 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h22;
  wire          compressDataVec_hitReq_42_34 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h22;
  wire          compressDataVec_hitReq_43_34 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h22;
  wire          compressDataVec_hitReq_44_34 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h22;
  wire          compressDataVec_hitReq_45_34 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h22;
  wire          compressDataVec_hitReq_46_34 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h22;
  wire          compressDataVec_hitReq_47_34 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h22;
  wire          compressDataVec_hitReq_48_34 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h22;
  wire          compressDataVec_hitReq_49_34 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h22;
  wire          compressDataVec_hitReq_50_34 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h22;
  wire          compressDataVec_hitReq_51_34 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h22;
  wire          compressDataVec_hitReq_52_34 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h22;
  wire          compressDataVec_hitReq_53_34 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h22;
  wire          compressDataVec_hitReq_54_34 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h22;
  wire          compressDataVec_hitReq_55_34 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h22;
  wire          compressDataVec_hitReq_56_34 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h22;
  wire          compressDataVec_hitReq_57_34 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h22;
  wire          compressDataVec_hitReq_58_34 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h22;
  wire          compressDataVec_hitReq_59_34 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h22;
  wire          compressDataVec_hitReq_60_34 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h22;
  wire          compressDataVec_hitReq_61_34 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h22;
  wire          compressDataVec_hitReq_62_34 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h22;
  wire          compressDataVec_hitReq_63_34 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h22;
  wire [7:0]    compressDataVec_selectReqData_34 =
    (compressDataVec_hitReq_0_34 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_34 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_34 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_34 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_34 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_34 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_34 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_34 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_34 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_34 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_34 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_34 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_34 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_34 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_34 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_34 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_34 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_34 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_34 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_34 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_34 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_34 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_34 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_34 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_34 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_34 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_34 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_34 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_34 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_34 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_34 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_34 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_34 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_34 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_34 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_34 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_34 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_34 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_34 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_34 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_34 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_34 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_34 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_34 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_34 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_34 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_34 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_34 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_34 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_34 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_34 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_34 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_34 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_34 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_34 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_34 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_34 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_34 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_34 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_34 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_34 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_34 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_34 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_34 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_34 = tailCount > 6'h22;
  wire          _GEN_1146 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h23;
  wire          compressDataVec_hitReq_0_35;
  assign compressDataVec_hitReq_0_35 = _GEN_1146;
  wire          compressDataVec_hitReq_0_163;
  assign compressDataVec_hitReq_0_163 = _GEN_1146;
  wire          _GEN_1147 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h23;
  wire          compressDataVec_hitReq_1_35;
  assign compressDataVec_hitReq_1_35 = _GEN_1147;
  wire          compressDataVec_hitReq_1_163;
  assign compressDataVec_hitReq_1_163 = _GEN_1147;
  wire          _GEN_1148 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h23;
  wire          compressDataVec_hitReq_2_35;
  assign compressDataVec_hitReq_2_35 = _GEN_1148;
  wire          compressDataVec_hitReq_2_163;
  assign compressDataVec_hitReq_2_163 = _GEN_1148;
  wire          _GEN_1149 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h23;
  wire          compressDataVec_hitReq_3_35;
  assign compressDataVec_hitReq_3_35 = _GEN_1149;
  wire          compressDataVec_hitReq_3_163;
  assign compressDataVec_hitReq_3_163 = _GEN_1149;
  wire          _GEN_1150 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h23;
  wire          compressDataVec_hitReq_4_35;
  assign compressDataVec_hitReq_4_35 = _GEN_1150;
  wire          compressDataVec_hitReq_4_163;
  assign compressDataVec_hitReq_4_163 = _GEN_1150;
  wire          _GEN_1151 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h23;
  wire          compressDataVec_hitReq_5_35;
  assign compressDataVec_hitReq_5_35 = _GEN_1151;
  wire          compressDataVec_hitReq_5_163;
  assign compressDataVec_hitReq_5_163 = _GEN_1151;
  wire          _GEN_1152 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h23;
  wire          compressDataVec_hitReq_6_35;
  assign compressDataVec_hitReq_6_35 = _GEN_1152;
  wire          compressDataVec_hitReq_6_163;
  assign compressDataVec_hitReq_6_163 = _GEN_1152;
  wire          _GEN_1153 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h23;
  wire          compressDataVec_hitReq_7_35;
  assign compressDataVec_hitReq_7_35 = _GEN_1153;
  wire          compressDataVec_hitReq_7_163;
  assign compressDataVec_hitReq_7_163 = _GEN_1153;
  wire          _GEN_1154 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h23;
  wire          compressDataVec_hitReq_8_35;
  assign compressDataVec_hitReq_8_35 = _GEN_1154;
  wire          compressDataVec_hitReq_8_163;
  assign compressDataVec_hitReq_8_163 = _GEN_1154;
  wire          _GEN_1155 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h23;
  wire          compressDataVec_hitReq_9_35;
  assign compressDataVec_hitReq_9_35 = _GEN_1155;
  wire          compressDataVec_hitReq_9_163;
  assign compressDataVec_hitReq_9_163 = _GEN_1155;
  wire          _GEN_1156 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h23;
  wire          compressDataVec_hitReq_10_35;
  assign compressDataVec_hitReq_10_35 = _GEN_1156;
  wire          compressDataVec_hitReq_10_163;
  assign compressDataVec_hitReq_10_163 = _GEN_1156;
  wire          _GEN_1157 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h23;
  wire          compressDataVec_hitReq_11_35;
  assign compressDataVec_hitReq_11_35 = _GEN_1157;
  wire          compressDataVec_hitReq_11_163;
  assign compressDataVec_hitReq_11_163 = _GEN_1157;
  wire          _GEN_1158 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h23;
  wire          compressDataVec_hitReq_12_35;
  assign compressDataVec_hitReq_12_35 = _GEN_1158;
  wire          compressDataVec_hitReq_12_163;
  assign compressDataVec_hitReq_12_163 = _GEN_1158;
  wire          _GEN_1159 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h23;
  wire          compressDataVec_hitReq_13_35;
  assign compressDataVec_hitReq_13_35 = _GEN_1159;
  wire          compressDataVec_hitReq_13_163;
  assign compressDataVec_hitReq_13_163 = _GEN_1159;
  wire          _GEN_1160 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h23;
  wire          compressDataVec_hitReq_14_35;
  assign compressDataVec_hitReq_14_35 = _GEN_1160;
  wire          compressDataVec_hitReq_14_163;
  assign compressDataVec_hitReq_14_163 = _GEN_1160;
  wire          _GEN_1161 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h23;
  wire          compressDataVec_hitReq_15_35;
  assign compressDataVec_hitReq_15_35 = _GEN_1161;
  wire          compressDataVec_hitReq_15_163;
  assign compressDataVec_hitReq_15_163 = _GEN_1161;
  wire          _GEN_1162 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h23;
  wire          compressDataVec_hitReq_16_35;
  assign compressDataVec_hitReq_16_35 = _GEN_1162;
  wire          compressDataVec_hitReq_16_163;
  assign compressDataVec_hitReq_16_163 = _GEN_1162;
  wire          _GEN_1163 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h23;
  wire          compressDataVec_hitReq_17_35;
  assign compressDataVec_hitReq_17_35 = _GEN_1163;
  wire          compressDataVec_hitReq_17_163;
  assign compressDataVec_hitReq_17_163 = _GEN_1163;
  wire          _GEN_1164 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h23;
  wire          compressDataVec_hitReq_18_35;
  assign compressDataVec_hitReq_18_35 = _GEN_1164;
  wire          compressDataVec_hitReq_18_163;
  assign compressDataVec_hitReq_18_163 = _GEN_1164;
  wire          _GEN_1165 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h23;
  wire          compressDataVec_hitReq_19_35;
  assign compressDataVec_hitReq_19_35 = _GEN_1165;
  wire          compressDataVec_hitReq_19_163;
  assign compressDataVec_hitReq_19_163 = _GEN_1165;
  wire          _GEN_1166 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h23;
  wire          compressDataVec_hitReq_20_35;
  assign compressDataVec_hitReq_20_35 = _GEN_1166;
  wire          compressDataVec_hitReq_20_163;
  assign compressDataVec_hitReq_20_163 = _GEN_1166;
  wire          _GEN_1167 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h23;
  wire          compressDataVec_hitReq_21_35;
  assign compressDataVec_hitReq_21_35 = _GEN_1167;
  wire          compressDataVec_hitReq_21_163;
  assign compressDataVec_hitReq_21_163 = _GEN_1167;
  wire          _GEN_1168 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h23;
  wire          compressDataVec_hitReq_22_35;
  assign compressDataVec_hitReq_22_35 = _GEN_1168;
  wire          compressDataVec_hitReq_22_163;
  assign compressDataVec_hitReq_22_163 = _GEN_1168;
  wire          _GEN_1169 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h23;
  wire          compressDataVec_hitReq_23_35;
  assign compressDataVec_hitReq_23_35 = _GEN_1169;
  wire          compressDataVec_hitReq_23_163;
  assign compressDataVec_hitReq_23_163 = _GEN_1169;
  wire          _GEN_1170 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h23;
  wire          compressDataVec_hitReq_24_35;
  assign compressDataVec_hitReq_24_35 = _GEN_1170;
  wire          compressDataVec_hitReq_24_163;
  assign compressDataVec_hitReq_24_163 = _GEN_1170;
  wire          _GEN_1171 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h23;
  wire          compressDataVec_hitReq_25_35;
  assign compressDataVec_hitReq_25_35 = _GEN_1171;
  wire          compressDataVec_hitReq_25_163;
  assign compressDataVec_hitReq_25_163 = _GEN_1171;
  wire          _GEN_1172 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h23;
  wire          compressDataVec_hitReq_26_35;
  assign compressDataVec_hitReq_26_35 = _GEN_1172;
  wire          compressDataVec_hitReq_26_163;
  assign compressDataVec_hitReq_26_163 = _GEN_1172;
  wire          _GEN_1173 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h23;
  wire          compressDataVec_hitReq_27_35;
  assign compressDataVec_hitReq_27_35 = _GEN_1173;
  wire          compressDataVec_hitReq_27_163;
  assign compressDataVec_hitReq_27_163 = _GEN_1173;
  wire          _GEN_1174 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h23;
  wire          compressDataVec_hitReq_28_35;
  assign compressDataVec_hitReq_28_35 = _GEN_1174;
  wire          compressDataVec_hitReq_28_163;
  assign compressDataVec_hitReq_28_163 = _GEN_1174;
  wire          _GEN_1175 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h23;
  wire          compressDataVec_hitReq_29_35;
  assign compressDataVec_hitReq_29_35 = _GEN_1175;
  wire          compressDataVec_hitReq_29_163;
  assign compressDataVec_hitReq_29_163 = _GEN_1175;
  wire          _GEN_1176 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h23;
  wire          compressDataVec_hitReq_30_35;
  assign compressDataVec_hitReq_30_35 = _GEN_1176;
  wire          compressDataVec_hitReq_30_163;
  assign compressDataVec_hitReq_30_163 = _GEN_1176;
  wire          _GEN_1177 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h23;
  wire          compressDataVec_hitReq_31_35;
  assign compressDataVec_hitReq_31_35 = _GEN_1177;
  wire          compressDataVec_hitReq_31_163;
  assign compressDataVec_hitReq_31_163 = _GEN_1177;
  wire          compressDataVec_hitReq_32_35 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h23;
  wire          compressDataVec_hitReq_33_35 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h23;
  wire          compressDataVec_hitReq_34_35 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h23;
  wire          compressDataVec_hitReq_35_35 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h23;
  wire          compressDataVec_hitReq_36_35 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h23;
  wire          compressDataVec_hitReq_37_35 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h23;
  wire          compressDataVec_hitReq_38_35 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h23;
  wire          compressDataVec_hitReq_39_35 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h23;
  wire          compressDataVec_hitReq_40_35 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h23;
  wire          compressDataVec_hitReq_41_35 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h23;
  wire          compressDataVec_hitReq_42_35 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h23;
  wire          compressDataVec_hitReq_43_35 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h23;
  wire          compressDataVec_hitReq_44_35 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h23;
  wire          compressDataVec_hitReq_45_35 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h23;
  wire          compressDataVec_hitReq_46_35 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h23;
  wire          compressDataVec_hitReq_47_35 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h23;
  wire          compressDataVec_hitReq_48_35 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h23;
  wire          compressDataVec_hitReq_49_35 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h23;
  wire          compressDataVec_hitReq_50_35 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h23;
  wire          compressDataVec_hitReq_51_35 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h23;
  wire          compressDataVec_hitReq_52_35 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h23;
  wire          compressDataVec_hitReq_53_35 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h23;
  wire          compressDataVec_hitReq_54_35 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h23;
  wire          compressDataVec_hitReq_55_35 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h23;
  wire          compressDataVec_hitReq_56_35 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h23;
  wire          compressDataVec_hitReq_57_35 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h23;
  wire          compressDataVec_hitReq_58_35 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h23;
  wire          compressDataVec_hitReq_59_35 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h23;
  wire          compressDataVec_hitReq_60_35 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h23;
  wire          compressDataVec_hitReq_61_35 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h23;
  wire          compressDataVec_hitReq_62_35 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h23;
  wire          compressDataVec_hitReq_63_35 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h23;
  wire [7:0]    compressDataVec_selectReqData_35 =
    (compressDataVec_hitReq_0_35 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_35 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_35 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_35 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_35 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_35 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_35 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_35 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_35 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_35 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_35 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_35 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_35 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_35 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_35 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_35 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_35 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_35 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_35 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_35 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_35 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_35 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_35 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_35 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_35 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_35 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_35 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_35 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_35 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_35 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_35 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_35 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_35 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_35 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_35 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_35 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_35 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_35 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_35 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_35 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_35 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_35 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_35 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_35 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_35 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_35 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_35 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_35 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_35 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_35 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_35 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_35 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_35 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_35 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_35 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_35 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_35 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_35 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_35 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_35 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_35 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_35 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_35 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_35 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_35 = tailCount > 6'h23;
  wire          _GEN_1178 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h24;
  wire          compressDataVec_hitReq_0_36;
  assign compressDataVec_hitReq_0_36 = _GEN_1178;
  wire          compressDataVec_hitReq_0_164;
  assign compressDataVec_hitReq_0_164 = _GEN_1178;
  wire          _GEN_1179 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h24;
  wire          compressDataVec_hitReq_1_36;
  assign compressDataVec_hitReq_1_36 = _GEN_1179;
  wire          compressDataVec_hitReq_1_164;
  assign compressDataVec_hitReq_1_164 = _GEN_1179;
  wire          _GEN_1180 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h24;
  wire          compressDataVec_hitReq_2_36;
  assign compressDataVec_hitReq_2_36 = _GEN_1180;
  wire          compressDataVec_hitReq_2_164;
  assign compressDataVec_hitReq_2_164 = _GEN_1180;
  wire          _GEN_1181 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h24;
  wire          compressDataVec_hitReq_3_36;
  assign compressDataVec_hitReq_3_36 = _GEN_1181;
  wire          compressDataVec_hitReq_3_164;
  assign compressDataVec_hitReq_3_164 = _GEN_1181;
  wire          _GEN_1182 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h24;
  wire          compressDataVec_hitReq_4_36;
  assign compressDataVec_hitReq_4_36 = _GEN_1182;
  wire          compressDataVec_hitReq_4_164;
  assign compressDataVec_hitReq_4_164 = _GEN_1182;
  wire          _GEN_1183 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h24;
  wire          compressDataVec_hitReq_5_36;
  assign compressDataVec_hitReq_5_36 = _GEN_1183;
  wire          compressDataVec_hitReq_5_164;
  assign compressDataVec_hitReq_5_164 = _GEN_1183;
  wire          _GEN_1184 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h24;
  wire          compressDataVec_hitReq_6_36;
  assign compressDataVec_hitReq_6_36 = _GEN_1184;
  wire          compressDataVec_hitReq_6_164;
  assign compressDataVec_hitReq_6_164 = _GEN_1184;
  wire          _GEN_1185 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h24;
  wire          compressDataVec_hitReq_7_36;
  assign compressDataVec_hitReq_7_36 = _GEN_1185;
  wire          compressDataVec_hitReq_7_164;
  assign compressDataVec_hitReq_7_164 = _GEN_1185;
  wire          _GEN_1186 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h24;
  wire          compressDataVec_hitReq_8_36;
  assign compressDataVec_hitReq_8_36 = _GEN_1186;
  wire          compressDataVec_hitReq_8_164;
  assign compressDataVec_hitReq_8_164 = _GEN_1186;
  wire          _GEN_1187 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h24;
  wire          compressDataVec_hitReq_9_36;
  assign compressDataVec_hitReq_9_36 = _GEN_1187;
  wire          compressDataVec_hitReq_9_164;
  assign compressDataVec_hitReq_9_164 = _GEN_1187;
  wire          _GEN_1188 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h24;
  wire          compressDataVec_hitReq_10_36;
  assign compressDataVec_hitReq_10_36 = _GEN_1188;
  wire          compressDataVec_hitReq_10_164;
  assign compressDataVec_hitReq_10_164 = _GEN_1188;
  wire          _GEN_1189 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h24;
  wire          compressDataVec_hitReq_11_36;
  assign compressDataVec_hitReq_11_36 = _GEN_1189;
  wire          compressDataVec_hitReq_11_164;
  assign compressDataVec_hitReq_11_164 = _GEN_1189;
  wire          _GEN_1190 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h24;
  wire          compressDataVec_hitReq_12_36;
  assign compressDataVec_hitReq_12_36 = _GEN_1190;
  wire          compressDataVec_hitReq_12_164;
  assign compressDataVec_hitReq_12_164 = _GEN_1190;
  wire          _GEN_1191 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h24;
  wire          compressDataVec_hitReq_13_36;
  assign compressDataVec_hitReq_13_36 = _GEN_1191;
  wire          compressDataVec_hitReq_13_164;
  assign compressDataVec_hitReq_13_164 = _GEN_1191;
  wire          _GEN_1192 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h24;
  wire          compressDataVec_hitReq_14_36;
  assign compressDataVec_hitReq_14_36 = _GEN_1192;
  wire          compressDataVec_hitReq_14_164;
  assign compressDataVec_hitReq_14_164 = _GEN_1192;
  wire          _GEN_1193 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h24;
  wire          compressDataVec_hitReq_15_36;
  assign compressDataVec_hitReq_15_36 = _GEN_1193;
  wire          compressDataVec_hitReq_15_164;
  assign compressDataVec_hitReq_15_164 = _GEN_1193;
  wire          _GEN_1194 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h24;
  wire          compressDataVec_hitReq_16_36;
  assign compressDataVec_hitReq_16_36 = _GEN_1194;
  wire          compressDataVec_hitReq_16_164;
  assign compressDataVec_hitReq_16_164 = _GEN_1194;
  wire          _GEN_1195 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h24;
  wire          compressDataVec_hitReq_17_36;
  assign compressDataVec_hitReq_17_36 = _GEN_1195;
  wire          compressDataVec_hitReq_17_164;
  assign compressDataVec_hitReq_17_164 = _GEN_1195;
  wire          _GEN_1196 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h24;
  wire          compressDataVec_hitReq_18_36;
  assign compressDataVec_hitReq_18_36 = _GEN_1196;
  wire          compressDataVec_hitReq_18_164;
  assign compressDataVec_hitReq_18_164 = _GEN_1196;
  wire          _GEN_1197 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h24;
  wire          compressDataVec_hitReq_19_36;
  assign compressDataVec_hitReq_19_36 = _GEN_1197;
  wire          compressDataVec_hitReq_19_164;
  assign compressDataVec_hitReq_19_164 = _GEN_1197;
  wire          _GEN_1198 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h24;
  wire          compressDataVec_hitReq_20_36;
  assign compressDataVec_hitReq_20_36 = _GEN_1198;
  wire          compressDataVec_hitReq_20_164;
  assign compressDataVec_hitReq_20_164 = _GEN_1198;
  wire          _GEN_1199 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h24;
  wire          compressDataVec_hitReq_21_36;
  assign compressDataVec_hitReq_21_36 = _GEN_1199;
  wire          compressDataVec_hitReq_21_164;
  assign compressDataVec_hitReq_21_164 = _GEN_1199;
  wire          _GEN_1200 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h24;
  wire          compressDataVec_hitReq_22_36;
  assign compressDataVec_hitReq_22_36 = _GEN_1200;
  wire          compressDataVec_hitReq_22_164;
  assign compressDataVec_hitReq_22_164 = _GEN_1200;
  wire          _GEN_1201 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h24;
  wire          compressDataVec_hitReq_23_36;
  assign compressDataVec_hitReq_23_36 = _GEN_1201;
  wire          compressDataVec_hitReq_23_164;
  assign compressDataVec_hitReq_23_164 = _GEN_1201;
  wire          _GEN_1202 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h24;
  wire          compressDataVec_hitReq_24_36;
  assign compressDataVec_hitReq_24_36 = _GEN_1202;
  wire          compressDataVec_hitReq_24_164;
  assign compressDataVec_hitReq_24_164 = _GEN_1202;
  wire          _GEN_1203 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h24;
  wire          compressDataVec_hitReq_25_36;
  assign compressDataVec_hitReq_25_36 = _GEN_1203;
  wire          compressDataVec_hitReq_25_164;
  assign compressDataVec_hitReq_25_164 = _GEN_1203;
  wire          _GEN_1204 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h24;
  wire          compressDataVec_hitReq_26_36;
  assign compressDataVec_hitReq_26_36 = _GEN_1204;
  wire          compressDataVec_hitReq_26_164;
  assign compressDataVec_hitReq_26_164 = _GEN_1204;
  wire          _GEN_1205 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h24;
  wire          compressDataVec_hitReq_27_36;
  assign compressDataVec_hitReq_27_36 = _GEN_1205;
  wire          compressDataVec_hitReq_27_164;
  assign compressDataVec_hitReq_27_164 = _GEN_1205;
  wire          _GEN_1206 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h24;
  wire          compressDataVec_hitReq_28_36;
  assign compressDataVec_hitReq_28_36 = _GEN_1206;
  wire          compressDataVec_hitReq_28_164;
  assign compressDataVec_hitReq_28_164 = _GEN_1206;
  wire          _GEN_1207 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h24;
  wire          compressDataVec_hitReq_29_36;
  assign compressDataVec_hitReq_29_36 = _GEN_1207;
  wire          compressDataVec_hitReq_29_164;
  assign compressDataVec_hitReq_29_164 = _GEN_1207;
  wire          _GEN_1208 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h24;
  wire          compressDataVec_hitReq_30_36;
  assign compressDataVec_hitReq_30_36 = _GEN_1208;
  wire          compressDataVec_hitReq_30_164;
  assign compressDataVec_hitReq_30_164 = _GEN_1208;
  wire          _GEN_1209 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h24;
  wire          compressDataVec_hitReq_31_36;
  assign compressDataVec_hitReq_31_36 = _GEN_1209;
  wire          compressDataVec_hitReq_31_164;
  assign compressDataVec_hitReq_31_164 = _GEN_1209;
  wire          compressDataVec_hitReq_32_36 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h24;
  wire          compressDataVec_hitReq_33_36 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h24;
  wire          compressDataVec_hitReq_34_36 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h24;
  wire          compressDataVec_hitReq_35_36 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h24;
  wire          compressDataVec_hitReq_36_36 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h24;
  wire          compressDataVec_hitReq_37_36 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h24;
  wire          compressDataVec_hitReq_38_36 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h24;
  wire          compressDataVec_hitReq_39_36 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h24;
  wire          compressDataVec_hitReq_40_36 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h24;
  wire          compressDataVec_hitReq_41_36 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h24;
  wire          compressDataVec_hitReq_42_36 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h24;
  wire          compressDataVec_hitReq_43_36 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h24;
  wire          compressDataVec_hitReq_44_36 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h24;
  wire          compressDataVec_hitReq_45_36 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h24;
  wire          compressDataVec_hitReq_46_36 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h24;
  wire          compressDataVec_hitReq_47_36 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h24;
  wire          compressDataVec_hitReq_48_36 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h24;
  wire          compressDataVec_hitReq_49_36 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h24;
  wire          compressDataVec_hitReq_50_36 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h24;
  wire          compressDataVec_hitReq_51_36 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h24;
  wire          compressDataVec_hitReq_52_36 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h24;
  wire          compressDataVec_hitReq_53_36 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h24;
  wire          compressDataVec_hitReq_54_36 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h24;
  wire          compressDataVec_hitReq_55_36 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h24;
  wire          compressDataVec_hitReq_56_36 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h24;
  wire          compressDataVec_hitReq_57_36 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h24;
  wire          compressDataVec_hitReq_58_36 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h24;
  wire          compressDataVec_hitReq_59_36 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h24;
  wire          compressDataVec_hitReq_60_36 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h24;
  wire          compressDataVec_hitReq_61_36 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h24;
  wire          compressDataVec_hitReq_62_36 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h24;
  wire          compressDataVec_hitReq_63_36 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h24;
  wire [7:0]    compressDataVec_selectReqData_36 =
    (compressDataVec_hitReq_0_36 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_36 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_36 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_36 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_36 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_36 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_36 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_36 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_36 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_36 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_36 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_36 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_36 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_36 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_36 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_36 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_36 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_36 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_36 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_36 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_36 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_36 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_36 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_36 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_36 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_36 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_36 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_36 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_36 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_36 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_36 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_36 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_36 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_36 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_36 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_36 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_36 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_36 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_36 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_36 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_36 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_36 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_36 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_36 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_36 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_36 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_36 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_36 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_36 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_36 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_36 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_36 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_36 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_36 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_36 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_36 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_36 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_36 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_36 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_36 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_36 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_36 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_36 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_36 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_36 = tailCount > 6'h24;
  wire          _GEN_1210 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h25;
  wire          compressDataVec_hitReq_0_37;
  assign compressDataVec_hitReq_0_37 = _GEN_1210;
  wire          compressDataVec_hitReq_0_165;
  assign compressDataVec_hitReq_0_165 = _GEN_1210;
  wire          _GEN_1211 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h25;
  wire          compressDataVec_hitReq_1_37;
  assign compressDataVec_hitReq_1_37 = _GEN_1211;
  wire          compressDataVec_hitReq_1_165;
  assign compressDataVec_hitReq_1_165 = _GEN_1211;
  wire          _GEN_1212 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h25;
  wire          compressDataVec_hitReq_2_37;
  assign compressDataVec_hitReq_2_37 = _GEN_1212;
  wire          compressDataVec_hitReq_2_165;
  assign compressDataVec_hitReq_2_165 = _GEN_1212;
  wire          _GEN_1213 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h25;
  wire          compressDataVec_hitReq_3_37;
  assign compressDataVec_hitReq_3_37 = _GEN_1213;
  wire          compressDataVec_hitReq_3_165;
  assign compressDataVec_hitReq_3_165 = _GEN_1213;
  wire          _GEN_1214 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h25;
  wire          compressDataVec_hitReq_4_37;
  assign compressDataVec_hitReq_4_37 = _GEN_1214;
  wire          compressDataVec_hitReq_4_165;
  assign compressDataVec_hitReq_4_165 = _GEN_1214;
  wire          _GEN_1215 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h25;
  wire          compressDataVec_hitReq_5_37;
  assign compressDataVec_hitReq_5_37 = _GEN_1215;
  wire          compressDataVec_hitReq_5_165;
  assign compressDataVec_hitReq_5_165 = _GEN_1215;
  wire          _GEN_1216 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h25;
  wire          compressDataVec_hitReq_6_37;
  assign compressDataVec_hitReq_6_37 = _GEN_1216;
  wire          compressDataVec_hitReq_6_165;
  assign compressDataVec_hitReq_6_165 = _GEN_1216;
  wire          _GEN_1217 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h25;
  wire          compressDataVec_hitReq_7_37;
  assign compressDataVec_hitReq_7_37 = _GEN_1217;
  wire          compressDataVec_hitReq_7_165;
  assign compressDataVec_hitReq_7_165 = _GEN_1217;
  wire          _GEN_1218 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h25;
  wire          compressDataVec_hitReq_8_37;
  assign compressDataVec_hitReq_8_37 = _GEN_1218;
  wire          compressDataVec_hitReq_8_165;
  assign compressDataVec_hitReq_8_165 = _GEN_1218;
  wire          _GEN_1219 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h25;
  wire          compressDataVec_hitReq_9_37;
  assign compressDataVec_hitReq_9_37 = _GEN_1219;
  wire          compressDataVec_hitReq_9_165;
  assign compressDataVec_hitReq_9_165 = _GEN_1219;
  wire          _GEN_1220 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h25;
  wire          compressDataVec_hitReq_10_37;
  assign compressDataVec_hitReq_10_37 = _GEN_1220;
  wire          compressDataVec_hitReq_10_165;
  assign compressDataVec_hitReq_10_165 = _GEN_1220;
  wire          _GEN_1221 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h25;
  wire          compressDataVec_hitReq_11_37;
  assign compressDataVec_hitReq_11_37 = _GEN_1221;
  wire          compressDataVec_hitReq_11_165;
  assign compressDataVec_hitReq_11_165 = _GEN_1221;
  wire          _GEN_1222 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h25;
  wire          compressDataVec_hitReq_12_37;
  assign compressDataVec_hitReq_12_37 = _GEN_1222;
  wire          compressDataVec_hitReq_12_165;
  assign compressDataVec_hitReq_12_165 = _GEN_1222;
  wire          _GEN_1223 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h25;
  wire          compressDataVec_hitReq_13_37;
  assign compressDataVec_hitReq_13_37 = _GEN_1223;
  wire          compressDataVec_hitReq_13_165;
  assign compressDataVec_hitReq_13_165 = _GEN_1223;
  wire          _GEN_1224 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h25;
  wire          compressDataVec_hitReq_14_37;
  assign compressDataVec_hitReq_14_37 = _GEN_1224;
  wire          compressDataVec_hitReq_14_165;
  assign compressDataVec_hitReq_14_165 = _GEN_1224;
  wire          _GEN_1225 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h25;
  wire          compressDataVec_hitReq_15_37;
  assign compressDataVec_hitReq_15_37 = _GEN_1225;
  wire          compressDataVec_hitReq_15_165;
  assign compressDataVec_hitReq_15_165 = _GEN_1225;
  wire          _GEN_1226 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h25;
  wire          compressDataVec_hitReq_16_37;
  assign compressDataVec_hitReq_16_37 = _GEN_1226;
  wire          compressDataVec_hitReq_16_165;
  assign compressDataVec_hitReq_16_165 = _GEN_1226;
  wire          _GEN_1227 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h25;
  wire          compressDataVec_hitReq_17_37;
  assign compressDataVec_hitReq_17_37 = _GEN_1227;
  wire          compressDataVec_hitReq_17_165;
  assign compressDataVec_hitReq_17_165 = _GEN_1227;
  wire          _GEN_1228 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h25;
  wire          compressDataVec_hitReq_18_37;
  assign compressDataVec_hitReq_18_37 = _GEN_1228;
  wire          compressDataVec_hitReq_18_165;
  assign compressDataVec_hitReq_18_165 = _GEN_1228;
  wire          _GEN_1229 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h25;
  wire          compressDataVec_hitReq_19_37;
  assign compressDataVec_hitReq_19_37 = _GEN_1229;
  wire          compressDataVec_hitReq_19_165;
  assign compressDataVec_hitReq_19_165 = _GEN_1229;
  wire          _GEN_1230 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h25;
  wire          compressDataVec_hitReq_20_37;
  assign compressDataVec_hitReq_20_37 = _GEN_1230;
  wire          compressDataVec_hitReq_20_165;
  assign compressDataVec_hitReq_20_165 = _GEN_1230;
  wire          _GEN_1231 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h25;
  wire          compressDataVec_hitReq_21_37;
  assign compressDataVec_hitReq_21_37 = _GEN_1231;
  wire          compressDataVec_hitReq_21_165;
  assign compressDataVec_hitReq_21_165 = _GEN_1231;
  wire          _GEN_1232 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h25;
  wire          compressDataVec_hitReq_22_37;
  assign compressDataVec_hitReq_22_37 = _GEN_1232;
  wire          compressDataVec_hitReq_22_165;
  assign compressDataVec_hitReq_22_165 = _GEN_1232;
  wire          _GEN_1233 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h25;
  wire          compressDataVec_hitReq_23_37;
  assign compressDataVec_hitReq_23_37 = _GEN_1233;
  wire          compressDataVec_hitReq_23_165;
  assign compressDataVec_hitReq_23_165 = _GEN_1233;
  wire          _GEN_1234 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h25;
  wire          compressDataVec_hitReq_24_37;
  assign compressDataVec_hitReq_24_37 = _GEN_1234;
  wire          compressDataVec_hitReq_24_165;
  assign compressDataVec_hitReq_24_165 = _GEN_1234;
  wire          _GEN_1235 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h25;
  wire          compressDataVec_hitReq_25_37;
  assign compressDataVec_hitReq_25_37 = _GEN_1235;
  wire          compressDataVec_hitReq_25_165;
  assign compressDataVec_hitReq_25_165 = _GEN_1235;
  wire          _GEN_1236 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h25;
  wire          compressDataVec_hitReq_26_37;
  assign compressDataVec_hitReq_26_37 = _GEN_1236;
  wire          compressDataVec_hitReq_26_165;
  assign compressDataVec_hitReq_26_165 = _GEN_1236;
  wire          _GEN_1237 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h25;
  wire          compressDataVec_hitReq_27_37;
  assign compressDataVec_hitReq_27_37 = _GEN_1237;
  wire          compressDataVec_hitReq_27_165;
  assign compressDataVec_hitReq_27_165 = _GEN_1237;
  wire          _GEN_1238 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h25;
  wire          compressDataVec_hitReq_28_37;
  assign compressDataVec_hitReq_28_37 = _GEN_1238;
  wire          compressDataVec_hitReq_28_165;
  assign compressDataVec_hitReq_28_165 = _GEN_1238;
  wire          _GEN_1239 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h25;
  wire          compressDataVec_hitReq_29_37;
  assign compressDataVec_hitReq_29_37 = _GEN_1239;
  wire          compressDataVec_hitReq_29_165;
  assign compressDataVec_hitReq_29_165 = _GEN_1239;
  wire          _GEN_1240 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h25;
  wire          compressDataVec_hitReq_30_37;
  assign compressDataVec_hitReq_30_37 = _GEN_1240;
  wire          compressDataVec_hitReq_30_165;
  assign compressDataVec_hitReq_30_165 = _GEN_1240;
  wire          _GEN_1241 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h25;
  wire          compressDataVec_hitReq_31_37;
  assign compressDataVec_hitReq_31_37 = _GEN_1241;
  wire          compressDataVec_hitReq_31_165;
  assign compressDataVec_hitReq_31_165 = _GEN_1241;
  wire          compressDataVec_hitReq_32_37 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h25;
  wire          compressDataVec_hitReq_33_37 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h25;
  wire          compressDataVec_hitReq_34_37 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h25;
  wire          compressDataVec_hitReq_35_37 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h25;
  wire          compressDataVec_hitReq_36_37 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h25;
  wire          compressDataVec_hitReq_37_37 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h25;
  wire          compressDataVec_hitReq_38_37 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h25;
  wire          compressDataVec_hitReq_39_37 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h25;
  wire          compressDataVec_hitReq_40_37 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h25;
  wire          compressDataVec_hitReq_41_37 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h25;
  wire          compressDataVec_hitReq_42_37 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h25;
  wire          compressDataVec_hitReq_43_37 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h25;
  wire          compressDataVec_hitReq_44_37 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h25;
  wire          compressDataVec_hitReq_45_37 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h25;
  wire          compressDataVec_hitReq_46_37 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h25;
  wire          compressDataVec_hitReq_47_37 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h25;
  wire          compressDataVec_hitReq_48_37 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h25;
  wire          compressDataVec_hitReq_49_37 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h25;
  wire          compressDataVec_hitReq_50_37 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h25;
  wire          compressDataVec_hitReq_51_37 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h25;
  wire          compressDataVec_hitReq_52_37 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h25;
  wire          compressDataVec_hitReq_53_37 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h25;
  wire          compressDataVec_hitReq_54_37 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h25;
  wire          compressDataVec_hitReq_55_37 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h25;
  wire          compressDataVec_hitReq_56_37 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h25;
  wire          compressDataVec_hitReq_57_37 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h25;
  wire          compressDataVec_hitReq_58_37 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h25;
  wire          compressDataVec_hitReq_59_37 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h25;
  wire          compressDataVec_hitReq_60_37 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h25;
  wire          compressDataVec_hitReq_61_37 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h25;
  wire          compressDataVec_hitReq_62_37 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h25;
  wire          compressDataVec_hitReq_63_37 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h25;
  wire [7:0]    compressDataVec_selectReqData_37 =
    (compressDataVec_hitReq_0_37 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_37 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_37 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_37 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_37 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_37 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_37 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_37 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_37 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_37 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_37 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_37 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_37 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_37 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_37 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_37 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_37 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_37 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_37 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_37 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_37 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_37 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_37 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_37 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_37 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_37 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_37 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_37 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_37 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_37 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_37 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_37 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_37 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_37 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_37 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_37 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_37 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_37 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_37 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_37 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_37 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_37 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_37 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_37 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_37 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_37 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_37 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_37 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_37 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_37 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_37 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_37 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_37 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_37 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_37 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_37 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_37 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_37 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_37 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_37 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_37 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_37 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_37 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_37 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_37 = tailCount > 6'h25;
  wire          _GEN_1242 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h26;
  wire          compressDataVec_hitReq_0_38;
  assign compressDataVec_hitReq_0_38 = _GEN_1242;
  wire          compressDataVec_hitReq_0_166;
  assign compressDataVec_hitReq_0_166 = _GEN_1242;
  wire          _GEN_1243 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h26;
  wire          compressDataVec_hitReq_1_38;
  assign compressDataVec_hitReq_1_38 = _GEN_1243;
  wire          compressDataVec_hitReq_1_166;
  assign compressDataVec_hitReq_1_166 = _GEN_1243;
  wire          _GEN_1244 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h26;
  wire          compressDataVec_hitReq_2_38;
  assign compressDataVec_hitReq_2_38 = _GEN_1244;
  wire          compressDataVec_hitReq_2_166;
  assign compressDataVec_hitReq_2_166 = _GEN_1244;
  wire          _GEN_1245 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h26;
  wire          compressDataVec_hitReq_3_38;
  assign compressDataVec_hitReq_3_38 = _GEN_1245;
  wire          compressDataVec_hitReq_3_166;
  assign compressDataVec_hitReq_3_166 = _GEN_1245;
  wire          _GEN_1246 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h26;
  wire          compressDataVec_hitReq_4_38;
  assign compressDataVec_hitReq_4_38 = _GEN_1246;
  wire          compressDataVec_hitReq_4_166;
  assign compressDataVec_hitReq_4_166 = _GEN_1246;
  wire          _GEN_1247 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h26;
  wire          compressDataVec_hitReq_5_38;
  assign compressDataVec_hitReq_5_38 = _GEN_1247;
  wire          compressDataVec_hitReq_5_166;
  assign compressDataVec_hitReq_5_166 = _GEN_1247;
  wire          _GEN_1248 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h26;
  wire          compressDataVec_hitReq_6_38;
  assign compressDataVec_hitReq_6_38 = _GEN_1248;
  wire          compressDataVec_hitReq_6_166;
  assign compressDataVec_hitReq_6_166 = _GEN_1248;
  wire          _GEN_1249 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h26;
  wire          compressDataVec_hitReq_7_38;
  assign compressDataVec_hitReq_7_38 = _GEN_1249;
  wire          compressDataVec_hitReq_7_166;
  assign compressDataVec_hitReq_7_166 = _GEN_1249;
  wire          _GEN_1250 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h26;
  wire          compressDataVec_hitReq_8_38;
  assign compressDataVec_hitReq_8_38 = _GEN_1250;
  wire          compressDataVec_hitReq_8_166;
  assign compressDataVec_hitReq_8_166 = _GEN_1250;
  wire          _GEN_1251 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h26;
  wire          compressDataVec_hitReq_9_38;
  assign compressDataVec_hitReq_9_38 = _GEN_1251;
  wire          compressDataVec_hitReq_9_166;
  assign compressDataVec_hitReq_9_166 = _GEN_1251;
  wire          _GEN_1252 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h26;
  wire          compressDataVec_hitReq_10_38;
  assign compressDataVec_hitReq_10_38 = _GEN_1252;
  wire          compressDataVec_hitReq_10_166;
  assign compressDataVec_hitReq_10_166 = _GEN_1252;
  wire          _GEN_1253 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h26;
  wire          compressDataVec_hitReq_11_38;
  assign compressDataVec_hitReq_11_38 = _GEN_1253;
  wire          compressDataVec_hitReq_11_166;
  assign compressDataVec_hitReq_11_166 = _GEN_1253;
  wire          _GEN_1254 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h26;
  wire          compressDataVec_hitReq_12_38;
  assign compressDataVec_hitReq_12_38 = _GEN_1254;
  wire          compressDataVec_hitReq_12_166;
  assign compressDataVec_hitReq_12_166 = _GEN_1254;
  wire          _GEN_1255 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h26;
  wire          compressDataVec_hitReq_13_38;
  assign compressDataVec_hitReq_13_38 = _GEN_1255;
  wire          compressDataVec_hitReq_13_166;
  assign compressDataVec_hitReq_13_166 = _GEN_1255;
  wire          _GEN_1256 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h26;
  wire          compressDataVec_hitReq_14_38;
  assign compressDataVec_hitReq_14_38 = _GEN_1256;
  wire          compressDataVec_hitReq_14_166;
  assign compressDataVec_hitReq_14_166 = _GEN_1256;
  wire          _GEN_1257 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h26;
  wire          compressDataVec_hitReq_15_38;
  assign compressDataVec_hitReq_15_38 = _GEN_1257;
  wire          compressDataVec_hitReq_15_166;
  assign compressDataVec_hitReq_15_166 = _GEN_1257;
  wire          _GEN_1258 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h26;
  wire          compressDataVec_hitReq_16_38;
  assign compressDataVec_hitReq_16_38 = _GEN_1258;
  wire          compressDataVec_hitReq_16_166;
  assign compressDataVec_hitReq_16_166 = _GEN_1258;
  wire          _GEN_1259 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h26;
  wire          compressDataVec_hitReq_17_38;
  assign compressDataVec_hitReq_17_38 = _GEN_1259;
  wire          compressDataVec_hitReq_17_166;
  assign compressDataVec_hitReq_17_166 = _GEN_1259;
  wire          _GEN_1260 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h26;
  wire          compressDataVec_hitReq_18_38;
  assign compressDataVec_hitReq_18_38 = _GEN_1260;
  wire          compressDataVec_hitReq_18_166;
  assign compressDataVec_hitReq_18_166 = _GEN_1260;
  wire          _GEN_1261 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h26;
  wire          compressDataVec_hitReq_19_38;
  assign compressDataVec_hitReq_19_38 = _GEN_1261;
  wire          compressDataVec_hitReq_19_166;
  assign compressDataVec_hitReq_19_166 = _GEN_1261;
  wire          _GEN_1262 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h26;
  wire          compressDataVec_hitReq_20_38;
  assign compressDataVec_hitReq_20_38 = _GEN_1262;
  wire          compressDataVec_hitReq_20_166;
  assign compressDataVec_hitReq_20_166 = _GEN_1262;
  wire          _GEN_1263 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h26;
  wire          compressDataVec_hitReq_21_38;
  assign compressDataVec_hitReq_21_38 = _GEN_1263;
  wire          compressDataVec_hitReq_21_166;
  assign compressDataVec_hitReq_21_166 = _GEN_1263;
  wire          _GEN_1264 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h26;
  wire          compressDataVec_hitReq_22_38;
  assign compressDataVec_hitReq_22_38 = _GEN_1264;
  wire          compressDataVec_hitReq_22_166;
  assign compressDataVec_hitReq_22_166 = _GEN_1264;
  wire          _GEN_1265 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h26;
  wire          compressDataVec_hitReq_23_38;
  assign compressDataVec_hitReq_23_38 = _GEN_1265;
  wire          compressDataVec_hitReq_23_166;
  assign compressDataVec_hitReq_23_166 = _GEN_1265;
  wire          _GEN_1266 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h26;
  wire          compressDataVec_hitReq_24_38;
  assign compressDataVec_hitReq_24_38 = _GEN_1266;
  wire          compressDataVec_hitReq_24_166;
  assign compressDataVec_hitReq_24_166 = _GEN_1266;
  wire          _GEN_1267 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h26;
  wire          compressDataVec_hitReq_25_38;
  assign compressDataVec_hitReq_25_38 = _GEN_1267;
  wire          compressDataVec_hitReq_25_166;
  assign compressDataVec_hitReq_25_166 = _GEN_1267;
  wire          _GEN_1268 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h26;
  wire          compressDataVec_hitReq_26_38;
  assign compressDataVec_hitReq_26_38 = _GEN_1268;
  wire          compressDataVec_hitReq_26_166;
  assign compressDataVec_hitReq_26_166 = _GEN_1268;
  wire          _GEN_1269 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h26;
  wire          compressDataVec_hitReq_27_38;
  assign compressDataVec_hitReq_27_38 = _GEN_1269;
  wire          compressDataVec_hitReq_27_166;
  assign compressDataVec_hitReq_27_166 = _GEN_1269;
  wire          _GEN_1270 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h26;
  wire          compressDataVec_hitReq_28_38;
  assign compressDataVec_hitReq_28_38 = _GEN_1270;
  wire          compressDataVec_hitReq_28_166;
  assign compressDataVec_hitReq_28_166 = _GEN_1270;
  wire          _GEN_1271 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h26;
  wire          compressDataVec_hitReq_29_38;
  assign compressDataVec_hitReq_29_38 = _GEN_1271;
  wire          compressDataVec_hitReq_29_166;
  assign compressDataVec_hitReq_29_166 = _GEN_1271;
  wire          _GEN_1272 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h26;
  wire          compressDataVec_hitReq_30_38;
  assign compressDataVec_hitReq_30_38 = _GEN_1272;
  wire          compressDataVec_hitReq_30_166;
  assign compressDataVec_hitReq_30_166 = _GEN_1272;
  wire          _GEN_1273 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h26;
  wire          compressDataVec_hitReq_31_38;
  assign compressDataVec_hitReq_31_38 = _GEN_1273;
  wire          compressDataVec_hitReq_31_166;
  assign compressDataVec_hitReq_31_166 = _GEN_1273;
  wire          compressDataVec_hitReq_32_38 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h26;
  wire          compressDataVec_hitReq_33_38 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h26;
  wire          compressDataVec_hitReq_34_38 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h26;
  wire          compressDataVec_hitReq_35_38 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h26;
  wire          compressDataVec_hitReq_36_38 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h26;
  wire          compressDataVec_hitReq_37_38 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h26;
  wire          compressDataVec_hitReq_38_38 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h26;
  wire          compressDataVec_hitReq_39_38 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h26;
  wire          compressDataVec_hitReq_40_38 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h26;
  wire          compressDataVec_hitReq_41_38 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h26;
  wire          compressDataVec_hitReq_42_38 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h26;
  wire          compressDataVec_hitReq_43_38 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h26;
  wire          compressDataVec_hitReq_44_38 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h26;
  wire          compressDataVec_hitReq_45_38 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h26;
  wire          compressDataVec_hitReq_46_38 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h26;
  wire          compressDataVec_hitReq_47_38 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h26;
  wire          compressDataVec_hitReq_48_38 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h26;
  wire          compressDataVec_hitReq_49_38 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h26;
  wire          compressDataVec_hitReq_50_38 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h26;
  wire          compressDataVec_hitReq_51_38 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h26;
  wire          compressDataVec_hitReq_52_38 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h26;
  wire          compressDataVec_hitReq_53_38 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h26;
  wire          compressDataVec_hitReq_54_38 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h26;
  wire          compressDataVec_hitReq_55_38 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h26;
  wire          compressDataVec_hitReq_56_38 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h26;
  wire          compressDataVec_hitReq_57_38 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h26;
  wire          compressDataVec_hitReq_58_38 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h26;
  wire          compressDataVec_hitReq_59_38 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h26;
  wire          compressDataVec_hitReq_60_38 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h26;
  wire          compressDataVec_hitReq_61_38 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h26;
  wire          compressDataVec_hitReq_62_38 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h26;
  wire          compressDataVec_hitReq_63_38 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h26;
  wire [7:0]    compressDataVec_selectReqData_38 =
    (compressDataVec_hitReq_0_38 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_38 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_38 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_38 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_38 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_38 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_38 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_38 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_38 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_38 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_38 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_38 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_38 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_38 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_38 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_38 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_38 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_38 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_38 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_38 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_38 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_38 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_38 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_38 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_38 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_38 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_38 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_38 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_38 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_38 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_38 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_38 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_38 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_38 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_38 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_38 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_38 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_38 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_38 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_38 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_38 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_38 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_38 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_38 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_38 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_38 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_38 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_38 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_38 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_38 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_38 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_38 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_38 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_38 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_38 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_38 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_38 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_38 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_38 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_38 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_38 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_38 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_38 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_38 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_38 = tailCount > 6'h26;
  wire          _GEN_1274 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h27;
  wire          compressDataVec_hitReq_0_39;
  assign compressDataVec_hitReq_0_39 = _GEN_1274;
  wire          compressDataVec_hitReq_0_167;
  assign compressDataVec_hitReq_0_167 = _GEN_1274;
  wire          _GEN_1275 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h27;
  wire          compressDataVec_hitReq_1_39;
  assign compressDataVec_hitReq_1_39 = _GEN_1275;
  wire          compressDataVec_hitReq_1_167;
  assign compressDataVec_hitReq_1_167 = _GEN_1275;
  wire          _GEN_1276 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h27;
  wire          compressDataVec_hitReq_2_39;
  assign compressDataVec_hitReq_2_39 = _GEN_1276;
  wire          compressDataVec_hitReq_2_167;
  assign compressDataVec_hitReq_2_167 = _GEN_1276;
  wire          _GEN_1277 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h27;
  wire          compressDataVec_hitReq_3_39;
  assign compressDataVec_hitReq_3_39 = _GEN_1277;
  wire          compressDataVec_hitReq_3_167;
  assign compressDataVec_hitReq_3_167 = _GEN_1277;
  wire          _GEN_1278 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h27;
  wire          compressDataVec_hitReq_4_39;
  assign compressDataVec_hitReq_4_39 = _GEN_1278;
  wire          compressDataVec_hitReq_4_167;
  assign compressDataVec_hitReq_4_167 = _GEN_1278;
  wire          _GEN_1279 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h27;
  wire          compressDataVec_hitReq_5_39;
  assign compressDataVec_hitReq_5_39 = _GEN_1279;
  wire          compressDataVec_hitReq_5_167;
  assign compressDataVec_hitReq_5_167 = _GEN_1279;
  wire          _GEN_1280 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h27;
  wire          compressDataVec_hitReq_6_39;
  assign compressDataVec_hitReq_6_39 = _GEN_1280;
  wire          compressDataVec_hitReq_6_167;
  assign compressDataVec_hitReq_6_167 = _GEN_1280;
  wire          _GEN_1281 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h27;
  wire          compressDataVec_hitReq_7_39;
  assign compressDataVec_hitReq_7_39 = _GEN_1281;
  wire          compressDataVec_hitReq_7_167;
  assign compressDataVec_hitReq_7_167 = _GEN_1281;
  wire          _GEN_1282 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h27;
  wire          compressDataVec_hitReq_8_39;
  assign compressDataVec_hitReq_8_39 = _GEN_1282;
  wire          compressDataVec_hitReq_8_167;
  assign compressDataVec_hitReq_8_167 = _GEN_1282;
  wire          _GEN_1283 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h27;
  wire          compressDataVec_hitReq_9_39;
  assign compressDataVec_hitReq_9_39 = _GEN_1283;
  wire          compressDataVec_hitReq_9_167;
  assign compressDataVec_hitReq_9_167 = _GEN_1283;
  wire          _GEN_1284 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h27;
  wire          compressDataVec_hitReq_10_39;
  assign compressDataVec_hitReq_10_39 = _GEN_1284;
  wire          compressDataVec_hitReq_10_167;
  assign compressDataVec_hitReq_10_167 = _GEN_1284;
  wire          _GEN_1285 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h27;
  wire          compressDataVec_hitReq_11_39;
  assign compressDataVec_hitReq_11_39 = _GEN_1285;
  wire          compressDataVec_hitReq_11_167;
  assign compressDataVec_hitReq_11_167 = _GEN_1285;
  wire          _GEN_1286 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h27;
  wire          compressDataVec_hitReq_12_39;
  assign compressDataVec_hitReq_12_39 = _GEN_1286;
  wire          compressDataVec_hitReq_12_167;
  assign compressDataVec_hitReq_12_167 = _GEN_1286;
  wire          _GEN_1287 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h27;
  wire          compressDataVec_hitReq_13_39;
  assign compressDataVec_hitReq_13_39 = _GEN_1287;
  wire          compressDataVec_hitReq_13_167;
  assign compressDataVec_hitReq_13_167 = _GEN_1287;
  wire          _GEN_1288 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h27;
  wire          compressDataVec_hitReq_14_39;
  assign compressDataVec_hitReq_14_39 = _GEN_1288;
  wire          compressDataVec_hitReq_14_167;
  assign compressDataVec_hitReq_14_167 = _GEN_1288;
  wire          _GEN_1289 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h27;
  wire          compressDataVec_hitReq_15_39;
  assign compressDataVec_hitReq_15_39 = _GEN_1289;
  wire          compressDataVec_hitReq_15_167;
  assign compressDataVec_hitReq_15_167 = _GEN_1289;
  wire          _GEN_1290 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h27;
  wire          compressDataVec_hitReq_16_39;
  assign compressDataVec_hitReq_16_39 = _GEN_1290;
  wire          compressDataVec_hitReq_16_167;
  assign compressDataVec_hitReq_16_167 = _GEN_1290;
  wire          _GEN_1291 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h27;
  wire          compressDataVec_hitReq_17_39;
  assign compressDataVec_hitReq_17_39 = _GEN_1291;
  wire          compressDataVec_hitReq_17_167;
  assign compressDataVec_hitReq_17_167 = _GEN_1291;
  wire          _GEN_1292 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h27;
  wire          compressDataVec_hitReq_18_39;
  assign compressDataVec_hitReq_18_39 = _GEN_1292;
  wire          compressDataVec_hitReq_18_167;
  assign compressDataVec_hitReq_18_167 = _GEN_1292;
  wire          _GEN_1293 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h27;
  wire          compressDataVec_hitReq_19_39;
  assign compressDataVec_hitReq_19_39 = _GEN_1293;
  wire          compressDataVec_hitReq_19_167;
  assign compressDataVec_hitReq_19_167 = _GEN_1293;
  wire          _GEN_1294 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h27;
  wire          compressDataVec_hitReq_20_39;
  assign compressDataVec_hitReq_20_39 = _GEN_1294;
  wire          compressDataVec_hitReq_20_167;
  assign compressDataVec_hitReq_20_167 = _GEN_1294;
  wire          _GEN_1295 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h27;
  wire          compressDataVec_hitReq_21_39;
  assign compressDataVec_hitReq_21_39 = _GEN_1295;
  wire          compressDataVec_hitReq_21_167;
  assign compressDataVec_hitReq_21_167 = _GEN_1295;
  wire          _GEN_1296 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h27;
  wire          compressDataVec_hitReq_22_39;
  assign compressDataVec_hitReq_22_39 = _GEN_1296;
  wire          compressDataVec_hitReq_22_167;
  assign compressDataVec_hitReq_22_167 = _GEN_1296;
  wire          _GEN_1297 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h27;
  wire          compressDataVec_hitReq_23_39;
  assign compressDataVec_hitReq_23_39 = _GEN_1297;
  wire          compressDataVec_hitReq_23_167;
  assign compressDataVec_hitReq_23_167 = _GEN_1297;
  wire          _GEN_1298 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h27;
  wire          compressDataVec_hitReq_24_39;
  assign compressDataVec_hitReq_24_39 = _GEN_1298;
  wire          compressDataVec_hitReq_24_167;
  assign compressDataVec_hitReq_24_167 = _GEN_1298;
  wire          _GEN_1299 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h27;
  wire          compressDataVec_hitReq_25_39;
  assign compressDataVec_hitReq_25_39 = _GEN_1299;
  wire          compressDataVec_hitReq_25_167;
  assign compressDataVec_hitReq_25_167 = _GEN_1299;
  wire          _GEN_1300 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h27;
  wire          compressDataVec_hitReq_26_39;
  assign compressDataVec_hitReq_26_39 = _GEN_1300;
  wire          compressDataVec_hitReq_26_167;
  assign compressDataVec_hitReq_26_167 = _GEN_1300;
  wire          _GEN_1301 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h27;
  wire          compressDataVec_hitReq_27_39;
  assign compressDataVec_hitReq_27_39 = _GEN_1301;
  wire          compressDataVec_hitReq_27_167;
  assign compressDataVec_hitReq_27_167 = _GEN_1301;
  wire          _GEN_1302 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h27;
  wire          compressDataVec_hitReq_28_39;
  assign compressDataVec_hitReq_28_39 = _GEN_1302;
  wire          compressDataVec_hitReq_28_167;
  assign compressDataVec_hitReq_28_167 = _GEN_1302;
  wire          _GEN_1303 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h27;
  wire          compressDataVec_hitReq_29_39;
  assign compressDataVec_hitReq_29_39 = _GEN_1303;
  wire          compressDataVec_hitReq_29_167;
  assign compressDataVec_hitReq_29_167 = _GEN_1303;
  wire          _GEN_1304 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h27;
  wire          compressDataVec_hitReq_30_39;
  assign compressDataVec_hitReq_30_39 = _GEN_1304;
  wire          compressDataVec_hitReq_30_167;
  assign compressDataVec_hitReq_30_167 = _GEN_1304;
  wire          _GEN_1305 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h27;
  wire          compressDataVec_hitReq_31_39;
  assign compressDataVec_hitReq_31_39 = _GEN_1305;
  wire          compressDataVec_hitReq_31_167;
  assign compressDataVec_hitReq_31_167 = _GEN_1305;
  wire          compressDataVec_hitReq_32_39 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h27;
  wire          compressDataVec_hitReq_33_39 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h27;
  wire          compressDataVec_hitReq_34_39 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h27;
  wire          compressDataVec_hitReq_35_39 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h27;
  wire          compressDataVec_hitReq_36_39 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h27;
  wire          compressDataVec_hitReq_37_39 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h27;
  wire          compressDataVec_hitReq_38_39 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h27;
  wire          compressDataVec_hitReq_39_39 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h27;
  wire          compressDataVec_hitReq_40_39 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h27;
  wire          compressDataVec_hitReq_41_39 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h27;
  wire          compressDataVec_hitReq_42_39 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h27;
  wire          compressDataVec_hitReq_43_39 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h27;
  wire          compressDataVec_hitReq_44_39 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h27;
  wire          compressDataVec_hitReq_45_39 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h27;
  wire          compressDataVec_hitReq_46_39 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h27;
  wire          compressDataVec_hitReq_47_39 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h27;
  wire          compressDataVec_hitReq_48_39 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h27;
  wire          compressDataVec_hitReq_49_39 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h27;
  wire          compressDataVec_hitReq_50_39 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h27;
  wire          compressDataVec_hitReq_51_39 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h27;
  wire          compressDataVec_hitReq_52_39 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h27;
  wire          compressDataVec_hitReq_53_39 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h27;
  wire          compressDataVec_hitReq_54_39 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h27;
  wire          compressDataVec_hitReq_55_39 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h27;
  wire          compressDataVec_hitReq_56_39 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h27;
  wire          compressDataVec_hitReq_57_39 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h27;
  wire          compressDataVec_hitReq_58_39 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h27;
  wire          compressDataVec_hitReq_59_39 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h27;
  wire          compressDataVec_hitReq_60_39 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h27;
  wire          compressDataVec_hitReq_61_39 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h27;
  wire          compressDataVec_hitReq_62_39 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h27;
  wire          compressDataVec_hitReq_63_39 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h27;
  wire [7:0]    compressDataVec_selectReqData_39 =
    (compressDataVec_hitReq_0_39 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_39 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_39 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_39 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_39 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_39 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_39 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_39 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_39 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_39 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_39 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_39 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_39 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_39 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_39 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_39 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_39 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_39 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_39 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_39 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_39 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_39 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_39 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_39 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_39 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_39 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_39 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_39 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_39 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_39 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_39 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_39 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_39 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_39 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_39 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_39 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_39 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_39 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_39 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_39 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_39 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_39 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_39 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_39 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_39 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_39 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_39 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_39 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_39 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_39 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_39 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_39 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_39 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_39 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_39 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_39 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_39 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_39 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_39 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_39 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_39 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_39 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_39 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_39 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_39 = tailCount > 6'h27;
  wire          _GEN_1306 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h28;
  wire          compressDataVec_hitReq_0_40;
  assign compressDataVec_hitReq_0_40 = _GEN_1306;
  wire          compressDataVec_hitReq_0_168;
  assign compressDataVec_hitReq_0_168 = _GEN_1306;
  wire          _GEN_1307 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h28;
  wire          compressDataVec_hitReq_1_40;
  assign compressDataVec_hitReq_1_40 = _GEN_1307;
  wire          compressDataVec_hitReq_1_168;
  assign compressDataVec_hitReq_1_168 = _GEN_1307;
  wire          _GEN_1308 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h28;
  wire          compressDataVec_hitReq_2_40;
  assign compressDataVec_hitReq_2_40 = _GEN_1308;
  wire          compressDataVec_hitReq_2_168;
  assign compressDataVec_hitReq_2_168 = _GEN_1308;
  wire          _GEN_1309 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h28;
  wire          compressDataVec_hitReq_3_40;
  assign compressDataVec_hitReq_3_40 = _GEN_1309;
  wire          compressDataVec_hitReq_3_168;
  assign compressDataVec_hitReq_3_168 = _GEN_1309;
  wire          _GEN_1310 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h28;
  wire          compressDataVec_hitReq_4_40;
  assign compressDataVec_hitReq_4_40 = _GEN_1310;
  wire          compressDataVec_hitReq_4_168;
  assign compressDataVec_hitReq_4_168 = _GEN_1310;
  wire          _GEN_1311 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h28;
  wire          compressDataVec_hitReq_5_40;
  assign compressDataVec_hitReq_5_40 = _GEN_1311;
  wire          compressDataVec_hitReq_5_168;
  assign compressDataVec_hitReq_5_168 = _GEN_1311;
  wire          _GEN_1312 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h28;
  wire          compressDataVec_hitReq_6_40;
  assign compressDataVec_hitReq_6_40 = _GEN_1312;
  wire          compressDataVec_hitReq_6_168;
  assign compressDataVec_hitReq_6_168 = _GEN_1312;
  wire          _GEN_1313 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h28;
  wire          compressDataVec_hitReq_7_40;
  assign compressDataVec_hitReq_7_40 = _GEN_1313;
  wire          compressDataVec_hitReq_7_168;
  assign compressDataVec_hitReq_7_168 = _GEN_1313;
  wire          _GEN_1314 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h28;
  wire          compressDataVec_hitReq_8_40;
  assign compressDataVec_hitReq_8_40 = _GEN_1314;
  wire          compressDataVec_hitReq_8_168;
  assign compressDataVec_hitReq_8_168 = _GEN_1314;
  wire          _GEN_1315 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h28;
  wire          compressDataVec_hitReq_9_40;
  assign compressDataVec_hitReq_9_40 = _GEN_1315;
  wire          compressDataVec_hitReq_9_168;
  assign compressDataVec_hitReq_9_168 = _GEN_1315;
  wire          _GEN_1316 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h28;
  wire          compressDataVec_hitReq_10_40;
  assign compressDataVec_hitReq_10_40 = _GEN_1316;
  wire          compressDataVec_hitReq_10_168;
  assign compressDataVec_hitReq_10_168 = _GEN_1316;
  wire          _GEN_1317 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h28;
  wire          compressDataVec_hitReq_11_40;
  assign compressDataVec_hitReq_11_40 = _GEN_1317;
  wire          compressDataVec_hitReq_11_168;
  assign compressDataVec_hitReq_11_168 = _GEN_1317;
  wire          _GEN_1318 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h28;
  wire          compressDataVec_hitReq_12_40;
  assign compressDataVec_hitReq_12_40 = _GEN_1318;
  wire          compressDataVec_hitReq_12_168;
  assign compressDataVec_hitReq_12_168 = _GEN_1318;
  wire          _GEN_1319 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h28;
  wire          compressDataVec_hitReq_13_40;
  assign compressDataVec_hitReq_13_40 = _GEN_1319;
  wire          compressDataVec_hitReq_13_168;
  assign compressDataVec_hitReq_13_168 = _GEN_1319;
  wire          _GEN_1320 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h28;
  wire          compressDataVec_hitReq_14_40;
  assign compressDataVec_hitReq_14_40 = _GEN_1320;
  wire          compressDataVec_hitReq_14_168;
  assign compressDataVec_hitReq_14_168 = _GEN_1320;
  wire          _GEN_1321 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h28;
  wire          compressDataVec_hitReq_15_40;
  assign compressDataVec_hitReq_15_40 = _GEN_1321;
  wire          compressDataVec_hitReq_15_168;
  assign compressDataVec_hitReq_15_168 = _GEN_1321;
  wire          _GEN_1322 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h28;
  wire          compressDataVec_hitReq_16_40;
  assign compressDataVec_hitReq_16_40 = _GEN_1322;
  wire          compressDataVec_hitReq_16_168;
  assign compressDataVec_hitReq_16_168 = _GEN_1322;
  wire          _GEN_1323 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h28;
  wire          compressDataVec_hitReq_17_40;
  assign compressDataVec_hitReq_17_40 = _GEN_1323;
  wire          compressDataVec_hitReq_17_168;
  assign compressDataVec_hitReq_17_168 = _GEN_1323;
  wire          _GEN_1324 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h28;
  wire          compressDataVec_hitReq_18_40;
  assign compressDataVec_hitReq_18_40 = _GEN_1324;
  wire          compressDataVec_hitReq_18_168;
  assign compressDataVec_hitReq_18_168 = _GEN_1324;
  wire          _GEN_1325 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h28;
  wire          compressDataVec_hitReq_19_40;
  assign compressDataVec_hitReq_19_40 = _GEN_1325;
  wire          compressDataVec_hitReq_19_168;
  assign compressDataVec_hitReq_19_168 = _GEN_1325;
  wire          _GEN_1326 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h28;
  wire          compressDataVec_hitReq_20_40;
  assign compressDataVec_hitReq_20_40 = _GEN_1326;
  wire          compressDataVec_hitReq_20_168;
  assign compressDataVec_hitReq_20_168 = _GEN_1326;
  wire          _GEN_1327 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h28;
  wire          compressDataVec_hitReq_21_40;
  assign compressDataVec_hitReq_21_40 = _GEN_1327;
  wire          compressDataVec_hitReq_21_168;
  assign compressDataVec_hitReq_21_168 = _GEN_1327;
  wire          _GEN_1328 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h28;
  wire          compressDataVec_hitReq_22_40;
  assign compressDataVec_hitReq_22_40 = _GEN_1328;
  wire          compressDataVec_hitReq_22_168;
  assign compressDataVec_hitReq_22_168 = _GEN_1328;
  wire          _GEN_1329 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h28;
  wire          compressDataVec_hitReq_23_40;
  assign compressDataVec_hitReq_23_40 = _GEN_1329;
  wire          compressDataVec_hitReq_23_168;
  assign compressDataVec_hitReq_23_168 = _GEN_1329;
  wire          _GEN_1330 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h28;
  wire          compressDataVec_hitReq_24_40;
  assign compressDataVec_hitReq_24_40 = _GEN_1330;
  wire          compressDataVec_hitReq_24_168;
  assign compressDataVec_hitReq_24_168 = _GEN_1330;
  wire          _GEN_1331 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h28;
  wire          compressDataVec_hitReq_25_40;
  assign compressDataVec_hitReq_25_40 = _GEN_1331;
  wire          compressDataVec_hitReq_25_168;
  assign compressDataVec_hitReq_25_168 = _GEN_1331;
  wire          _GEN_1332 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h28;
  wire          compressDataVec_hitReq_26_40;
  assign compressDataVec_hitReq_26_40 = _GEN_1332;
  wire          compressDataVec_hitReq_26_168;
  assign compressDataVec_hitReq_26_168 = _GEN_1332;
  wire          _GEN_1333 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h28;
  wire          compressDataVec_hitReq_27_40;
  assign compressDataVec_hitReq_27_40 = _GEN_1333;
  wire          compressDataVec_hitReq_27_168;
  assign compressDataVec_hitReq_27_168 = _GEN_1333;
  wire          _GEN_1334 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h28;
  wire          compressDataVec_hitReq_28_40;
  assign compressDataVec_hitReq_28_40 = _GEN_1334;
  wire          compressDataVec_hitReq_28_168;
  assign compressDataVec_hitReq_28_168 = _GEN_1334;
  wire          _GEN_1335 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h28;
  wire          compressDataVec_hitReq_29_40;
  assign compressDataVec_hitReq_29_40 = _GEN_1335;
  wire          compressDataVec_hitReq_29_168;
  assign compressDataVec_hitReq_29_168 = _GEN_1335;
  wire          _GEN_1336 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h28;
  wire          compressDataVec_hitReq_30_40;
  assign compressDataVec_hitReq_30_40 = _GEN_1336;
  wire          compressDataVec_hitReq_30_168;
  assign compressDataVec_hitReq_30_168 = _GEN_1336;
  wire          _GEN_1337 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h28;
  wire          compressDataVec_hitReq_31_40;
  assign compressDataVec_hitReq_31_40 = _GEN_1337;
  wire          compressDataVec_hitReq_31_168;
  assign compressDataVec_hitReq_31_168 = _GEN_1337;
  wire          compressDataVec_hitReq_32_40 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h28;
  wire          compressDataVec_hitReq_33_40 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h28;
  wire          compressDataVec_hitReq_34_40 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h28;
  wire          compressDataVec_hitReq_35_40 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h28;
  wire          compressDataVec_hitReq_36_40 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h28;
  wire          compressDataVec_hitReq_37_40 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h28;
  wire          compressDataVec_hitReq_38_40 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h28;
  wire          compressDataVec_hitReq_39_40 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h28;
  wire          compressDataVec_hitReq_40_40 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h28;
  wire          compressDataVec_hitReq_41_40 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h28;
  wire          compressDataVec_hitReq_42_40 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h28;
  wire          compressDataVec_hitReq_43_40 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h28;
  wire          compressDataVec_hitReq_44_40 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h28;
  wire          compressDataVec_hitReq_45_40 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h28;
  wire          compressDataVec_hitReq_46_40 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h28;
  wire          compressDataVec_hitReq_47_40 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h28;
  wire          compressDataVec_hitReq_48_40 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h28;
  wire          compressDataVec_hitReq_49_40 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h28;
  wire          compressDataVec_hitReq_50_40 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h28;
  wire          compressDataVec_hitReq_51_40 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h28;
  wire          compressDataVec_hitReq_52_40 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h28;
  wire          compressDataVec_hitReq_53_40 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h28;
  wire          compressDataVec_hitReq_54_40 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h28;
  wire          compressDataVec_hitReq_55_40 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h28;
  wire          compressDataVec_hitReq_56_40 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h28;
  wire          compressDataVec_hitReq_57_40 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h28;
  wire          compressDataVec_hitReq_58_40 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h28;
  wire          compressDataVec_hitReq_59_40 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h28;
  wire          compressDataVec_hitReq_60_40 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h28;
  wire          compressDataVec_hitReq_61_40 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h28;
  wire          compressDataVec_hitReq_62_40 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h28;
  wire          compressDataVec_hitReq_63_40 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h28;
  wire [7:0]    compressDataVec_selectReqData_40 =
    (compressDataVec_hitReq_0_40 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_40 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_40 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_40 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_40 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_40 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_40 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_40 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_40 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_40 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_40 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_40 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_40 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_40 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_40 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_40 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_40 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_40 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_40 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_40 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_40 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_40 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_40 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_40 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_40 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_40 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_40 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_40 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_40 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_40 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_40 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_40 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_40 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_40 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_40 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_40 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_40 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_40 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_40 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_40 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_40 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_40 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_40 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_40 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_40 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_40 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_40 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_40 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_40 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_40 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_40 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_40 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_40 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_40 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_40 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_40 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_40 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_40 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_40 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_40 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_40 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_40 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_40 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_40 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_40 = tailCount > 6'h28;
  wire          _GEN_1338 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h29;
  wire          compressDataVec_hitReq_0_41;
  assign compressDataVec_hitReq_0_41 = _GEN_1338;
  wire          compressDataVec_hitReq_0_169;
  assign compressDataVec_hitReq_0_169 = _GEN_1338;
  wire          _GEN_1339 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h29;
  wire          compressDataVec_hitReq_1_41;
  assign compressDataVec_hitReq_1_41 = _GEN_1339;
  wire          compressDataVec_hitReq_1_169;
  assign compressDataVec_hitReq_1_169 = _GEN_1339;
  wire          _GEN_1340 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h29;
  wire          compressDataVec_hitReq_2_41;
  assign compressDataVec_hitReq_2_41 = _GEN_1340;
  wire          compressDataVec_hitReq_2_169;
  assign compressDataVec_hitReq_2_169 = _GEN_1340;
  wire          _GEN_1341 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h29;
  wire          compressDataVec_hitReq_3_41;
  assign compressDataVec_hitReq_3_41 = _GEN_1341;
  wire          compressDataVec_hitReq_3_169;
  assign compressDataVec_hitReq_3_169 = _GEN_1341;
  wire          _GEN_1342 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h29;
  wire          compressDataVec_hitReq_4_41;
  assign compressDataVec_hitReq_4_41 = _GEN_1342;
  wire          compressDataVec_hitReq_4_169;
  assign compressDataVec_hitReq_4_169 = _GEN_1342;
  wire          _GEN_1343 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h29;
  wire          compressDataVec_hitReq_5_41;
  assign compressDataVec_hitReq_5_41 = _GEN_1343;
  wire          compressDataVec_hitReq_5_169;
  assign compressDataVec_hitReq_5_169 = _GEN_1343;
  wire          _GEN_1344 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h29;
  wire          compressDataVec_hitReq_6_41;
  assign compressDataVec_hitReq_6_41 = _GEN_1344;
  wire          compressDataVec_hitReq_6_169;
  assign compressDataVec_hitReq_6_169 = _GEN_1344;
  wire          _GEN_1345 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h29;
  wire          compressDataVec_hitReq_7_41;
  assign compressDataVec_hitReq_7_41 = _GEN_1345;
  wire          compressDataVec_hitReq_7_169;
  assign compressDataVec_hitReq_7_169 = _GEN_1345;
  wire          _GEN_1346 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h29;
  wire          compressDataVec_hitReq_8_41;
  assign compressDataVec_hitReq_8_41 = _GEN_1346;
  wire          compressDataVec_hitReq_8_169;
  assign compressDataVec_hitReq_8_169 = _GEN_1346;
  wire          _GEN_1347 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h29;
  wire          compressDataVec_hitReq_9_41;
  assign compressDataVec_hitReq_9_41 = _GEN_1347;
  wire          compressDataVec_hitReq_9_169;
  assign compressDataVec_hitReq_9_169 = _GEN_1347;
  wire          _GEN_1348 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h29;
  wire          compressDataVec_hitReq_10_41;
  assign compressDataVec_hitReq_10_41 = _GEN_1348;
  wire          compressDataVec_hitReq_10_169;
  assign compressDataVec_hitReq_10_169 = _GEN_1348;
  wire          _GEN_1349 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h29;
  wire          compressDataVec_hitReq_11_41;
  assign compressDataVec_hitReq_11_41 = _GEN_1349;
  wire          compressDataVec_hitReq_11_169;
  assign compressDataVec_hitReq_11_169 = _GEN_1349;
  wire          _GEN_1350 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h29;
  wire          compressDataVec_hitReq_12_41;
  assign compressDataVec_hitReq_12_41 = _GEN_1350;
  wire          compressDataVec_hitReq_12_169;
  assign compressDataVec_hitReq_12_169 = _GEN_1350;
  wire          _GEN_1351 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h29;
  wire          compressDataVec_hitReq_13_41;
  assign compressDataVec_hitReq_13_41 = _GEN_1351;
  wire          compressDataVec_hitReq_13_169;
  assign compressDataVec_hitReq_13_169 = _GEN_1351;
  wire          _GEN_1352 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h29;
  wire          compressDataVec_hitReq_14_41;
  assign compressDataVec_hitReq_14_41 = _GEN_1352;
  wire          compressDataVec_hitReq_14_169;
  assign compressDataVec_hitReq_14_169 = _GEN_1352;
  wire          _GEN_1353 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h29;
  wire          compressDataVec_hitReq_15_41;
  assign compressDataVec_hitReq_15_41 = _GEN_1353;
  wire          compressDataVec_hitReq_15_169;
  assign compressDataVec_hitReq_15_169 = _GEN_1353;
  wire          _GEN_1354 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h29;
  wire          compressDataVec_hitReq_16_41;
  assign compressDataVec_hitReq_16_41 = _GEN_1354;
  wire          compressDataVec_hitReq_16_169;
  assign compressDataVec_hitReq_16_169 = _GEN_1354;
  wire          _GEN_1355 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h29;
  wire          compressDataVec_hitReq_17_41;
  assign compressDataVec_hitReq_17_41 = _GEN_1355;
  wire          compressDataVec_hitReq_17_169;
  assign compressDataVec_hitReq_17_169 = _GEN_1355;
  wire          _GEN_1356 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h29;
  wire          compressDataVec_hitReq_18_41;
  assign compressDataVec_hitReq_18_41 = _GEN_1356;
  wire          compressDataVec_hitReq_18_169;
  assign compressDataVec_hitReq_18_169 = _GEN_1356;
  wire          _GEN_1357 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h29;
  wire          compressDataVec_hitReq_19_41;
  assign compressDataVec_hitReq_19_41 = _GEN_1357;
  wire          compressDataVec_hitReq_19_169;
  assign compressDataVec_hitReq_19_169 = _GEN_1357;
  wire          _GEN_1358 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h29;
  wire          compressDataVec_hitReq_20_41;
  assign compressDataVec_hitReq_20_41 = _GEN_1358;
  wire          compressDataVec_hitReq_20_169;
  assign compressDataVec_hitReq_20_169 = _GEN_1358;
  wire          _GEN_1359 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h29;
  wire          compressDataVec_hitReq_21_41;
  assign compressDataVec_hitReq_21_41 = _GEN_1359;
  wire          compressDataVec_hitReq_21_169;
  assign compressDataVec_hitReq_21_169 = _GEN_1359;
  wire          _GEN_1360 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h29;
  wire          compressDataVec_hitReq_22_41;
  assign compressDataVec_hitReq_22_41 = _GEN_1360;
  wire          compressDataVec_hitReq_22_169;
  assign compressDataVec_hitReq_22_169 = _GEN_1360;
  wire          _GEN_1361 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h29;
  wire          compressDataVec_hitReq_23_41;
  assign compressDataVec_hitReq_23_41 = _GEN_1361;
  wire          compressDataVec_hitReq_23_169;
  assign compressDataVec_hitReq_23_169 = _GEN_1361;
  wire          _GEN_1362 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h29;
  wire          compressDataVec_hitReq_24_41;
  assign compressDataVec_hitReq_24_41 = _GEN_1362;
  wire          compressDataVec_hitReq_24_169;
  assign compressDataVec_hitReq_24_169 = _GEN_1362;
  wire          _GEN_1363 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h29;
  wire          compressDataVec_hitReq_25_41;
  assign compressDataVec_hitReq_25_41 = _GEN_1363;
  wire          compressDataVec_hitReq_25_169;
  assign compressDataVec_hitReq_25_169 = _GEN_1363;
  wire          _GEN_1364 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h29;
  wire          compressDataVec_hitReq_26_41;
  assign compressDataVec_hitReq_26_41 = _GEN_1364;
  wire          compressDataVec_hitReq_26_169;
  assign compressDataVec_hitReq_26_169 = _GEN_1364;
  wire          _GEN_1365 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h29;
  wire          compressDataVec_hitReq_27_41;
  assign compressDataVec_hitReq_27_41 = _GEN_1365;
  wire          compressDataVec_hitReq_27_169;
  assign compressDataVec_hitReq_27_169 = _GEN_1365;
  wire          _GEN_1366 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h29;
  wire          compressDataVec_hitReq_28_41;
  assign compressDataVec_hitReq_28_41 = _GEN_1366;
  wire          compressDataVec_hitReq_28_169;
  assign compressDataVec_hitReq_28_169 = _GEN_1366;
  wire          _GEN_1367 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h29;
  wire          compressDataVec_hitReq_29_41;
  assign compressDataVec_hitReq_29_41 = _GEN_1367;
  wire          compressDataVec_hitReq_29_169;
  assign compressDataVec_hitReq_29_169 = _GEN_1367;
  wire          _GEN_1368 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h29;
  wire          compressDataVec_hitReq_30_41;
  assign compressDataVec_hitReq_30_41 = _GEN_1368;
  wire          compressDataVec_hitReq_30_169;
  assign compressDataVec_hitReq_30_169 = _GEN_1368;
  wire          _GEN_1369 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h29;
  wire          compressDataVec_hitReq_31_41;
  assign compressDataVec_hitReq_31_41 = _GEN_1369;
  wire          compressDataVec_hitReq_31_169;
  assign compressDataVec_hitReq_31_169 = _GEN_1369;
  wire          compressDataVec_hitReq_32_41 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h29;
  wire          compressDataVec_hitReq_33_41 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h29;
  wire          compressDataVec_hitReq_34_41 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h29;
  wire          compressDataVec_hitReq_35_41 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h29;
  wire          compressDataVec_hitReq_36_41 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h29;
  wire          compressDataVec_hitReq_37_41 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h29;
  wire          compressDataVec_hitReq_38_41 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h29;
  wire          compressDataVec_hitReq_39_41 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h29;
  wire          compressDataVec_hitReq_40_41 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h29;
  wire          compressDataVec_hitReq_41_41 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h29;
  wire          compressDataVec_hitReq_42_41 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h29;
  wire          compressDataVec_hitReq_43_41 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h29;
  wire          compressDataVec_hitReq_44_41 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h29;
  wire          compressDataVec_hitReq_45_41 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h29;
  wire          compressDataVec_hitReq_46_41 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h29;
  wire          compressDataVec_hitReq_47_41 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h29;
  wire          compressDataVec_hitReq_48_41 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h29;
  wire          compressDataVec_hitReq_49_41 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h29;
  wire          compressDataVec_hitReq_50_41 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h29;
  wire          compressDataVec_hitReq_51_41 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h29;
  wire          compressDataVec_hitReq_52_41 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h29;
  wire          compressDataVec_hitReq_53_41 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h29;
  wire          compressDataVec_hitReq_54_41 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h29;
  wire          compressDataVec_hitReq_55_41 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h29;
  wire          compressDataVec_hitReq_56_41 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h29;
  wire          compressDataVec_hitReq_57_41 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h29;
  wire          compressDataVec_hitReq_58_41 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h29;
  wire          compressDataVec_hitReq_59_41 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h29;
  wire          compressDataVec_hitReq_60_41 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h29;
  wire          compressDataVec_hitReq_61_41 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h29;
  wire          compressDataVec_hitReq_62_41 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h29;
  wire          compressDataVec_hitReq_63_41 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h29;
  wire [7:0]    compressDataVec_selectReqData_41 =
    (compressDataVec_hitReq_0_41 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_41 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_41 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_41 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_41 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_41 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_41 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_41 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_41 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_41 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_41 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_41 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_41 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_41 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_41 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_41 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_41 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_41 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_41 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_41 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_41 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_41 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_41 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_41 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_41 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_41 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_41 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_41 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_41 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_41 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_41 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_41 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_41 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_41 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_41 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_41 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_41 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_41 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_41 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_41 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_41 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_41 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_41 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_41 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_41 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_41 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_41 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_41 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_41 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_41 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_41 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_41 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_41 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_41 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_41 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_41 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_41 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_41 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_41 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_41 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_41 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_41 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_41 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_41 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_41 = tailCount > 6'h29;
  wire          _GEN_1370 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h2A;
  wire          compressDataVec_hitReq_0_42;
  assign compressDataVec_hitReq_0_42 = _GEN_1370;
  wire          compressDataVec_hitReq_0_170;
  assign compressDataVec_hitReq_0_170 = _GEN_1370;
  wire          _GEN_1371 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h2A;
  wire          compressDataVec_hitReq_1_42;
  assign compressDataVec_hitReq_1_42 = _GEN_1371;
  wire          compressDataVec_hitReq_1_170;
  assign compressDataVec_hitReq_1_170 = _GEN_1371;
  wire          _GEN_1372 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h2A;
  wire          compressDataVec_hitReq_2_42;
  assign compressDataVec_hitReq_2_42 = _GEN_1372;
  wire          compressDataVec_hitReq_2_170;
  assign compressDataVec_hitReq_2_170 = _GEN_1372;
  wire          _GEN_1373 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h2A;
  wire          compressDataVec_hitReq_3_42;
  assign compressDataVec_hitReq_3_42 = _GEN_1373;
  wire          compressDataVec_hitReq_3_170;
  assign compressDataVec_hitReq_3_170 = _GEN_1373;
  wire          _GEN_1374 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h2A;
  wire          compressDataVec_hitReq_4_42;
  assign compressDataVec_hitReq_4_42 = _GEN_1374;
  wire          compressDataVec_hitReq_4_170;
  assign compressDataVec_hitReq_4_170 = _GEN_1374;
  wire          _GEN_1375 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h2A;
  wire          compressDataVec_hitReq_5_42;
  assign compressDataVec_hitReq_5_42 = _GEN_1375;
  wire          compressDataVec_hitReq_5_170;
  assign compressDataVec_hitReq_5_170 = _GEN_1375;
  wire          _GEN_1376 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h2A;
  wire          compressDataVec_hitReq_6_42;
  assign compressDataVec_hitReq_6_42 = _GEN_1376;
  wire          compressDataVec_hitReq_6_170;
  assign compressDataVec_hitReq_6_170 = _GEN_1376;
  wire          _GEN_1377 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h2A;
  wire          compressDataVec_hitReq_7_42;
  assign compressDataVec_hitReq_7_42 = _GEN_1377;
  wire          compressDataVec_hitReq_7_170;
  assign compressDataVec_hitReq_7_170 = _GEN_1377;
  wire          _GEN_1378 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h2A;
  wire          compressDataVec_hitReq_8_42;
  assign compressDataVec_hitReq_8_42 = _GEN_1378;
  wire          compressDataVec_hitReq_8_170;
  assign compressDataVec_hitReq_8_170 = _GEN_1378;
  wire          _GEN_1379 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h2A;
  wire          compressDataVec_hitReq_9_42;
  assign compressDataVec_hitReq_9_42 = _GEN_1379;
  wire          compressDataVec_hitReq_9_170;
  assign compressDataVec_hitReq_9_170 = _GEN_1379;
  wire          _GEN_1380 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h2A;
  wire          compressDataVec_hitReq_10_42;
  assign compressDataVec_hitReq_10_42 = _GEN_1380;
  wire          compressDataVec_hitReq_10_170;
  assign compressDataVec_hitReq_10_170 = _GEN_1380;
  wire          _GEN_1381 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h2A;
  wire          compressDataVec_hitReq_11_42;
  assign compressDataVec_hitReq_11_42 = _GEN_1381;
  wire          compressDataVec_hitReq_11_170;
  assign compressDataVec_hitReq_11_170 = _GEN_1381;
  wire          _GEN_1382 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h2A;
  wire          compressDataVec_hitReq_12_42;
  assign compressDataVec_hitReq_12_42 = _GEN_1382;
  wire          compressDataVec_hitReq_12_170;
  assign compressDataVec_hitReq_12_170 = _GEN_1382;
  wire          _GEN_1383 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h2A;
  wire          compressDataVec_hitReq_13_42;
  assign compressDataVec_hitReq_13_42 = _GEN_1383;
  wire          compressDataVec_hitReq_13_170;
  assign compressDataVec_hitReq_13_170 = _GEN_1383;
  wire          _GEN_1384 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h2A;
  wire          compressDataVec_hitReq_14_42;
  assign compressDataVec_hitReq_14_42 = _GEN_1384;
  wire          compressDataVec_hitReq_14_170;
  assign compressDataVec_hitReq_14_170 = _GEN_1384;
  wire          _GEN_1385 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h2A;
  wire          compressDataVec_hitReq_15_42;
  assign compressDataVec_hitReq_15_42 = _GEN_1385;
  wire          compressDataVec_hitReq_15_170;
  assign compressDataVec_hitReq_15_170 = _GEN_1385;
  wire          _GEN_1386 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h2A;
  wire          compressDataVec_hitReq_16_42;
  assign compressDataVec_hitReq_16_42 = _GEN_1386;
  wire          compressDataVec_hitReq_16_170;
  assign compressDataVec_hitReq_16_170 = _GEN_1386;
  wire          _GEN_1387 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h2A;
  wire          compressDataVec_hitReq_17_42;
  assign compressDataVec_hitReq_17_42 = _GEN_1387;
  wire          compressDataVec_hitReq_17_170;
  assign compressDataVec_hitReq_17_170 = _GEN_1387;
  wire          _GEN_1388 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h2A;
  wire          compressDataVec_hitReq_18_42;
  assign compressDataVec_hitReq_18_42 = _GEN_1388;
  wire          compressDataVec_hitReq_18_170;
  assign compressDataVec_hitReq_18_170 = _GEN_1388;
  wire          _GEN_1389 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h2A;
  wire          compressDataVec_hitReq_19_42;
  assign compressDataVec_hitReq_19_42 = _GEN_1389;
  wire          compressDataVec_hitReq_19_170;
  assign compressDataVec_hitReq_19_170 = _GEN_1389;
  wire          _GEN_1390 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h2A;
  wire          compressDataVec_hitReq_20_42;
  assign compressDataVec_hitReq_20_42 = _GEN_1390;
  wire          compressDataVec_hitReq_20_170;
  assign compressDataVec_hitReq_20_170 = _GEN_1390;
  wire          _GEN_1391 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h2A;
  wire          compressDataVec_hitReq_21_42;
  assign compressDataVec_hitReq_21_42 = _GEN_1391;
  wire          compressDataVec_hitReq_21_170;
  assign compressDataVec_hitReq_21_170 = _GEN_1391;
  wire          _GEN_1392 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h2A;
  wire          compressDataVec_hitReq_22_42;
  assign compressDataVec_hitReq_22_42 = _GEN_1392;
  wire          compressDataVec_hitReq_22_170;
  assign compressDataVec_hitReq_22_170 = _GEN_1392;
  wire          _GEN_1393 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h2A;
  wire          compressDataVec_hitReq_23_42;
  assign compressDataVec_hitReq_23_42 = _GEN_1393;
  wire          compressDataVec_hitReq_23_170;
  assign compressDataVec_hitReq_23_170 = _GEN_1393;
  wire          _GEN_1394 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h2A;
  wire          compressDataVec_hitReq_24_42;
  assign compressDataVec_hitReq_24_42 = _GEN_1394;
  wire          compressDataVec_hitReq_24_170;
  assign compressDataVec_hitReq_24_170 = _GEN_1394;
  wire          _GEN_1395 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h2A;
  wire          compressDataVec_hitReq_25_42;
  assign compressDataVec_hitReq_25_42 = _GEN_1395;
  wire          compressDataVec_hitReq_25_170;
  assign compressDataVec_hitReq_25_170 = _GEN_1395;
  wire          _GEN_1396 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h2A;
  wire          compressDataVec_hitReq_26_42;
  assign compressDataVec_hitReq_26_42 = _GEN_1396;
  wire          compressDataVec_hitReq_26_170;
  assign compressDataVec_hitReq_26_170 = _GEN_1396;
  wire          _GEN_1397 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h2A;
  wire          compressDataVec_hitReq_27_42;
  assign compressDataVec_hitReq_27_42 = _GEN_1397;
  wire          compressDataVec_hitReq_27_170;
  assign compressDataVec_hitReq_27_170 = _GEN_1397;
  wire          _GEN_1398 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h2A;
  wire          compressDataVec_hitReq_28_42;
  assign compressDataVec_hitReq_28_42 = _GEN_1398;
  wire          compressDataVec_hitReq_28_170;
  assign compressDataVec_hitReq_28_170 = _GEN_1398;
  wire          _GEN_1399 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h2A;
  wire          compressDataVec_hitReq_29_42;
  assign compressDataVec_hitReq_29_42 = _GEN_1399;
  wire          compressDataVec_hitReq_29_170;
  assign compressDataVec_hitReq_29_170 = _GEN_1399;
  wire          _GEN_1400 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h2A;
  wire          compressDataVec_hitReq_30_42;
  assign compressDataVec_hitReq_30_42 = _GEN_1400;
  wire          compressDataVec_hitReq_30_170;
  assign compressDataVec_hitReq_30_170 = _GEN_1400;
  wire          _GEN_1401 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h2A;
  wire          compressDataVec_hitReq_31_42;
  assign compressDataVec_hitReq_31_42 = _GEN_1401;
  wire          compressDataVec_hitReq_31_170;
  assign compressDataVec_hitReq_31_170 = _GEN_1401;
  wire          compressDataVec_hitReq_32_42 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h2A;
  wire          compressDataVec_hitReq_33_42 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h2A;
  wire          compressDataVec_hitReq_34_42 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h2A;
  wire          compressDataVec_hitReq_35_42 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h2A;
  wire          compressDataVec_hitReq_36_42 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h2A;
  wire          compressDataVec_hitReq_37_42 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h2A;
  wire          compressDataVec_hitReq_38_42 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h2A;
  wire          compressDataVec_hitReq_39_42 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h2A;
  wire          compressDataVec_hitReq_40_42 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h2A;
  wire          compressDataVec_hitReq_41_42 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h2A;
  wire          compressDataVec_hitReq_42_42 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h2A;
  wire          compressDataVec_hitReq_43_42 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h2A;
  wire          compressDataVec_hitReq_44_42 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h2A;
  wire          compressDataVec_hitReq_45_42 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h2A;
  wire          compressDataVec_hitReq_46_42 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h2A;
  wire          compressDataVec_hitReq_47_42 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h2A;
  wire          compressDataVec_hitReq_48_42 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h2A;
  wire          compressDataVec_hitReq_49_42 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h2A;
  wire          compressDataVec_hitReq_50_42 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h2A;
  wire          compressDataVec_hitReq_51_42 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h2A;
  wire          compressDataVec_hitReq_52_42 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h2A;
  wire          compressDataVec_hitReq_53_42 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h2A;
  wire          compressDataVec_hitReq_54_42 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h2A;
  wire          compressDataVec_hitReq_55_42 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h2A;
  wire          compressDataVec_hitReq_56_42 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h2A;
  wire          compressDataVec_hitReq_57_42 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h2A;
  wire          compressDataVec_hitReq_58_42 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h2A;
  wire          compressDataVec_hitReq_59_42 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h2A;
  wire          compressDataVec_hitReq_60_42 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h2A;
  wire          compressDataVec_hitReq_61_42 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h2A;
  wire          compressDataVec_hitReq_62_42 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h2A;
  wire          compressDataVec_hitReq_63_42 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h2A;
  wire [7:0]    compressDataVec_selectReqData_42 =
    (compressDataVec_hitReq_0_42 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_42 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_42 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_42 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_42 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_42 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_42 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_42 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_42 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_42 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_42 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_42 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_42 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_42 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_42 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_42 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_42 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_42 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_42 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_42 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_42 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_42 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_42 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_42 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_42 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_42 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_42 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_42 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_42 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_42 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_42 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_42 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_42 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_42 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_42 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_42 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_42 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_42 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_42 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_42 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_42 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_42 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_42 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_42 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_42 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_42 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_42 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_42 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_42 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_42 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_42 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_42 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_42 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_42 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_42 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_42 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_42 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_42 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_42 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_42 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_42 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_42 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_42 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_42 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_42 = tailCount > 6'h2A;
  wire          _GEN_1402 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h2B;
  wire          compressDataVec_hitReq_0_43;
  assign compressDataVec_hitReq_0_43 = _GEN_1402;
  wire          compressDataVec_hitReq_0_171;
  assign compressDataVec_hitReq_0_171 = _GEN_1402;
  wire          _GEN_1403 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h2B;
  wire          compressDataVec_hitReq_1_43;
  assign compressDataVec_hitReq_1_43 = _GEN_1403;
  wire          compressDataVec_hitReq_1_171;
  assign compressDataVec_hitReq_1_171 = _GEN_1403;
  wire          _GEN_1404 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h2B;
  wire          compressDataVec_hitReq_2_43;
  assign compressDataVec_hitReq_2_43 = _GEN_1404;
  wire          compressDataVec_hitReq_2_171;
  assign compressDataVec_hitReq_2_171 = _GEN_1404;
  wire          _GEN_1405 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h2B;
  wire          compressDataVec_hitReq_3_43;
  assign compressDataVec_hitReq_3_43 = _GEN_1405;
  wire          compressDataVec_hitReq_3_171;
  assign compressDataVec_hitReq_3_171 = _GEN_1405;
  wire          _GEN_1406 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h2B;
  wire          compressDataVec_hitReq_4_43;
  assign compressDataVec_hitReq_4_43 = _GEN_1406;
  wire          compressDataVec_hitReq_4_171;
  assign compressDataVec_hitReq_4_171 = _GEN_1406;
  wire          _GEN_1407 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h2B;
  wire          compressDataVec_hitReq_5_43;
  assign compressDataVec_hitReq_5_43 = _GEN_1407;
  wire          compressDataVec_hitReq_5_171;
  assign compressDataVec_hitReq_5_171 = _GEN_1407;
  wire          _GEN_1408 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h2B;
  wire          compressDataVec_hitReq_6_43;
  assign compressDataVec_hitReq_6_43 = _GEN_1408;
  wire          compressDataVec_hitReq_6_171;
  assign compressDataVec_hitReq_6_171 = _GEN_1408;
  wire          _GEN_1409 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h2B;
  wire          compressDataVec_hitReq_7_43;
  assign compressDataVec_hitReq_7_43 = _GEN_1409;
  wire          compressDataVec_hitReq_7_171;
  assign compressDataVec_hitReq_7_171 = _GEN_1409;
  wire          _GEN_1410 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h2B;
  wire          compressDataVec_hitReq_8_43;
  assign compressDataVec_hitReq_8_43 = _GEN_1410;
  wire          compressDataVec_hitReq_8_171;
  assign compressDataVec_hitReq_8_171 = _GEN_1410;
  wire          _GEN_1411 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h2B;
  wire          compressDataVec_hitReq_9_43;
  assign compressDataVec_hitReq_9_43 = _GEN_1411;
  wire          compressDataVec_hitReq_9_171;
  assign compressDataVec_hitReq_9_171 = _GEN_1411;
  wire          _GEN_1412 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h2B;
  wire          compressDataVec_hitReq_10_43;
  assign compressDataVec_hitReq_10_43 = _GEN_1412;
  wire          compressDataVec_hitReq_10_171;
  assign compressDataVec_hitReq_10_171 = _GEN_1412;
  wire          _GEN_1413 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h2B;
  wire          compressDataVec_hitReq_11_43;
  assign compressDataVec_hitReq_11_43 = _GEN_1413;
  wire          compressDataVec_hitReq_11_171;
  assign compressDataVec_hitReq_11_171 = _GEN_1413;
  wire          _GEN_1414 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h2B;
  wire          compressDataVec_hitReq_12_43;
  assign compressDataVec_hitReq_12_43 = _GEN_1414;
  wire          compressDataVec_hitReq_12_171;
  assign compressDataVec_hitReq_12_171 = _GEN_1414;
  wire          _GEN_1415 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h2B;
  wire          compressDataVec_hitReq_13_43;
  assign compressDataVec_hitReq_13_43 = _GEN_1415;
  wire          compressDataVec_hitReq_13_171;
  assign compressDataVec_hitReq_13_171 = _GEN_1415;
  wire          _GEN_1416 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h2B;
  wire          compressDataVec_hitReq_14_43;
  assign compressDataVec_hitReq_14_43 = _GEN_1416;
  wire          compressDataVec_hitReq_14_171;
  assign compressDataVec_hitReq_14_171 = _GEN_1416;
  wire          _GEN_1417 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h2B;
  wire          compressDataVec_hitReq_15_43;
  assign compressDataVec_hitReq_15_43 = _GEN_1417;
  wire          compressDataVec_hitReq_15_171;
  assign compressDataVec_hitReq_15_171 = _GEN_1417;
  wire          _GEN_1418 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h2B;
  wire          compressDataVec_hitReq_16_43;
  assign compressDataVec_hitReq_16_43 = _GEN_1418;
  wire          compressDataVec_hitReq_16_171;
  assign compressDataVec_hitReq_16_171 = _GEN_1418;
  wire          _GEN_1419 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h2B;
  wire          compressDataVec_hitReq_17_43;
  assign compressDataVec_hitReq_17_43 = _GEN_1419;
  wire          compressDataVec_hitReq_17_171;
  assign compressDataVec_hitReq_17_171 = _GEN_1419;
  wire          _GEN_1420 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h2B;
  wire          compressDataVec_hitReq_18_43;
  assign compressDataVec_hitReq_18_43 = _GEN_1420;
  wire          compressDataVec_hitReq_18_171;
  assign compressDataVec_hitReq_18_171 = _GEN_1420;
  wire          _GEN_1421 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h2B;
  wire          compressDataVec_hitReq_19_43;
  assign compressDataVec_hitReq_19_43 = _GEN_1421;
  wire          compressDataVec_hitReq_19_171;
  assign compressDataVec_hitReq_19_171 = _GEN_1421;
  wire          _GEN_1422 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h2B;
  wire          compressDataVec_hitReq_20_43;
  assign compressDataVec_hitReq_20_43 = _GEN_1422;
  wire          compressDataVec_hitReq_20_171;
  assign compressDataVec_hitReq_20_171 = _GEN_1422;
  wire          _GEN_1423 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h2B;
  wire          compressDataVec_hitReq_21_43;
  assign compressDataVec_hitReq_21_43 = _GEN_1423;
  wire          compressDataVec_hitReq_21_171;
  assign compressDataVec_hitReq_21_171 = _GEN_1423;
  wire          _GEN_1424 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h2B;
  wire          compressDataVec_hitReq_22_43;
  assign compressDataVec_hitReq_22_43 = _GEN_1424;
  wire          compressDataVec_hitReq_22_171;
  assign compressDataVec_hitReq_22_171 = _GEN_1424;
  wire          _GEN_1425 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h2B;
  wire          compressDataVec_hitReq_23_43;
  assign compressDataVec_hitReq_23_43 = _GEN_1425;
  wire          compressDataVec_hitReq_23_171;
  assign compressDataVec_hitReq_23_171 = _GEN_1425;
  wire          _GEN_1426 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h2B;
  wire          compressDataVec_hitReq_24_43;
  assign compressDataVec_hitReq_24_43 = _GEN_1426;
  wire          compressDataVec_hitReq_24_171;
  assign compressDataVec_hitReq_24_171 = _GEN_1426;
  wire          _GEN_1427 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h2B;
  wire          compressDataVec_hitReq_25_43;
  assign compressDataVec_hitReq_25_43 = _GEN_1427;
  wire          compressDataVec_hitReq_25_171;
  assign compressDataVec_hitReq_25_171 = _GEN_1427;
  wire          _GEN_1428 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h2B;
  wire          compressDataVec_hitReq_26_43;
  assign compressDataVec_hitReq_26_43 = _GEN_1428;
  wire          compressDataVec_hitReq_26_171;
  assign compressDataVec_hitReq_26_171 = _GEN_1428;
  wire          _GEN_1429 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h2B;
  wire          compressDataVec_hitReq_27_43;
  assign compressDataVec_hitReq_27_43 = _GEN_1429;
  wire          compressDataVec_hitReq_27_171;
  assign compressDataVec_hitReq_27_171 = _GEN_1429;
  wire          _GEN_1430 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h2B;
  wire          compressDataVec_hitReq_28_43;
  assign compressDataVec_hitReq_28_43 = _GEN_1430;
  wire          compressDataVec_hitReq_28_171;
  assign compressDataVec_hitReq_28_171 = _GEN_1430;
  wire          _GEN_1431 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h2B;
  wire          compressDataVec_hitReq_29_43;
  assign compressDataVec_hitReq_29_43 = _GEN_1431;
  wire          compressDataVec_hitReq_29_171;
  assign compressDataVec_hitReq_29_171 = _GEN_1431;
  wire          _GEN_1432 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h2B;
  wire          compressDataVec_hitReq_30_43;
  assign compressDataVec_hitReq_30_43 = _GEN_1432;
  wire          compressDataVec_hitReq_30_171;
  assign compressDataVec_hitReq_30_171 = _GEN_1432;
  wire          _GEN_1433 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h2B;
  wire          compressDataVec_hitReq_31_43;
  assign compressDataVec_hitReq_31_43 = _GEN_1433;
  wire          compressDataVec_hitReq_31_171;
  assign compressDataVec_hitReq_31_171 = _GEN_1433;
  wire          compressDataVec_hitReq_32_43 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h2B;
  wire          compressDataVec_hitReq_33_43 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h2B;
  wire          compressDataVec_hitReq_34_43 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h2B;
  wire          compressDataVec_hitReq_35_43 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h2B;
  wire          compressDataVec_hitReq_36_43 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h2B;
  wire          compressDataVec_hitReq_37_43 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h2B;
  wire          compressDataVec_hitReq_38_43 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h2B;
  wire          compressDataVec_hitReq_39_43 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h2B;
  wire          compressDataVec_hitReq_40_43 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h2B;
  wire          compressDataVec_hitReq_41_43 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h2B;
  wire          compressDataVec_hitReq_42_43 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h2B;
  wire          compressDataVec_hitReq_43_43 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h2B;
  wire          compressDataVec_hitReq_44_43 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h2B;
  wire          compressDataVec_hitReq_45_43 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h2B;
  wire          compressDataVec_hitReq_46_43 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h2B;
  wire          compressDataVec_hitReq_47_43 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h2B;
  wire          compressDataVec_hitReq_48_43 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h2B;
  wire          compressDataVec_hitReq_49_43 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h2B;
  wire          compressDataVec_hitReq_50_43 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h2B;
  wire          compressDataVec_hitReq_51_43 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h2B;
  wire          compressDataVec_hitReq_52_43 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h2B;
  wire          compressDataVec_hitReq_53_43 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h2B;
  wire          compressDataVec_hitReq_54_43 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h2B;
  wire          compressDataVec_hitReq_55_43 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h2B;
  wire          compressDataVec_hitReq_56_43 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h2B;
  wire          compressDataVec_hitReq_57_43 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h2B;
  wire          compressDataVec_hitReq_58_43 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h2B;
  wire          compressDataVec_hitReq_59_43 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h2B;
  wire          compressDataVec_hitReq_60_43 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h2B;
  wire          compressDataVec_hitReq_61_43 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h2B;
  wire          compressDataVec_hitReq_62_43 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h2B;
  wire          compressDataVec_hitReq_63_43 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h2B;
  wire [7:0]    compressDataVec_selectReqData_43 =
    (compressDataVec_hitReq_0_43 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_43 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_43 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_43 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_43 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_43 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_43 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_43 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_43 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_43 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_43 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_43 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_43 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_43 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_43 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_43 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_43 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_43 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_43 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_43 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_43 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_43 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_43 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_43 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_43 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_43 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_43 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_43 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_43 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_43 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_43 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_43 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_43 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_43 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_43 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_43 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_43 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_43 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_43 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_43 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_43 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_43 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_43 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_43 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_43 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_43 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_43 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_43 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_43 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_43 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_43 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_43 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_43 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_43 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_43 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_43 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_43 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_43 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_43 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_43 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_43 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_43 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_43 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_43 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_43 = tailCount > 6'h2B;
  wire          _GEN_1434 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h2C;
  wire          compressDataVec_hitReq_0_44;
  assign compressDataVec_hitReq_0_44 = _GEN_1434;
  wire          compressDataVec_hitReq_0_172;
  assign compressDataVec_hitReq_0_172 = _GEN_1434;
  wire          _GEN_1435 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h2C;
  wire          compressDataVec_hitReq_1_44;
  assign compressDataVec_hitReq_1_44 = _GEN_1435;
  wire          compressDataVec_hitReq_1_172;
  assign compressDataVec_hitReq_1_172 = _GEN_1435;
  wire          _GEN_1436 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h2C;
  wire          compressDataVec_hitReq_2_44;
  assign compressDataVec_hitReq_2_44 = _GEN_1436;
  wire          compressDataVec_hitReq_2_172;
  assign compressDataVec_hitReq_2_172 = _GEN_1436;
  wire          _GEN_1437 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h2C;
  wire          compressDataVec_hitReq_3_44;
  assign compressDataVec_hitReq_3_44 = _GEN_1437;
  wire          compressDataVec_hitReq_3_172;
  assign compressDataVec_hitReq_3_172 = _GEN_1437;
  wire          _GEN_1438 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h2C;
  wire          compressDataVec_hitReq_4_44;
  assign compressDataVec_hitReq_4_44 = _GEN_1438;
  wire          compressDataVec_hitReq_4_172;
  assign compressDataVec_hitReq_4_172 = _GEN_1438;
  wire          _GEN_1439 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h2C;
  wire          compressDataVec_hitReq_5_44;
  assign compressDataVec_hitReq_5_44 = _GEN_1439;
  wire          compressDataVec_hitReq_5_172;
  assign compressDataVec_hitReq_5_172 = _GEN_1439;
  wire          _GEN_1440 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h2C;
  wire          compressDataVec_hitReq_6_44;
  assign compressDataVec_hitReq_6_44 = _GEN_1440;
  wire          compressDataVec_hitReq_6_172;
  assign compressDataVec_hitReq_6_172 = _GEN_1440;
  wire          _GEN_1441 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h2C;
  wire          compressDataVec_hitReq_7_44;
  assign compressDataVec_hitReq_7_44 = _GEN_1441;
  wire          compressDataVec_hitReq_7_172;
  assign compressDataVec_hitReq_7_172 = _GEN_1441;
  wire          _GEN_1442 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h2C;
  wire          compressDataVec_hitReq_8_44;
  assign compressDataVec_hitReq_8_44 = _GEN_1442;
  wire          compressDataVec_hitReq_8_172;
  assign compressDataVec_hitReq_8_172 = _GEN_1442;
  wire          _GEN_1443 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h2C;
  wire          compressDataVec_hitReq_9_44;
  assign compressDataVec_hitReq_9_44 = _GEN_1443;
  wire          compressDataVec_hitReq_9_172;
  assign compressDataVec_hitReq_9_172 = _GEN_1443;
  wire          _GEN_1444 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h2C;
  wire          compressDataVec_hitReq_10_44;
  assign compressDataVec_hitReq_10_44 = _GEN_1444;
  wire          compressDataVec_hitReq_10_172;
  assign compressDataVec_hitReq_10_172 = _GEN_1444;
  wire          _GEN_1445 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h2C;
  wire          compressDataVec_hitReq_11_44;
  assign compressDataVec_hitReq_11_44 = _GEN_1445;
  wire          compressDataVec_hitReq_11_172;
  assign compressDataVec_hitReq_11_172 = _GEN_1445;
  wire          _GEN_1446 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h2C;
  wire          compressDataVec_hitReq_12_44;
  assign compressDataVec_hitReq_12_44 = _GEN_1446;
  wire          compressDataVec_hitReq_12_172;
  assign compressDataVec_hitReq_12_172 = _GEN_1446;
  wire          _GEN_1447 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h2C;
  wire          compressDataVec_hitReq_13_44;
  assign compressDataVec_hitReq_13_44 = _GEN_1447;
  wire          compressDataVec_hitReq_13_172;
  assign compressDataVec_hitReq_13_172 = _GEN_1447;
  wire          _GEN_1448 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h2C;
  wire          compressDataVec_hitReq_14_44;
  assign compressDataVec_hitReq_14_44 = _GEN_1448;
  wire          compressDataVec_hitReq_14_172;
  assign compressDataVec_hitReq_14_172 = _GEN_1448;
  wire          _GEN_1449 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h2C;
  wire          compressDataVec_hitReq_15_44;
  assign compressDataVec_hitReq_15_44 = _GEN_1449;
  wire          compressDataVec_hitReq_15_172;
  assign compressDataVec_hitReq_15_172 = _GEN_1449;
  wire          _GEN_1450 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h2C;
  wire          compressDataVec_hitReq_16_44;
  assign compressDataVec_hitReq_16_44 = _GEN_1450;
  wire          compressDataVec_hitReq_16_172;
  assign compressDataVec_hitReq_16_172 = _GEN_1450;
  wire          _GEN_1451 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h2C;
  wire          compressDataVec_hitReq_17_44;
  assign compressDataVec_hitReq_17_44 = _GEN_1451;
  wire          compressDataVec_hitReq_17_172;
  assign compressDataVec_hitReq_17_172 = _GEN_1451;
  wire          _GEN_1452 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h2C;
  wire          compressDataVec_hitReq_18_44;
  assign compressDataVec_hitReq_18_44 = _GEN_1452;
  wire          compressDataVec_hitReq_18_172;
  assign compressDataVec_hitReq_18_172 = _GEN_1452;
  wire          _GEN_1453 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h2C;
  wire          compressDataVec_hitReq_19_44;
  assign compressDataVec_hitReq_19_44 = _GEN_1453;
  wire          compressDataVec_hitReq_19_172;
  assign compressDataVec_hitReq_19_172 = _GEN_1453;
  wire          _GEN_1454 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h2C;
  wire          compressDataVec_hitReq_20_44;
  assign compressDataVec_hitReq_20_44 = _GEN_1454;
  wire          compressDataVec_hitReq_20_172;
  assign compressDataVec_hitReq_20_172 = _GEN_1454;
  wire          _GEN_1455 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h2C;
  wire          compressDataVec_hitReq_21_44;
  assign compressDataVec_hitReq_21_44 = _GEN_1455;
  wire          compressDataVec_hitReq_21_172;
  assign compressDataVec_hitReq_21_172 = _GEN_1455;
  wire          _GEN_1456 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h2C;
  wire          compressDataVec_hitReq_22_44;
  assign compressDataVec_hitReq_22_44 = _GEN_1456;
  wire          compressDataVec_hitReq_22_172;
  assign compressDataVec_hitReq_22_172 = _GEN_1456;
  wire          _GEN_1457 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h2C;
  wire          compressDataVec_hitReq_23_44;
  assign compressDataVec_hitReq_23_44 = _GEN_1457;
  wire          compressDataVec_hitReq_23_172;
  assign compressDataVec_hitReq_23_172 = _GEN_1457;
  wire          _GEN_1458 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h2C;
  wire          compressDataVec_hitReq_24_44;
  assign compressDataVec_hitReq_24_44 = _GEN_1458;
  wire          compressDataVec_hitReq_24_172;
  assign compressDataVec_hitReq_24_172 = _GEN_1458;
  wire          _GEN_1459 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h2C;
  wire          compressDataVec_hitReq_25_44;
  assign compressDataVec_hitReq_25_44 = _GEN_1459;
  wire          compressDataVec_hitReq_25_172;
  assign compressDataVec_hitReq_25_172 = _GEN_1459;
  wire          _GEN_1460 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h2C;
  wire          compressDataVec_hitReq_26_44;
  assign compressDataVec_hitReq_26_44 = _GEN_1460;
  wire          compressDataVec_hitReq_26_172;
  assign compressDataVec_hitReq_26_172 = _GEN_1460;
  wire          _GEN_1461 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h2C;
  wire          compressDataVec_hitReq_27_44;
  assign compressDataVec_hitReq_27_44 = _GEN_1461;
  wire          compressDataVec_hitReq_27_172;
  assign compressDataVec_hitReq_27_172 = _GEN_1461;
  wire          _GEN_1462 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h2C;
  wire          compressDataVec_hitReq_28_44;
  assign compressDataVec_hitReq_28_44 = _GEN_1462;
  wire          compressDataVec_hitReq_28_172;
  assign compressDataVec_hitReq_28_172 = _GEN_1462;
  wire          _GEN_1463 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h2C;
  wire          compressDataVec_hitReq_29_44;
  assign compressDataVec_hitReq_29_44 = _GEN_1463;
  wire          compressDataVec_hitReq_29_172;
  assign compressDataVec_hitReq_29_172 = _GEN_1463;
  wire          _GEN_1464 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h2C;
  wire          compressDataVec_hitReq_30_44;
  assign compressDataVec_hitReq_30_44 = _GEN_1464;
  wire          compressDataVec_hitReq_30_172;
  assign compressDataVec_hitReq_30_172 = _GEN_1464;
  wire          _GEN_1465 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h2C;
  wire          compressDataVec_hitReq_31_44;
  assign compressDataVec_hitReq_31_44 = _GEN_1465;
  wire          compressDataVec_hitReq_31_172;
  assign compressDataVec_hitReq_31_172 = _GEN_1465;
  wire          compressDataVec_hitReq_32_44 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h2C;
  wire          compressDataVec_hitReq_33_44 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h2C;
  wire          compressDataVec_hitReq_34_44 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h2C;
  wire          compressDataVec_hitReq_35_44 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h2C;
  wire          compressDataVec_hitReq_36_44 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h2C;
  wire          compressDataVec_hitReq_37_44 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h2C;
  wire          compressDataVec_hitReq_38_44 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h2C;
  wire          compressDataVec_hitReq_39_44 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h2C;
  wire          compressDataVec_hitReq_40_44 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h2C;
  wire          compressDataVec_hitReq_41_44 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h2C;
  wire          compressDataVec_hitReq_42_44 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h2C;
  wire          compressDataVec_hitReq_43_44 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h2C;
  wire          compressDataVec_hitReq_44_44 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h2C;
  wire          compressDataVec_hitReq_45_44 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h2C;
  wire          compressDataVec_hitReq_46_44 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h2C;
  wire          compressDataVec_hitReq_47_44 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h2C;
  wire          compressDataVec_hitReq_48_44 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h2C;
  wire          compressDataVec_hitReq_49_44 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h2C;
  wire          compressDataVec_hitReq_50_44 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h2C;
  wire          compressDataVec_hitReq_51_44 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h2C;
  wire          compressDataVec_hitReq_52_44 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h2C;
  wire          compressDataVec_hitReq_53_44 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h2C;
  wire          compressDataVec_hitReq_54_44 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h2C;
  wire          compressDataVec_hitReq_55_44 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h2C;
  wire          compressDataVec_hitReq_56_44 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h2C;
  wire          compressDataVec_hitReq_57_44 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h2C;
  wire          compressDataVec_hitReq_58_44 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h2C;
  wire          compressDataVec_hitReq_59_44 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h2C;
  wire          compressDataVec_hitReq_60_44 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h2C;
  wire          compressDataVec_hitReq_61_44 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h2C;
  wire          compressDataVec_hitReq_62_44 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h2C;
  wire          compressDataVec_hitReq_63_44 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h2C;
  wire [7:0]    compressDataVec_selectReqData_44 =
    (compressDataVec_hitReq_0_44 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_44 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_44 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_44 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_44 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_44 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_44 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_44 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_44 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_44 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_44 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_44 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_44 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_44 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_44 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_44 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_44 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_44 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_44 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_44 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_44 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_44 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_44 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_44 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_44 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_44 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_44 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_44 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_44 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_44 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_44 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_44 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_44 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_44 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_44 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_44 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_44 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_44 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_44 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_44 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_44 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_44 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_44 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_44 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_44 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_44 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_44 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_44 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_44 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_44 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_44 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_44 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_44 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_44 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_44 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_44 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_44 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_44 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_44 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_44 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_44 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_44 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_44 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_44 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_44 = tailCount > 6'h2C;
  wire          _GEN_1466 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h2D;
  wire          compressDataVec_hitReq_0_45;
  assign compressDataVec_hitReq_0_45 = _GEN_1466;
  wire          compressDataVec_hitReq_0_173;
  assign compressDataVec_hitReq_0_173 = _GEN_1466;
  wire          _GEN_1467 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h2D;
  wire          compressDataVec_hitReq_1_45;
  assign compressDataVec_hitReq_1_45 = _GEN_1467;
  wire          compressDataVec_hitReq_1_173;
  assign compressDataVec_hitReq_1_173 = _GEN_1467;
  wire          _GEN_1468 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h2D;
  wire          compressDataVec_hitReq_2_45;
  assign compressDataVec_hitReq_2_45 = _GEN_1468;
  wire          compressDataVec_hitReq_2_173;
  assign compressDataVec_hitReq_2_173 = _GEN_1468;
  wire          _GEN_1469 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h2D;
  wire          compressDataVec_hitReq_3_45;
  assign compressDataVec_hitReq_3_45 = _GEN_1469;
  wire          compressDataVec_hitReq_3_173;
  assign compressDataVec_hitReq_3_173 = _GEN_1469;
  wire          _GEN_1470 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h2D;
  wire          compressDataVec_hitReq_4_45;
  assign compressDataVec_hitReq_4_45 = _GEN_1470;
  wire          compressDataVec_hitReq_4_173;
  assign compressDataVec_hitReq_4_173 = _GEN_1470;
  wire          _GEN_1471 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h2D;
  wire          compressDataVec_hitReq_5_45;
  assign compressDataVec_hitReq_5_45 = _GEN_1471;
  wire          compressDataVec_hitReq_5_173;
  assign compressDataVec_hitReq_5_173 = _GEN_1471;
  wire          _GEN_1472 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h2D;
  wire          compressDataVec_hitReq_6_45;
  assign compressDataVec_hitReq_6_45 = _GEN_1472;
  wire          compressDataVec_hitReq_6_173;
  assign compressDataVec_hitReq_6_173 = _GEN_1472;
  wire          _GEN_1473 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h2D;
  wire          compressDataVec_hitReq_7_45;
  assign compressDataVec_hitReq_7_45 = _GEN_1473;
  wire          compressDataVec_hitReq_7_173;
  assign compressDataVec_hitReq_7_173 = _GEN_1473;
  wire          _GEN_1474 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h2D;
  wire          compressDataVec_hitReq_8_45;
  assign compressDataVec_hitReq_8_45 = _GEN_1474;
  wire          compressDataVec_hitReq_8_173;
  assign compressDataVec_hitReq_8_173 = _GEN_1474;
  wire          _GEN_1475 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h2D;
  wire          compressDataVec_hitReq_9_45;
  assign compressDataVec_hitReq_9_45 = _GEN_1475;
  wire          compressDataVec_hitReq_9_173;
  assign compressDataVec_hitReq_9_173 = _GEN_1475;
  wire          _GEN_1476 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h2D;
  wire          compressDataVec_hitReq_10_45;
  assign compressDataVec_hitReq_10_45 = _GEN_1476;
  wire          compressDataVec_hitReq_10_173;
  assign compressDataVec_hitReq_10_173 = _GEN_1476;
  wire          _GEN_1477 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h2D;
  wire          compressDataVec_hitReq_11_45;
  assign compressDataVec_hitReq_11_45 = _GEN_1477;
  wire          compressDataVec_hitReq_11_173;
  assign compressDataVec_hitReq_11_173 = _GEN_1477;
  wire          _GEN_1478 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h2D;
  wire          compressDataVec_hitReq_12_45;
  assign compressDataVec_hitReq_12_45 = _GEN_1478;
  wire          compressDataVec_hitReq_12_173;
  assign compressDataVec_hitReq_12_173 = _GEN_1478;
  wire          _GEN_1479 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h2D;
  wire          compressDataVec_hitReq_13_45;
  assign compressDataVec_hitReq_13_45 = _GEN_1479;
  wire          compressDataVec_hitReq_13_173;
  assign compressDataVec_hitReq_13_173 = _GEN_1479;
  wire          _GEN_1480 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h2D;
  wire          compressDataVec_hitReq_14_45;
  assign compressDataVec_hitReq_14_45 = _GEN_1480;
  wire          compressDataVec_hitReq_14_173;
  assign compressDataVec_hitReq_14_173 = _GEN_1480;
  wire          _GEN_1481 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h2D;
  wire          compressDataVec_hitReq_15_45;
  assign compressDataVec_hitReq_15_45 = _GEN_1481;
  wire          compressDataVec_hitReq_15_173;
  assign compressDataVec_hitReq_15_173 = _GEN_1481;
  wire          _GEN_1482 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h2D;
  wire          compressDataVec_hitReq_16_45;
  assign compressDataVec_hitReq_16_45 = _GEN_1482;
  wire          compressDataVec_hitReq_16_173;
  assign compressDataVec_hitReq_16_173 = _GEN_1482;
  wire          _GEN_1483 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h2D;
  wire          compressDataVec_hitReq_17_45;
  assign compressDataVec_hitReq_17_45 = _GEN_1483;
  wire          compressDataVec_hitReq_17_173;
  assign compressDataVec_hitReq_17_173 = _GEN_1483;
  wire          _GEN_1484 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h2D;
  wire          compressDataVec_hitReq_18_45;
  assign compressDataVec_hitReq_18_45 = _GEN_1484;
  wire          compressDataVec_hitReq_18_173;
  assign compressDataVec_hitReq_18_173 = _GEN_1484;
  wire          _GEN_1485 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h2D;
  wire          compressDataVec_hitReq_19_45;
  assign compressDataVec_hitReq_19_45 = _GEN_1485;
  wire          compressDataVec_hitReq_19_173;
  assign compressDataVec_hitReq_19_173 = _GEN_1485;
  wire          _GEN_1486 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h2D;
  wire          compressDataVec_hitReq_20_45;
  assign compressDataVec_hitReq_20_45 = _GEN_1486;
  wire          compressDataVec_hitReq_20_173;
  assign compressDataVec_hitReq_20_173 = _GEN_1486;
  wire          _GEN_1487 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h2D;
  wire          compressDataVec_hitReq_21_45;
  assign compressDataVec_hitReq_21_45 = _GEN_1487;
  wire          compressDataVec_hitReq_21_173;
  assign compressDataVec_hitReq_21_173 = _GEN_1487;
  wire          _GEN_1488 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h2D;
  wire          compressDataVec_hitReq_22_45;
  assign compressDataVec_hitReq_22_45 = _GEN_1488;
  wire          compressDataVec_hitReq_22_173;
  assign compressDataVec_hitReq_22_173 = _GEN_1488;
  wire          _GEN_1489 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h2D;
  wire          compressDataVec_hitReq_23_45;
  assign compressDataVec_hitReq_23_45 = _GEN_1489;
  wire          compressDataVec_hitReq_23_173;
  assign compressDataVec_hitReq_23_173 = _GEN_1489;
  wire          _GEN_1490 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h2D;
  wire          compressDataVec_hitReq_24_45;
  assign compressDataVec_hitReq_24_45 = _GEN_1490;
  wire          compressDataVec_hitReq_24_173;
  assign compressDataVec_hitReq_24_173 = _GEN_1490;
  wire          _GEN_1491 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h2D;
  wire          compressDataVec_hitReq_25_45;
  assign compressDataVec_hitReq_25_45 = _GEN_1491;
  wire          compressDataVec_hitReq_25_173;
  assign compressDataVec_hitReq_25_173 = _GEN_1491;
  wire          _GEN_1492 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h2D;
  wire          compressDataVec_hitReq_26_45;
  assign compressDataVec_hitReq_26_45 = _GEN_1492;
  wire          compressDataVec_hitReq_26_173;
  assign compressDataVec_hitReq_26_173 = _GEN_1492;
  wire          _GEN_1493 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h2D;
  wire          compressDataVec_hitReq_27_45;
  assign compressDataVec_hitReq_27_45 = _GEN_1493;
  wire          compressDataVec_hitReq_27_173;
  assign compressDataVec_hitReq_27_173 = _GEN_1493;
  wire          _GEN_1494 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h2D;
  wire          compressDataVec_hitReq_28_45;
  assign compressDataVec_hitReq_28_45 = _GEN_1494;
  wire          compressDataVec_hitReq_28_173;
  assign compressDataVec_hitReq_28_173 = _GEN_1494;
  wire          _GEN_1495 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h2D;
  wire          compressDataVec_hitReq_29_45;
  assign compressDataVec_hitReq_29_45 = _GEN_1495;
  wire          compressDataVec_hitReq_29_173;
  assign compressDataVec_hitReq_29_173 = _GEN_1495;
  wire          _GEN_1496 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h2D;
  wire          compressDataVec_hitReq_30_45;
  assign compressDataVec_hitReq_30_45 = _GEN_1496;
  wire          compressDataVec_hitReq_30_173;
  assign compressDataVec_hitReq_30_173 = _GEN_1496;
  wire          _GEN_1497 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h2D;
  wire          compressDataVec_hitReq_31_45;
  assign compressDataVec_hitReq_31_45 = _GEN_1497;
  wire          compressDataVec_hitReq_31_173;
  assign compressDataVec_hitReq_31_173 = _GEN_1497;
  wire          compressDataVec_hitReq_32_45 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h2D;
  wire          compressDataVec_hitReq_33_45 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h2D;
  wire          compressDataVec_hitReq_34_45 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h2D;
  wire          compressDataVec_hitReq_35_45 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h2D;
  wire          compressDataVec_hitReq_36_45 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h2D;
  wire          compressDataVec_hitReq_37_45 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h2D;
  wire          compressDataVec_hitReq_38_45 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h2D;
  wire          compressDataVec_hitReq_39_45 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h2D;
  wire          compressDataVec_hitReq_40_45 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h2D;
  wire          compressDataVec_hitReq_41_45 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h2D;
  wire          compressDataVec_hitReq_42_45 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h2D;
  wire          compressDataVec_hitReq_43_45 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h2D;
  wire          compressDataVec_hitReq_44_45 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h2D;
  wire          compressDataVec_hitReq_45_45 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h2D;
  wire          compressDataVec_hitReq_46_45 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h2D;
  wire          compressDataVec_hitReq_47_45 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h2D;
  wire          compressDataVec_hitReq_48_45 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h2D;
  wire          compressDataVec_hitReq_49_45 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h2D;
  wire          compressDataVec_hitReq_50_45 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h2D;
  wire          compressDataVec_hitReq_51_45 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h2D;
  wire          compressDataVec_hitReq_52_45 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h2D;
  wire          compressDataVec_hitReq_53_45 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h2D;
  wire          compressDataVec_hitReq_54_45 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h2D;
  wire          compressDataVec_hitReq_55_45 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h2D;
  wire          compressDataVec_hitReq_56_45 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h2D;
  wire          compressDataVec_hitReq_57_45 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h2D;
  wire          compressDataVec_hitReq_58_45 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h2D;
  wire          compressDataVec_hitReq_59_45 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h2D;
  wire          compressDataVec_hitReq_60_45 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h2D;
  wire          compressDataVec_hitReq_61_45 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h2D;
  wire          compressDataVec_hitReq_62_45 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h2D;
  wire          compressDataVec_hitReq_63_45 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h2D;
  wire [7:0]    compressDataVec_selectReqData_45 =
    (compressDataVec_hitReq_0_45 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_45 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_45 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_45 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_45 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_45 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_45 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_45 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_45 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_45 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_45 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_45 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_45 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_45 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_45 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_45 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_45 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_45 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_45 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_45 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_45 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_45 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_45 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_45 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_45 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_45 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_45 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_45 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_45 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_45 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_45 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_45 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_45 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_45 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_45 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_45 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_45 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_45 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_45 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_45 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_45 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_45 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_45 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_45 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_45 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_45 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_45 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_45 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_45 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_45 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_45 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_45 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_45 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_45 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_45 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_45 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_45 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_45 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_45 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_45 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_45 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_45 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_45 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_45 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_45 = tailCount > 6'h2D;
  wire          _GEN_1498 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h2E;
  wire          compressDataVec_hitReq_0_46;
  assign compressDataVec_hitReq_0_46 = _GEN_1498;
  wire          compressDataVec_hitReq_0_174;
  assign compressDataVec_hitReq_0_174 = _GEN_1498;
  wire          _GEN_1499 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h2E;
  wire          compressDataVec_hitReq_1_46;
  assign compressDataVec_hitReq_1_46 = _GEN_1499;
  wire          compressDataVec_hitReq_1_174;
  assign compressDataVec_hitReq_1_174 = _GEN_1499;
  wire          _GEN_1500 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h2E;
  wire          compressDataVec_hitReq_2_46;
  assign compressDataVec_hitReq_2_46 = _GEN_1500;
  wire          compressDataVec_hitReq_2_174;
  assign compressDataVec_hitReq_2_174 = _GEN_1500;
  wire          _GEN_1501 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h2E;
  wire          compressDataVec_hitReq_3_46;
  assign compressDataVec_hitReq_3_46 = _GEN_1501;
  wire          compressDataVec_hitReq_3_174;
  assign compressDataVec_hitReq_3_174 = _GEN_1501;
  wire          _GEN_1502 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h2E;
  wire          compressDataVec_hitReq_4_46;
  assign compressDataVec_hitReq_4_46 = _GEN_1502;
  wire          compressDataVec_hitReq_4_174;
  assign compressDataVec_hitReq_4_174 = _GEN_1502;
  wire          _GEN_1503 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h2E;
  wire          compressDataVec_hitReq_5_46;
  assign compressDataVec_hitReq_5_46 = _GEN_1503;
  wire          compressDataVec_hitReq_5_174;
  assign compressDataVec_hitReq_5_174 = _GEN_1503;
  wire          _GEN_1504 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h2E;
  wire          compressDataVec_hitReq_6_46;
  assign compressDataVec_hitReq_6_46 = _GEN_1504;
  wire          compressDataVec_hitReq_6_174;
  assign compressDataVec_hitReq_6_174 = _GEN_1504;
  wire          _GEN_1505 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h2E;
  wire          compressDataVec_hitReq_7_46;
  assign compressDataVec_hitReq_7_46 = _GEN_1505;
  wire          compressDataVec_hitReq_7_174;
  assign compressDataVec_hitReq_7_174 = _GEN_1505;
  wire          _GEN_1506 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h2E;
  wire          compressDataVec_hitReq_8_46;
  assign compressDataVec_hitReq_8_46 = _GEN_1506;
  wire          compressDataVec_hitReq_8_174;
  assign compressDataVec_hitReq_8_174 = _GEN_1506;
  wire          _GEN_1507 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h2E;
  wire          compressDataVec_hitReq_9_46;
  assign compressDataVec_hitReq_9_46 = _GEN_1507;
  wire          compressDataVec_hitReq_9_174;
  assign compressDataVec_hitReq_9_174 = _GEN_1507;
  wire          _GEN_1508 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h2E;
  wire          compressDataVec_hitReq_10_46;
  assign compressDataVec_hitReq_10_46 = _GEN_1508;
  wire          compressDataVec_hitReq_10_174;
  assign compressDataVec_hitReq_10_174 = _GEN_1508;
  wire          _GEN_1509 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h2E;
  wire          compressDataVec_hitReq_11_46;
  assign compressDataVec_hitReq_11_46 = _GEN_1509;
  wire          compressDataVec_hitReq_11_174;
  assign compressDataVec_hitReq_11_174 = _GEN_1509;
  wire          _GEN_1510 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h2E;
  wire          compressDataVec_hitReq_12_46;
  assign compressDataVec_hitReq_12_46 = _GEN_1510;
  wire          compressDataVec_hitReq_12_174;
  assign compressDataVec_hitReq_12_174 = _GEN_1510;
  wire          _GEN_1511 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h2E;
  wire          compressDataVec_hitReq_13_46;
  assign compressDataVec_hitReq_13_46 = _GEN_1511;
  wire          compressDataVec_hitReq_13_174;
  assign compressDataVec_hitReq_13_174 = _GEN_1511;
  wire          _GEN_1512 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h2E;
  wire          compressDataVec_hitReq_14_46;
  assign compressDataVec_hitReq_14_46 = _GEN_1512;
  wire          compressDataVec_hitReq_14_174;
  assign compressDataVec_hitReq_14_174 = _GEN_1512;
  wire          _GEN_1513 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h2E;
  wire          compressDataVec_hitReq_15_46;
  assign compressDataVec_hitReq_15_46 = _GEN_1513;
  wire          compressDataVec_hitReq_15_174;
  assign compressDataVec_hitReq_15_174 = _GEN_1513;
  wire          _GEN_1514 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h2E;
  wire          compressDataVec_hitReq_16_46;
  assign compressDataVec_hitReq_16_46 = _GEN_1514;
  wire          compressDataVec_hitReq_16_174;
  assign compressDataVec_hitReq_16_174 = _GEN_1514;
  wire          _GEN_1515 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h2E;
  wire          compressDataVec_hitReq_17_46;
  assign compressDataVec_hitReq_17_46 = _GEN_1515;
  wire          compressDataVec_hitReq_17_174;
  assign compressDataVec_hitReq_17_174 = _GEN_1515;
  wire          _GEN_1516 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h2E;
  wire          compressDataVec_hitReq_18_46;
  assign compressDataVec_hitReq_18_46 = _GEN_1516;
  wire          compressDataVec_hitReq_18_174;
  assign compressDataVec_hitReq_18_174 = _GEN_1516;
  wire          _GEN_1517 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h2E;
  wire          compressDataVec_hitReq_19_46;
  assign compressDataVec_hitReq_19_46 = _GEN_1517;
  wire          compressDataVec_hitReq_19_174;
  assign compressDataVec_hitReq_19_174 = _GEN_1517;
  wire          _GEN_1518 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h2E;
  wire          compressDataVec_hitReq_20_46;
  assign compressDataVec_hitReq_20_46 = _GEN_1518;
  wire          compressDataVec_hitReq_20_174;
  assign compressDataVec_hitReq_20_174 = _GEN_1518;
  wire          _GEN_1519 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h2E;
  wire          compressDataVec_hitReq_21_46;
  assign compressDataVec_hitReq_21_46 = _GEN_1519;
  wire          compressDataVec_hitReq_21_174;
  assign compressDataVec_hitReq_21_174 = _GEN_1519;
  wire          _GEN_1520 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h2E;
  wire          compressDataVec_hitReq_22_46;
  assign compressDataVec_hitReq_22_46 = _GEN_1520;
  wire          compressDataVec_hitReq_22_174;
  assign compressDataVec_hitReq_22_174 = _GEN_1520;
  wire          _GEN_1521 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h2E;
  wire          compressDataVec_hitReq_23_46;
  assign compressDataVec_hitReq_23_46 = _GEN_1521;
  wire          compressDataVec_hitReq_23_174;
  assign compressDataVec_hitReq_23_174 = _GEN_1521;
  wire          _GEN_1522 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h2E;
  wire          compressDataVec_hitReq_24_46;
  assign compressDataVec_hitReq_24_46 = _GEN_1522;
  wire          compressDataVec_hitReq_24_174;
  assign compressDataVec_hitReq_24_174 = _GEN_1522;
  wire          _GEN_1523 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h2E;
  wire          compressDataVec_hitReq_25_46;
  assign compressDataVec_hitReq_25_46 = _GEN_1523;
  wire          compressDataVec_hitReq_25_174;
  assign compressDataVec_hitReq_25_174 = _GEN_1523;
  wire          _GEN_1524 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h2E;
  wire          compressDataVec_hitReq_26_46;
  assign compressDataVec_hitReq_26_46 = _GEN_1524;
  wire          compressDataVec_hitReq_26_174;
  assign compressDataVec_hitReq_26_174 = _GEN_1524;
  wire          _GEN_1525 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h2E;
  wire          compressDataVec_hitReq_27_46;
  assign compressDataVec_hitReq_27_46 = _GEN_1525;
  wire          compressDataVec_hitReq_27_174;
  assign compressDataVec_hitReq_27_174 = _GEN_1525;
  wire          _GEN_1526 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h2E;
  wire          compressDataVec_hitReq_28_46;
  assign compressDataVec_hitReq_28_46 = _GEN_1526;
  wire          compressDataVec_hitReq_28_174;
  assign compressDataVec_hitReq_28_174 = _GEN_1526;
  wire          _GEN_1527 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h2E;
  wire          compressDataVec_hitReq_29_46;
  assign compressDataVec_hitReq_29_46 = _GEN_1527;
  wire          compressDataVec_hitReq_29_174;
  assign compressDataVec_hitReq_29_174 = _GEN_1527;
  wire          _GEN_1528 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h2E;
  wire          compressDataVec_hitReq_30_46;
  assign compressDataVec_hitReq_30_46 = _GEN_1528;
  wire          compressDataVec_hitReq_30_174;
  assign compressDataVec_hitReq_30_174 = _GEN_1528;
  wire          _GEN_1529 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h2E;
  wire          compressDataVec_hitReq_31_46;
  assign compressDataVec_hitReq_31_46 = _GEN_1529;
  wire          compressDataVec_hitReq_31_174;
  assign compressDataVec_hitReq_31_174 = _GEN_1529;
  wire          compressDataVec_hitReq_32_46 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h2E;
  wire          compressDataVec_hitReq_33_46 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h2E;
  wire          compressDataVec_hitReq_34_46 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h2E;
  wire          compressDataVec_hitReq_35_46 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h2E;
  wire          compressDataVec_hitReq_36_46 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h2E;
  wire          compressDataVec_hitReq_37_46 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h2E;
  wire          compressDataVec_hitReq_38_46 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h2E;
  wire          compressDataVec_hitReq_39_46 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h2E;
  wire          compressDataVec_hitReq_40_46 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h2E;
  wire          compressDataVec_hitReq_41_46 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h2E;
  wire          compressDataVec_hitReq_42_46 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h2E;
  wire          compressDataVec_hitReq_43_46 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h2E;
  wire          compressDataVec_hitReq_44_46 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h2E;
  wire          compressDataVec_hitReq_45_46 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h2E;
  wire          compressDataVec_hitReq_46_46 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h2E;
  wire          compressDataVec_hitReq_47_46 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h2E;
  wire          compressDataVec_hitReq_48_46 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h2E;
  wire          compressDataVec_hitReq_49_46 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h2E;
  wire          compressDataVec_hitReq_50_46 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h2E;
  wire          compressDataVec_hitReq_51_46 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h2E;
  wire          compressDataVec_hitReq_52_46 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h2E;
  wire          compressDataVec_hitReq_53_46 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h2E;
  wire          compressDataVec_hitReq_54_46 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h2E;
  wire          compressDataVec_hitReq_55_46 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h2E;
  wire          compressDataVec_hitReq_56_46 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h2E;
  wire          compressDataVec_hitReq_57_46 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h2E;
  wire          compressDataVec_hitReq_58_46 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h2E;
  wire          compressDataVec_hitReq_59_46 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h2E;
  wire          compressDataVec_hitReq_60_46 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h2E;
  wire          compressDataVec_hitReq_61_46 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h2E;
  wire          compressDataVec_hitReq_62_46 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h2E;
  wire          compressDataVec_hitReq_63_46 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h2E;
  wire [7:0]    compressDataVec_selectReqData_46 =
    (compressDataVec_hitReq_0_46 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_46 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_46 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_46 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_46 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_46 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_46 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_46 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_46 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_46 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_46 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_46 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_46 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_46 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_46 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_46 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_46 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_46 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_46 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_46 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_46 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_46 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_46 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_46 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_46 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_46 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_46 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_46 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_46 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_46 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_46 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_46 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_46 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_46 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_46 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_46 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_46 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_46 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_46 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_46 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_46 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_46 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_46 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_46 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_46 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_46 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_46 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_46 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_46 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_46 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_46 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_46 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_46 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_46 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_46 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_46 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_46 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_46 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_46 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_46 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_46 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_46 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_46 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_46 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_46 = tailCount > 6'h2E;
  wire          _GEN_1530 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h2F;
  wire          compressDataVec_hitReq_0_47;
  assign compressDataVec_hitReq_0_47 = _GEN_1530;
  wire          compressDataVec_hitReq_0_175;
  assign compressDataVec_hitReq_0_175 = _GEN_1530;
  wire          _GEN_1531 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h2F;
  wire          compressDataVec_hitReq_1_47;
  assign compressDataVec_hitReq_1_47 = _GEN_1531;
  wire          compressDataVec_hitReq_1_175;
  assign compressDataVec_hitReq_1_175 = _GEN_1531;
  wire          _GEN_1532 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h2F;
  wire          compressDataVec_hitReq_2_47;
  assign compressDataVec_hitReq_2_47 = _GEN_1532;
  wire          compressDataVec_hitReq_2_175;
  assign compressDataVec_hitReq_2_175 = _GEN_1532;
  wire          _GEN_1533 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h2F;
  wire          compressDataVec_hitReq_3_47;
  assign compressDataVec_hitReq_3_47 = _GEN_1533;
  wire          compressDataVec_hitReq_3_175;
  assign compressDataVec_hitReq_3_175 = _GEN_1533;
  wire          _GEN_1534 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h2F;
  wire          compressDataVec_hitReq_4_47;
  assign compressDataVec_hitReq_4_47 = _GEN_1534;
  wire          compressDataVec_hitReq_4_175;
  assign compressDataVec_hitReq_4_175 = _GEN_1534;
  wire          _GEN_1535 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h2F;
  wire          compressDataVec_hitReq_5_47;
  assign compressDataVec_hitReq_5_47 = _GEN_1535;
  wire          compressDataVec_hitReq_5_175;
  assign compressDataVec_hitReq_5_175 = _GEN_1535;
  wire          _GEN_1536 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h2F;
  wire          compressDataVec_hitReq_6_47;
  assign compressDataVec_hitReq_6_47 = _GEN_1536;
  wire          compressDataVec_hitReq_6_175;
  assign compressDataVec_hitReq_6_175 = _GEN_1536;
  wire          _GEN_1537 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h2F;
  wire          compressDataVec_hitReq_7_47;
  assign compressDataVec_hitReq_7_47 = _GEN_1537;
  wire          compressDataVec_hitReq_7_175;
  assign compressDataVec_hitReq_7_175 = _GEN_1537;
  wire          _GEN_1538 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h2F;
  wire          compressDataVec_hitReq_8_47;
  assign compressDataVec_hitReq_8_47 = _GEN_1538;
  wire          compressDataVec_hitReq_8_175;
  assign compressDataVec_hitReq_8_175 = _GEN_1538;
  wire          _GEN_1539 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h2F;
  wire          compressDataVec_hitReq_9_47;
  assign compressDataVec_hitReq_9_47 = _GEN_1539;
  wire          compressDataVec_hitReq_9_175;
  assign compressDataVec_hitReq_9_175 = _GEN_1539;
  wire          _GEN_1540 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h2F;
  wire          compressDataVec_hitReq_10_47;
  assign compressDataVec_hitReq_10_47 = _GEN_1540;
  wire          compressDataVec_hitReq_10_175;
  assign compressDataVec_hitReq_10_175 = _GEN_1540;
  wire          _GEN_1541 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h2F;
  wire          compressDataVec_hitReq_11_47;
  assign compressDataVec_hitReq_11_47 = _GEN_1541;
  wire          compressDataVec_hitReq_11_175;
  assign compressDataVec_hitReq_11_175 = _GEN_1541;
  wire          _GEN_1542 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h2F;
  wire          compressDataVec_hitReq_12_47;
  assign compressDataVec_hitReq_12_47 = _GEN_1542;
  wire          compressDataVec_hitReq_12_175;
  assign compressDataVec_hitReq_12_175 = _GEN_1542;
  wire          _GEN_1543 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h2F;
  wire          compressDataVec_hitReq_13_47;
  assign compressDataVec_hitReq_13_47 = _GEN_1543;
  wire          compressDataVec_hitReq_13_175;
  assign compressDataVec_hitReq_13_175 = _GEN_1543;
  wire          _GEN_1544 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h2F;
  wire          compressDataVec_hitReq_14_47;
  assign compressDataVec_hitReq_14_47 = _GEN_1544;
  wire          compressDataVec_hitReq_14_175;
  assign compressDataVec_hitReq_14_175 = _GEN_1544;
  wire          _GEN_1545 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h2F;
  wire          compressDataVec_hitReq_15_47;
  assign compressDataVec_hitReq_15_47 = _GEN_1545;
  wire          compressDataVec_hitReq_15_175;
  assign compressDataVec_hitReq_15_175 = _GEN_1545;
  wire          _GEN_1546 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h2F;
  wire          compressDataVec_hitReq_16_47;
  assign compressDataVec_hitReq_16_47 = _GEN_1546;
  wire          compressDataVec_hitReq_16_175;
  assign compressDataVec_hitReq_16_175 = _GEN_1546;
  wire          _GEN_1547 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h2F;
  wire          compressDataVec_hitReq_17_47;
  assign compressDataVec_hitReq_17_47 = _GEN_1547;
  wire          compressDataVec_hitReq_17_175;
  assign compressDataVec_hitReq_17_175 = _GEN_1547;
  wire          _GEN_1548 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h2F;
  wire          compressDataVec_hitReq_18_47;
  assign compressDataVec_hitReq_18_47 = _GEN_1548;
  wire          compressDataVec_hitReq_18_175;
  assign compressDataVec_hitReq_18_175 = _GEN_1548;
  wire          _GEN_1549 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h2F;
  wire          compressDataVec_hitReq_19_47;
  assign compressDataVec_hitReq_19_47 = _GEN_1549;
  wire          compressDataVec_hitReq_19_175;
  assign compressDataVec_hitReq_19_175 = _GEN_1549;
  wire          _GEN_1550 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h2F;
  wire          compressDataVec_hitReq_20_47;
  assign compressDataVec_hitReq_20_47 = _GEN_1550;
  wire          compressDataVec_hitReq_20_175;
  assign compressDataVec_hitReq_20_175 = _GEN_1550;
  wire          _GEN_1551 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h2F;
  wire          compressDataVec_hitReq_21_47;
  assign compressDataVec_hitReq_21_47 = _GEN_1551;
  wire          compressDataVec_hitReq_21_175;
  assign compressDataVec_hitReq_21_175 = _GEN_1551;
  wire          _GEN_1552 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h2F;
  wire          compressDataVec_hitReq_22_47;
  assign compressDataVec_hitReq_22_47 = _GEN_1552;
  wire          compressDataVec_hitReq_22_175;
  assign compressDataVec_hitReq_22_175 = _GEN_1552;
  wire          _GEN_1553 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h2F;
  wire          compressDataVec_hitReq_23_47;
  assign compressDataVec_hitReq_23_47 = _GEN_1553;
  wire          compressDataVec_hitReq_23_175;
  assign compressDataVec_hitReq_23_175 = _GEN_1553;
  wire          _GEN_1554 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h2F;
  wire          compressDataVec_hitReq_24_47;
  assign compressDataVec_hitReq_24_47 = _GEN_1554;
  wire          compressDataVec_hitReq_24_175;
  assign compressDataVec_hitReq_24_175 = _GEN_1554;
  wire          _GEN_1555 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h2F;
  wire          compressDataVec_hitReq_25_47;
  assign compressDataVec_hitReq_25_47 = _GEN_1555;
  wire          compressDataVec_hitReq_25_175;
  assign compressDataVec_hitReq_25_175 = _GEN_1555;
  wire          _GEN_1556 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h2F;
  wire          compressDataVec_hitReq_26_47;
  assign compressDataVec_hitReq_26_47 = _GEN_1556;
  wire          compressDataVec_hitReq_26_175;
  assign compressDataVec_hitReq_26_175 = _GEN_1556;
  wire          _GEN_1557 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h2F;
  wire          compressDataVec_hitReq_27_47;
  assign compressDataVec_hitReq_27_47 = _GEN_1557;
  wire          compressDataVec_hitReq_27_175;
  assign compressDataVec_hitReq_27_175 = _GEN_1557;
  wire          _GEN_1558 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h2F;
  wire          compressDataVec_hitReq_28_47;
  assign compressDataVec_hitReq_28_47 = _GEN_1558;
  wire          compressDataVec_hitReq_28_175;
  assign compressDataVec_hitReq_28_175 = _GEN_1558;
  wire          _GEN_1559 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h2F;
  wire          compressDataVec_hitReq_29_47;
  assign compressDataVec_hitReq_29_47 = _GEN_1559;
  wire          compressDataVec_hitReq_29_175;
  assign compressDataVec_hitReq_29_175 = _GEN_1559;
  wire          _GEN_1560 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h2F;
  wire          compressDataVec_hitReq_30_47;
  assign compressDataVec_hitReq_30_47 = _GEN_1560;
  wire          compressDataVec_hitReq_30_175;
  assign compressDataVec_hitReq_30_175 = _GEN_1560;
  wire          _GEN_1561 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h2F;
  wire          compressDataVec_hitReq_31_47;
  assign compressDataVec_hitReq_31_47 = _GEN_1561;
  wire          compressDataVec_hitReq_31_175;
  assign compressDataVec_hitReq_31_175 = _GEN_1561;
  wire          compressDataVec_hitReq_32_47 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h2F;
  wire          compressDataVec_hitReq_33_47 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h2F;
  wire          compressDataVec_hitReq_34_47 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h2F;
  wire          compressDataVec_hitReq_35_47 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h2F;
  wire          compressDataVec_hitReq_36_47 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h2F;
  wire          compressDataVec_hitReq_37_47 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h2F;
  wire          compressDataVec_hitReq_38_47 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h2F;
  wire          compressDataVec_hitReq_39_47 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h2F;
  wire          compressDataVec_hitReq_40_47 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h2F;
  wire          compressDataVec_hitReq_41_47 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h2F;
  wire          compressDataVec_hitReq_42_47 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h2F;
  wire          compressDataVec_hitReq_43_47 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h2F;
  wire          compressDataVec_hitReq_44_47 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h2F;
  wire          compressDataVec_hitReq_45_47 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h2F;
  wire          compressDataVec_hitReq_46_47 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h2F;
  wire          compressDataVec_hitReq_47_47 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h2F;
  wire          compressDataVec_hitReq_48_47 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h2F;
  wire          compressDataVec_hitReq_49_47 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h2F;
  wire          compressDataVec_hitReq_50_47 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h2F;
  wire          compressDataVec_hitReq_51_47 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h2F;
  wire          compressDataVec_hitReq_52_47 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h2F;
  wire          compressDataVec_hitReq_53_47 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h2F;
  wire          compressDataVec_hitReq_54_47 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h2F;
  wire          compressDataVec_hitReq_55_47 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h2F;
  wire          compressDataVec_hitReq_56_47 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h2F;
  wire          compressDataVec_hitReq_57_47 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h2F;
  wire          compressDataVec_hitReq_58_47 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h2F;
  wire          compressDataVec_hitReq_59_47 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h2F;
  wire          compressDataVec_hitReq_60_47 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h2F;
  wire          compressDataVec_hitReq_61_47 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h2F;
  wire          compressDataVec_hitReq_62_47 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h2F;
  wire          compressDataVec_hitReq_63_47 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h2F;
  wire [7:0]    compressDataVec_selectReqData_47 =
    (compressDataVec_hitReq_0_47 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_47 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_47 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_47 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_47 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_47 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_47 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_47 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_47 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_47 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_47 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_47 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_47 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_47 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_47 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_47 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_47 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_47 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_47 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_47 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_47 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_47 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_47 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_47 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_47 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_47 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_47 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_47 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_47 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_47 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_47 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_47 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_47 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_47 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_47 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_47 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_47 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_47 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_47 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_47 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_47 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_47 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_47 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_47 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_47 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_47 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_47 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_47 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_47 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_47 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_47 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_47 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_47 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_47 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_47 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_47 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_47 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_47 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_47 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_47 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_47 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_47 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_47 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_47 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_47 = tailCount > 6'h2F;
  wire          _GEN_1562 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h30;
  wire          compressDataVec_hitReq_0_48;
  assign compressDataVec_hitReq_0_48 = _GEN_1562;
  wire          compressDataVec_hitReq_0_176;
  assign compressDataVec_hitReq_0_176 = _GEN_1562;
  wire          _GEN_1563 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h30;
  wire          compressDataVec_hitReq_1_48;
  assign compressDataVec_hitReq_1_48 = _GEN_1563;
  wire          compressDataVec_hitReq_1_176;
  assign compressDataVec_hitReq_1_176 = _GEN_1563;
  wire          _GEN_1564 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h30;
  wire          compressDataVec_hitReq_2_48;
  assign compressDataVec_hitReq_2_48 = _GEN_1564;
  wire          compressDataVec_hitReq_2_176;
  assign compressDataVec_hitReq_2_176 = _GEN_1564;
  wire          _GEN_1565 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h30;
  wire          compressDataVec_hitReq_3_48;
  assign compressDataVec_hitReq_3_48 = _GEN_1565;
  wire          compressDataVec_hitReq_3_176;
  assign compressDataVec_hitReq_3_176 = _GEN_1565;
  wire          _GEN_1566 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h30;
  wire          compressDataVec_hitReq_4_48;
  assign compressDataVec_hitReq_4_48 = _GEN_1566;
  wire          compressDataVec_hitReq_4_176;
  assign compressDataVec_hitReq_4_176 = _GEN_1566;
  wire          _GEN_1567 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h30;
  wire          compressDataVec_hitReq_5_48;
  assign compressDataVec_hitReq_5_48 = _GEN_1567;
  wire          compressDataVec_hitReq_5_176;
  assign compressDataVec_hitReq_5_176 = _GEN_1567;
  wire          _GEN_1568 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h30;
  wire          compressDataVec_hitReq_6_48;
  assign compressDataVec_hitReq_6_48 = _GEN_1568;
  wire          compressDataVec_hitReq_6_176;
  assign compressDataVec_hitReq_6_176 = _GEN_1568;
  wire          _GEN_1569 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h30;
  wire          compressDataVec_hitReq_7_48;
  assign compressDataVec_hitReq_7_48 = _GEN_1569;
  wire          compressDataVec_hitReq_7_176;
  assign compressDataVec_hitReq_7_176 = _GEN_1569;
  wire          _GEN_1570 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h30;
  wire          compressDataVec_hitReq_8_48;
  assign compressDataVec_hitReq_8_48 = _GEN_1570;
  wire          compressDataVec_hitReq_8_176;
  assign compressDataVec_hitReq_8_176 = _GEN_1570;
  wire          _GEN_1571 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h30;
  wire          compressDataVec_hitReq_9_48;
  assign compressDataVec_hitReq_9_48 = _GEN_1571;
  wire          compressDataVec_hitReq_9_176;
  assign compressDataVec_hitReq_9_176 = _GEN_1571;
  wire          _GEN_1572 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h30;
  wire          compressDataVec_hitReq_10_48;
  assign compressDataVec_hitReq_10_48 = _GEN_1572;
  wire          compressDataVec_hitReq_10_176;
  assign compressDataVec_hitReq_10_176 = _GEN_1572;
  wire          _GEN_1573 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h30;
  wire          compressDataVec_hitReq_11_48;
  assign compressDataVec_hitReq_11_48 = _GEN_1573;
  wire          compressDataVec_hitReq_11_176;
  assign compressDataVec_hitReq_11_176 = _GEN_1573;
  wire          _GEN_1574 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h30;
  wire          compressDataVec_hitReq_12_48;
  assign compressDataVec_hitReq_12_48 = _GEN_1574;
  wire          compressDataVec_hitReq_12_176;
  assign compressDataVec_hitReq_12_176 = _GEN_1574;
  wire          _GEN_1575 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h30;
  wire          compressDataVec_hitReq_13_48;
  assign compressDataVec_hitReq_13_48 = _GEN_1575;
  wire          compressDataVec_hitReq_13_176;
  assign compressDataVec_hitReq_13_176 = _GEN_1575;
  wire          _GEN_1576 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h30;
  wire          compressDataVec_hitReq_14_48;
  assign compressDataVec_hitReq_14_48 = _GEN_1576;
  wire          compressDataVec_hitReq_14_176;
  assign compressDataVec_hitReq_14_176 = _GEN_1576;
  wire          _GEN_1577 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h30;
  wire          compressDataVec_hitReq_15_48;
  assign compressDataVec_hitReq_15_48 = _GEN_1577;
  wire          compressDataVec_hitReq_15_176;
  assign compressDataVec_hitReq_15_176 = _GEN_1577;
  wire          _GEN_1578 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h30;
  wire          compressDataVec_hitReq_16_48;
  assign compressDataVec_hitReq_16_48 = _GEN_1578;
  wire          compressDataVec_hitReq_16_176;
  assign compressDataVec_hitReq_16_176 = _GEN_1578;
  wire          _GEN_1579 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h30;
  wire          compressDataVec_hitReq_17_48;
  assign compressDataVec_hitReq_17_48 = _GEN_1579;
  wire          compressDataVec_hitReq_17_176;
  assign compressDataVec_hitReq_17_176 = _GEN_1579;
  wire          _GEN_1580 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h30;
  wire          compressDataVec_hitReq_18_48;
  assign compressDataVec_hitReq_18_48 = _GEN_1580;
  wire          compressDataVec_hitReq_18_176;
  assign compressDataVec_hitReq_18_176 = _GEN_1580;
  wire          _GEN_1581 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h30;
  wire          compressDataVec_hitReq_19_48;
  assign compressDataVec_hitReq_19_48 = _GEN_1581;
  wire          compressDataVec_hitReq_19_176;
  assign compressDataVec_hitReq_19_176 = _GEN_1581;
  wire          _GEN_1582 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h30;
  wire          compressDataVec_hitReq_20_48;
  assign compressDataVec_hitReq_20_48 = _GEN_1582;
  wire          compressDataVec_hitReq_20_176;
  assign compressDataVec_hitReq_20_176 = _GEN_1582;
  wire          _GEN_1583 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h30;
  wire          compressDataVec_hitReq_21_48;
  assign compressDataVec_hitReq_21_48 = _GEN_1583;
  wire          compressDataVec_hitReq_21_176;
  assign compressDataVec_hitReq_21_176 = _GEN_1583;
  wire          _GEN_1584 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h30;
  wire          compressDataVec_hitReq_22_48;
  assign compressDataVec_hitReq_22_48 = _GEN_1584;
  wire          compressDataVec_hitReq_22_176;
  assign compressDataVec_hitReq_22_176 = _GEN_1584;
  wire          _GEN_1585 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h30;
  wire          compressDataVec_hitReq_23_48;
  assign compressDataVec_hitReq_23_48 = _GEN_1585;
  wire          compressDataVec_hitReq_23_176;
  assign compressDataVec_hitReq_23_176 = _GEN_1585;
  wire          _GEN_1586 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h30;
  wire          compressDataVec_hitReq_24_48;
  assign compressDataVec_hitReq_24_48 = _GEN_1586;
  wire          compressDataVec_hitReq_24_176;
  assign compressDataVec_hitReq_24_176 = _GEN_1586;
  wire          _GEN_1587 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h30;
  wire          compressDataVec_hitReq_25_48;
  assign compressDataVec_hitReq_25_48 = _GEN_1587;
  wire          compressDataVec_hitReq_25_176;
  assign compressDataVec_hitReq_25_176 = _GEN_1587;
  wire          _GEN_1588 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h30;
  wire          compressDataVec_hitReq_26_48;
  assign compressDataVec_hitReq_26_48 = _GEN_1588;
  wire          compressDataVec_hitReq_26_176;
  assign compressDataVec_hitReq_26_176 = _GEN_1588;
  wire          _GEN_1589 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h30;
  wire          compressDataVec_hitReq_27_48;
  assign compressDataVec_hitReq_27_48 = _GEN_1589;
  wire          compressDataVec_hitReq_27_176;
  assign compressDataVec_hitReq_27_176 = _GEN_1589;
  wire          _GEN_1590 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h30;
  wire          compressDataVec_hitReq_28_48;
  assign compressDataVec_hitReq_28_48 = _GEN_1590;
  wire          compressDataVec_hitReq_28_176;
  assign compressDataVec_hitReq_28_176 = _GEN_1590;
  wire          _GEN_1591 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h30;
  wire          compressDataVec_hitReq_29_48;
  assign compressDataVec_hitReq_29_48 = _GEN_1591;
  wire          compressDataVec_hitReq_29_176;
  assign compressDataVec_hitReq_29_176 = _GEN_1591;
  wire          _GEN_1592 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h30;
  wire          compressDataVec_hitReq_30_48;
  assign compressDataVec_hitReq_30_48 = _GEN_1592;
  wire          compressDataVec_hitReq_30_176;
  assign compressDataVec_hitReq_30_176 = _GEN_1592;
  wire          _GEN_1593 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h30;
  wire          compressDataVec_hitReq_31_48;
  assign compressDataVec_hitReq_31_48 = _GEN_1593;
  wire          compressDataVec_hitReq_31_176;
  assign compressDataVec_hitReq_31_176 = _GEN_1593;
  wire          compressDataVec_hitReq_32_48 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h30;
  wire          compressDataVec_hitReq_33_48 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h30;
  wire          compressDataVec_hitReq_34_48 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h30;
  wire          compressDataVec_hitReq_35_48 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h30;
  wire          compressDataVec_hitReq_36_48 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h30;
  wire          compressDataVec_hitReq_37_48 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h30;
  wire          compressDataVec_hitReq_38_48 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h30;
  wire          compressDataVec_hitReq_39_48 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h30;
  wire          compressDataVec_hitReq_40_48 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h30;
  wire          compressDataVec_hitReq_41_48 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h30;
  wire          compressDataVec_hitReq_42_48 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h30;
  wire          compressDataVec_hitReq_43_48 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h30;
  wire          compressDataVec_hitReq_44_48 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h30;
  wire          compressDataVec_hitReq_45_48 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h30;
  wire          compressDataVec_hitReq_46_48 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h30;
  wire          compressDataVec_hitReq_47_48 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h30;
  wire          compressDataVec_hitReq_48_48 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h30;
  wire          compressDataVec_hitReq_49_48 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h30;
  wire          compressDataVec_hitReq_50_48 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h30;
  wire          compressDataVec_hitReq_51_48 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h30;
  wire          compressDataVec_hitReq_52_48 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h30;
  wire          compressDataVec_hitReq_53_48 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h30;
  wire          compressDataVec_hitReq_54_48 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h30;
  wire          compressDataVec_hitReq_55_48 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h30;
  wire          compressDataVec_hitReq_56_48 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h30;
  wire          compressDataVec_hitReq_57_48 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h30;
  wire          compressDataVec_hitReq_58_48 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h30;
  wire          compressDataVec_hitReq_59_48 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h30;
  wire          compressDataVec_hitReq_60_48 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h30;
  wire          compressDataVec_hitReq_61_48 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h30;
  wire          compressDataVec_hitReq_62_48 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h30;
  wire          compressDataVec_hitReq_63_48 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h30;
  wire [7:0]    compressDataVec_selectReqData_48 =
    (compressDataVec_hitReq_0_48 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_48 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_48 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_48 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_48 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_48 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_48 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_48 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_48 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_48 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_48 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_48 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_48 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_48 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_48 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_48 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_48 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_48 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_48 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_48 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_48 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_48 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_48 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_48 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_48 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_48 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_48 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_48 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_48 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_48 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_48 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_48 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_48 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_48 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_48 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_48 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_48 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_48 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_48 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_48 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_48 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_48 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_48 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_48 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_48 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_48 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_48 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_48 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_48 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_48 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_48 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_48 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_48 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_48 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_48 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_48 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_48 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_48 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_48 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_48 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_48 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_48 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_48 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_48 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_48 = tailCount > 6'h30;
  wire          _GEN_1594 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h31;
  wire          compressDataVec_hitReq_0_49;
  assign compressDataVec_hitReq_0_49 = _GEN_1594;
  wire          compressDataVec_hitReq_0_177;
  assign compressDataVec_hitReq_0_177 = _GEN_1594;
  wire          _GEN_1595 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h31;
  wire          compressDataVec_hitReq_1_49;
  assign compressDataVec_hitReq_1_49 = _GEN_1595;
  wire          compressDataVec_hitReq_1_177;
  assign compressDataVec_hitReq_1_177 = _GEN_1595;
  wire          _GEN_1596 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h31;
  wire          compressDataVec_hitReq_2_49;
  assign compressDataVec_hitReq_2_49 = _GEN_1596;
  wire          compressDataVec_hitReq_2_177;
  assign compressDataVec_hitReq_2_177 = _GEN_1596;
  wire          _GEN_1597 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h31;
  wire          compressDataVec_hitReq_3_49;
  assign compressDataVec_hitReq_3_49 = _GEN_1597;
  wire          compressDataVec_hitReq_3_177;
  assign compressDataVec_hitReq_3_177 = _GEN_1597;
  wire          _GEN_1598 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h31;
  wire          compressDataVec_hitReq_4_49;
  assign compressDataVec_hitReq_4_49 = _GEN_1598;
  wire          compressDataVec_hitReq_4_177;
  assign compressDataVec_hitReq_4_177 = _GEN_1598;
  wire          _GEN_1599 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h31;
  wire          compressDataVec_hitReq_5_49;
  assign compressDataVec_hitReq_5_49 = _GEN_1599;
  wire          compressDataVec_hitReq_5_177;
  assign compressDataVec_hitReq_5_177 = _GEN_1599;
  wire          _GEN_1600 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h31;
  wire          compressDataVec_hitReq_6_49;
  assign compressDataVec_hitReq_6_49 = _GEN_1600;
  wire          compressDataVec_hitReq_6_177;
  assign compressDataVec_hitReq_6_177 = _GEN_1600;
  wire          _GEN_1601 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h31;
  wire          compressDataVec_hitReq_7_49;
  assign compressDataVec_hitReq_7_49 = _GEN_1601;
  wire          compressDataVec_hitReq_7_177;
  assign compressDataVec_hitReq_7_177 = _GEN_1601;
  wire          _GEN_1602 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h31;
  wire          compressDataVec_hitReq_8_49;
  assign compressDataVec_hitReq_8_49 = _GEN_1602;
  wire          compressDataVec_hitReq_8_177;
  assign compressDataVec_hitReq_8_177 = _GEN_1602;
  wire          _GEN_1603 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h31;
  wire          compressDataVec_hitReq_9_49;
  assign compressDataVec_hitReq_9_49 = _GEN_1603;
  wire          compressDataVec_hitReq_9_177;
  assign compressDataVec_hitReq_9_177 = _GEN_1603;
  wire          _GEN_1604 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h31;
  wire          compressDataVec_hitReq_10_49;
  assign compressDataVec_hitReq_10_49 = _GEN_1604;
  wire          compressDataVec_hitReq_10_177;
  assign compressDataVec_hitReq_10_177 = _GEN_1604;
  wire          _GEN_1605 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h31;
  wire          compressDataVec_hitReq_11_49;
  assign compressDataVec_hitReq_11_49 = _GEN_1605;
  wire          compressDataVec_hitReq_11_177;
  assign compressDataVec_hitReq_11_177 = _GEN_1605;
  wire          _GEN_1606 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h31;
  wire          compressDataVec_hitReq_12_49;
  assign compressDataVec_hitReq_12_49 = _GEN_1606;
  wire          compressDataVec_hitReq_12_177;
  assign compressDataVec_hitReq_12_177 = _GEN_1606;
  wire          _GEN_1607 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h31;
  wire          compressDataVec_hitReq_13_49;
  assign compressDataVec_hitReq_13_49 = _GEN_1607;
  wire          compressDataVec_hitReq_13_177;
  assign compressDataVec_hitReq_13_177 = _GEN_1607;
  wire          _GEN_1608 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h31;
  wire          compressDataVec_hitReq_14_49;
  assign compressDataVec_hitReq_14_49 = _GEN_1608;
  wire          compressDataVec_hitReq_14_177;
  assign compressDataVec_hitReq_14_177 = _GEN_1608;
  wire          _GEN_1609 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h31;
  wire          compressDataVec_hitReq_15_49;
  assign compressDataVec_hitReq_15_49 = _GEN_1609;
  wire          compressDataVec_hitReq_15_177;
  assign compressDataVec_hitReq_15_177 = _GEN_1609;
  wire          _GEN_1610 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h31;
  wire          compressDataVec_hitReq_16_49;
  assign compressDataVec_hitReq_16_49 = _GEN_1610;
  wire          compressDataVec_hitReq_16_177;
  assign compressDataVec_hitReq_16_177 = _GEN_1610;
  wire          _GEN_1611 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h31;
  wire          compressDataVec_hitReq_17_49;
  assign compressDataVec_hitReq_17_49 = _GEN_1611;
  wire          compressDataVec_hitReq_17_177;
  assign compressDataVec_hitReq_17_177 = _GEN_1611;
  wire          _GEN_1612 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h31;
  wire          compressDataVec_hitReq_18_49;
  assign compressDataVec_hitReq_18_49 = _GEN_1612;
  wire          compressDataVec_hitReq_18_177;
  assign compressDataVec_hitReq_18_177 = _GEN_1612;
  wire          _GEN_1613 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h31;
  wire          compressDataVec_hitReq_19_49;
  assign compressDataVec_hitReq_19_49 = _GEN_1613;
  wire          compressDataVec_hitReq_19_177;
  assign compressDataVec_hitReq_19_177 = _GEN_1613;
  wire          _GEN_1614 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h31;
  wire          compressDataVec_hitReq_20_49;
  assign compressDataVec_hitReq_20_49 = _GEN_1614;
  wire          compressDataVec_hitReq_20_177;
  assign compressDataVec_hitReq_20_177 = _GEN_1614;
  wire          _GEN_1615 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h31;
  wire          compressDataVec_hitReq_21_49;
  assign compressDataVec_hitReq_21_49 = _GEN_1615;
  wire          compressDataVec_hitReq_21_177;
  assign compressDataVec_hitReq_21_177 = _GEN_1615;
  wire          _GEN_1616 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h31;
  wire          compressDataVec_hitReq_22_49;
  assign compressDataVec_hitReq_22_49 = _GEN_1616;
  wire          compressDataVec_hitReq_22_177;
  assign compressDataVec_hitReq_22_177 = _GEN_1616;
  wire          _GEN_1617 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h31;
  wire          compressDataVec_hitReq_23_49;
  assign compressDataVec_hitReq_23_49 = _GEN_1617;
  wire          compressDataVec_hitReq_23_177;
  assign compressDataVec_hitReq_23_177 = _GEN_1617;
  wire          _GEN_1618 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h31;
  wire          compressDataVec_hitReq_24_49;
  assign compressDataVec_hitReq_24_49 = _GEN_1618;
  wire          compressDataVec_hitReq_24_177;
  assign compressDataVec_hitReq_24_177 = _GEN_1618;
  wire          _GEN_1619 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h31;
  wire          compressDataVec_hitReq_25_49;
  assign compressDataVec_hitReq_25_49 = _GEN_1619;
  wire          compressDataVec_hitReq_25_177;
  assign compressDataVec_hitReq_25_177 = _GEN_1619;
  wire          _GEN_1620 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h31;
  wire          compressDataVec_hitReq_26_49;
  assign compressDataVec_hitReq_26_49 = _GEN_1620;
  wire          compressDataVec_hitReq_26_177;
  assign compressDataVec_hitReq_26_177 = _GEN_1620;
  wire          _GEN_1621 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h31;
  wire          compressDataVec_hitReq_27_49;
  assign compressDataVec_hitReq_27_49 = _GEN_1621;
  wire          compressDataVec_hitReq_27_177;
  assign compressDataVec_hitReq_27_177 = _GEN_1621;
  wire          _GEN_1622 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h31;
  wire          compressDataVec_hitReq_28_49;
  assign compressDataVec_hitReq_28_49 = _GEN_1622;
  wire          compressDataVec_hitReq_28_177;
  assign compressDataVec_hitReq_28_177 = _GEN_1622;
  wire          _GEN_1623 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h31;
  wire          compressDataVec_hitReq_29_49;
  assign compressDataVec_hitReq_29_49 = _GEN_1623;
  wire          compressDataVec_hitReq_29_177;
  assign compressDataVec_hitReq_29_177 = _GEN_1623;
  wire          _GEN_1624 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h31;
  wire          compressDataVec_hitReq_30_49;
  assign compressDataVec_hitReq_30_49 = _GEN_1624;
  wire          compressDataVec_hitReq_30_177;
  assign compressDataVec_hitReq_30_177 = _GEN_1624;
  wire          _GEN_1625 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h31;
  wire          compressDataVec_hitReq_31_49;
  assign compressDataVec_hitReq_31_49 = _GEN_1625;
  wire          compressDataVec_hitReq_31_177;
  assign compressDataVec_hitReq_31_177 = _GEN_1625;
  wire          compressDataVec_hitReq_32_49 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h31;
  wire          compressDataVec_hitReq_33_49 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h31;
  wire          compressDataVec_hitReq_34_49 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h31;
  wire          compressDataVec_hitReq_35_49 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h31;
  wire          compressDataVec_hitReq_36_49 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h31;
  wire          compressDataVec_hitReq_37_49 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h31;
  wire          compressDataVec_hitReq_38_49 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h31;
  wire          compressDataVec_hitReq_39_49 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h31;
  wire          compressDataVec_hitReq_40_49 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h31;
  wire          compressDataVec_hitReq_41_49 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h31;
  wire          compressDataVec_hitReq_42_49 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h31;
  wire          compressDataVec_hitReq_43_49 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h31;
  wire          compressDataVec_hitReq_44_49 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h31;
  wire          compressDataVec_hitReq_45_49 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h31;
  wire          compressDataVec_hitReq_46_49 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h31;
  wire          compressDataVec_hitReq_47_49 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h31;
  wire          compressDataVec_hitReq_48_49 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h31;
  wire          compressDataVec_hitReq_49_49 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h31;
  wire          compressDataVec_hitReq_50_49 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h31;
  wire          compressDataVec_hitReq_51_49 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h31;
  wire          compressDataVec_hitReq_52_49 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h31;
  wire          compressDataVec_hitReq_53_49 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h31;
  wire          compressDataVec_hitReq_54_49 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h31;
  wire          compressDataVec_hitReq_55_49 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h31;
  wire          compressDataVec_hitReq_56_49 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h31;
  wire          compressDataVec_hitReq_57_49 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h31;
  wire          compressDataVec_hitReq_58_49 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h31;
  wire          compressDataVec_hitReq_59_49 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h31;
  wire          compressDataVec_hitReq_60_49 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h31;
  wire          compressDataVec_hitReq_61_49 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h31;
  wire          compressDataVec_hitReq_62_49 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h31;
  wire          compressDataVec_hitReq_63_49 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h31;
  wire [7:0]    compressDataVec_selectReqData_49 =
    (compressDataVec_hitReq_0_49 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_49 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_49 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_49 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_49 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_49 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_49 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_49 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_49 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_49 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_49 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_49 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_49 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_49 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_49 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_49 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_49 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_49 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_49 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_49 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_49 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_49 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_49 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_49 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_49 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_49 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_49 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_49 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_49 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_49 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_49 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_49 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_49 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_49 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_49 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_49 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_49 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_49 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_49 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_49 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_49 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_49 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_49 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_49 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_49 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_49 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_49 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_49 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_49 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_49 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_49 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_49 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_49 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_49 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_49 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_49 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_49 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_49 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_49 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_49 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_49 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_49 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_49 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_49 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_49 = tailCount > 6'h31;
  wire          _GEN_1626 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h32;
  wire          compressDataVec_hitReq_0_50;
  assign compressDataVec_hitReq_0_50 = _GEN_1626;
  wire          compressDataVec_hitReq_0_178;
  assign compressDataVec_hitReq_0_178 = _GEN_1626;
  wire          _GEN_1627 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h32;
  wire          compressDataVec_hitReq_1_50;
  assign compressDataVec_hitReq_1_50 = _GEN_1627;
  wire          compressDataVec_hitReq_1_178;
  assign compressDataVec_hitReq_1_178 = _GEN_1627;
  wire          _GEN_1628 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h32;
  wire          compressDataVec_hitReq_2_50;
  assign compressDataVec_hitReq_2_50 = _GEN_1628;
  wire          compressDataVec_hitReq_2_178;
  assign compressDataVec_hitReq_2_178 = _GEN_1628;
  wire          _GEN_1629 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h32;
  wire          compressDataVec_hitReq_3_50;
  assign compressDataVec_hitReq_3_50 = _GEN_1629;
  wire          compressDataVec_hitReq_3_178;
  assign compressDataVec_hitReq_3_178 = _GEN_1629;
  wire          _GEN_1630 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h32;
  wire          compressDataVec_hitReq_4_50;
  assign compressDataVec_hitReq_4_50 = _GEN_1630;
  wire          compressDataVec_hitReq_4_178;
  assign compressDataVec_hitReq_4_178 = _GEN_1630;
  wire          _GEN_1631 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h32;
  wire          compressDataVec_hitReq_5_50;
  assign compressDataVec_hitReq_5_50 = _GEN_1631;
  wire          compressDataVec_hitReq_5_178;
  assign compressDataVec_hitReq_5_178 = _GEN_1631;
  wire          _GEN_1632 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h32;
  wire          compressDataVec_hitReq_6_50;
  assign compressDataVec_hitReq_6_50 = _GEN_1632;
  wire          compressDataVec_hitReq_6_178;
  assign compressDataVec_hitReq_6_178 = _GEN_1632;
  wire          _GEN_1633 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h32;
  wire          compressDataVec_hitReq_7_50;
  assign compressDataVec_hitReq_7_50 = _GEN_1633;
  wire          compressDataVec_hitReq_7_178;
  assign compressDataVec_hitReq_7_178 = _GEN_1633;
  wire          _GEN_1634 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h32;
  wire          compressDataVec_hitReq_8_50;
  assign compressDataVec_hitReq_8_50 = _GEN_1634;
  wire          compressDataVec_hitReq_8_178;
  assign compressDataVec_hitReq_8_178 = _GEN_1634;
  wire          _GEN_1635 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h32;
  wire          compressDataVec_hitReq_9_50;
  assign compressDataVec_hitReq_9_50 = _GEN_1635;
  wire          compressDataVec_hitReq_9_178;
  assign compressDataVec_hitReq_9_178 = _GEN_1635;
  wire          _GEN_1636 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h32;
  wire          compressDataVec_hitReq_10_50;
  assign compressDataVec_hitReq_10_50 = _GEN_1636;
  wire          compressDataVec_hitReq_10_178;
  assign compressDataVec_hitReq_10_178 = _GEN_1636;
  wire          _GEN_1637 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h32;
  wire          compressDataVec_hitReq_11_50;
  assign compressDataVec_hitReq_11_50 = _GEN_1637;
  wire          compressDataVec_hitReq_11_178;
  assign compressDataVec_hitReq_11_178 = _GEN_1637;
  wire          _GEN_1638 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h32;
  wire          compressDataVec_hitReq_12_50;
  assign compressDataVec_hitReq_12_50 = _GEN_1638;
  wire          compressDataVec_hitReq_12_178;
  assign compressDataVec_hitReq_12_178 = _GEN_1638;
  wire          _GEN_1639 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h32;
  wire          compressDataVec_hitReq_13_50;
  assign compressDataVec_hitReq_13_50 = _GEN_1639;
  wire          compressDataVec_hitReq_13_178;
  assign compressDataVec_hitReq_13_178 = _GEN_1639;
  wire          _GEN_1640 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h32;
  wire          compressDataVec_hitReq_14_50;
  assign compressDataVec_hitReq_14_50 = _GEN_1640;
  wire          compressDataVec_hitReq_14_178;
  assign compressDataVec_hitReq_14_178 = _GEN_1640;
  wire          _GEN_1641 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h32;
  wire          compressDataVec_hitReq_15_50;
  assign compressDataVec_hitReq_15_50 = _GEN_1641;
  wire          compressDataVec_hitReq_15_178;
  assign compressDataVec_hitReq_15_178 = _GEN_1641;
  wire          _GEN_1642 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h32;
  wire          compressDataVec_hitReq_16_50;
  assign compressDataVec_hitReq_16_50 = _GEN_1642;
  wire          compressDataVec_hitReq_16_178;
  assign compressDataVec_hitReq_16_178 = _GEN_1642;
  wire          _GEN_1643 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h32;
  wire          compressDataVec_hitReq_17_50;
  assign compressDataVec_hitReq_17_50 = _GEN_1643;
  wire          compressDataVec_hitReq_17_178;
  assign compressDataVec_hitReq_17_178 = _GEN_1643;
  wire          _GEN_1644 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h32;
  wire          compressDataVec_hitReq_18_50;
  assign compressDataVec_hitReq_18_50 = _GEN_1644;
  wire          compressDataVec_hitReq_18_178;
  assign compressDataVec_hitReq_18_178 = _GEN_1644;
  wire          _GEN_1645 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h32;
  wire          compressDataVec_hitReq_19_50;
  assign compressDataVec_hitReq_19_50 = _GEN_1645;
  wire          compressDataVec_hitReq_19_178;
  assign compressDataVec_hitReq_19_178 = _GEN_1645;
  wire          _GEN_1646 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h32;
  wire          compressDataVec_hitReq_20_50;
  assign compressDataVec_hitReq_20_50 = _GEN_1646;
  wire          compressDataVec_hitReq_20_178;
  assign compressDataVec_hitReq_20_178 = _GEN_1646;
  wire          _GEN_1647 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h32;
  wire          compressDataVec_hitReq_21_50;
  assign compressDataVec_hitReq_21_50 = _GEN_1647;
  wire          compressDataVec_hitReq_21_178;
  assign compressDataVec_hitReq_21_178 = _GEN_1647;
  wire          _GEN_1648 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h32;
  wire          compressDataVec_hitReq_22_50;
  assign compressDataVec_hitReq_22_50 = _GEN_1648;
  wire          compressDataVec_hitReq_22_178;
  assign compressDataVec_hitReq_22_178 = _GEN_1648;
  wire          _GEN_1649 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h32;
  wire          compressDataVec_hitReq_23_50;
  assign compressDataVec_hitReq_23_50 = _GEN_1649;
  wire          compressDataVec_hitReq_23_178;
  assign compressDataVec_hitReq_23_178 = _GEN_1649;
  wire          _GEN_1650 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h32;
  wire          compressDataVec_hitReq_24_50;
  assign compressDataVec_hitReq_24_50 = _GEN_1650;
  wire          compressDataVec_hitReq_24_178;
  assign compressDataVec_hitReq_24_178 = _GEN_1650;
  wire          _GEN_1651 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h32;
  wire          compressDataVec_hitReq_25_50;
  assign compressDataVec_hitReq_25_50 = _GEN_1651;
  wire          compressDataVec_hitReq_25_178;
  assign compressDataVec_hitReq_25_178 = _GEN_1651;
  wire          _GEN_1652 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h32;
  wire          compressDataVec_hitReq_26_50;
  assign compressDataVec_hitReq_26_50 = _GEN_1652;
  wire          compressDataVec_hitReq_26_178;
  assign compressDataVec_hitReq_26_178 = _GEN_1652;
  wire          _GEN_1653 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h32;
  wire          compressDataVec_hitReq_27_50;
  assign compressDataVec_hitReq_27_50 = _GEN_1653;
  wire          compressDataVec_hitReq_27_178;
  assign compressDataVec_hitReq_27_178 = _GEN_1653;
  wire          _GEN_1654 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h32;
  wire          compressDataVec_hitReq_28_50;
  assign compressDataVec_hitReq_28_50 = _GEN_1654;
  wire          compressDataVec_hitReq_28_178;
  assign compressDataVec_hitReq_28_178 = _GEN_1654;
  wire          _GEN_1655 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h32;
  wire          compressDataVec_hitReq_29_50;
  assign compressDataVec_hitReq_29_50 = _GEN_1655;
  wire          compressDataVec_hitReq_29_178;
  assign compressDataVec_hitReq_29_178 = _GEN_1655;
  wire          _GEN_1656 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h32;
  wire          compressDataVec_hitReq_30_50;
  assign compressDataVec_hitReq_30_50 = _GEN_1656;
  wire          compressDataVec_hitReq_30_178;
  assign compressDataVec_hitReq_30_178 = _GEN_1656;
  wire          _GEN_1657 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h32;
  wire          compressDataVec_hitReq_31_50;
  assign compressDataVec_hitReq_31_50 = _GEN_1657;
  wire          compressDataVec_hitReq_31_178;
  assign compressDataVec_hitReq_31_178 = _GEN_1657;
  wire          compressDataVec_hitReq_32_50 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h32;
  wire          compressDataVec_hitReq_33_50 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h32;
  wire          compressDataVec_hitReq_34_50 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h32;
  wire          compressDataVec_hitReq_35_50 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h32;
  wire          compressDataVec_hitReq_36_50 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h32;
  wire          compressDataVec_hitReq_37_50 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h32;
  wire          compressDataVec_hitReq_38_50 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h32;
  wire          compressDataVec_hitReq_39_50 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h32;
  wire          compressDataVec_hitReq_40_50 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h32;
  wire          compressDataVec_hitReq_41_50 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h32;
  wire          compressDataVec_hitReq_42_50 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h32;
  wire          compressDataVec_hitReq_43_50 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h32;
  wire          compressDataVec_hitReq_44_50 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h32;
  wire          compressDataVec_hitReq_45_50 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h32;
  wire          compressDataVec_hitReq_46_50 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h32;
  wire          compressDataVec_hitReq_47_50 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h32;
  wire          compressDataVec_hitReq_48_50 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h32;
  wire          compressDataVec_hitReq_49_50 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h32;
  wire          compressDataVec_hitReq_50_50 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h32;
  wire          compressDataVec_hitReq_51_50 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h32;
  wire          compressDataVec_hitReq_52_50 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h32;
  wire          compressDataVec_hitReq_53_50 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h32;
  wire          compressDataVec_hitReq_54_50 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h32;
  wire          compressDataVec_hitReq_55_50 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h32;
  wire          compressDataVec_hitReq_56_50 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h32;
  wire          compressDataVec_hitReq_57_50 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h32;
  wire          compressDataVec_hitReq_58_50 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h32;
  wire          compressDataVec_hitReq_59_50 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h32;
  wire          compressDataVec_hitReq_60_50 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h32;
  wire          compressDataVec_hitReq_61_50 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h32;
  wire          compressDataVec_hitReq_62_50 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h32;
  wire          compressDataVec_hitReq_63_50 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h32;
  wire [7:0]    compressDataVec_selectReqData_50 =
    (compressDataVec_hitReq_0_50 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_50 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_50 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_50 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_50 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_50 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_50 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_50 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_50 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_50 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_50 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_50 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_50 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_50 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_50 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_50 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_50 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_50 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_50 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_50 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_50 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_50 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_50 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_50 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_50 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_50 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_50 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_50 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_50 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_50 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_50 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_50 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_50 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_50 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_50 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_50 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_50 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_50 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_50 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_50 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_50 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_50 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_50 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_50 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_50 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_50 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_50 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_50 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_50 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_50 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_50 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_50 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_50 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_50 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_50 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_50 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_50 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_50 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_50 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_50 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_50 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_50 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_50 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_50 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_50 = tailCount > 6'h32;
  wire          _GEN_1658 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h33;
  wire          compressDataVec_hitReq_0_51;
  assign compressDataVec_hitReq_0_51 = _GEN_1658;
  wire          compressDataVec_hitReq_0_179;
  assign compressDataVec_hitReq_0_179 = _GEN_1658;
  wire          _GEN_1659 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h33;
  wire          compressDataVec_hitReq_1_51;
  assign compressDataVec_hitReq_1_51 = _GEN_1659;
  wire          compressDataVec_hitReq_1_179;
  assign compressDataVec_hitReq_1_179 = _GEN_1659;
  wire          _GEN_1660 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h33;
  wire          compressDataVec_hitReq_2_51;
  assign compressDataVec_hitReq_2_51 = _GEN_1660;
  wire          compressDataVec_hitReq_2_179;
  assign compressDataVec_hitReq_2_179 = _GEN_1660;
  wire          _GEN_1661 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h33;
  wire          compressDataVec_hitReq_3_51;
  assign compressDataVec_hitReq_3_51 = _GEN_1661;
  wire          compressDataVec_hitReq_3_179;
  assign compressDataVec_hitReq_3_179 = _GEN_1661;
  wire          _GEN_1662 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h33;
  wire          compressDataVec_hitReq_4_51;
  assign compressDataVec_hitReq_4_51 = _GEN_1662;
  wire          compressDataVec_hitReq_4_179;
  assign compressDataVec_hitReq_4_179 = _GEN_1662;
  wire          _GEN_1663 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h33;
  wire          compressDataVec_hitReq_5_51;
  assign compressDataVec_hitReq_5_51 = _GEN_1663;
  wire          compressDataVec_hitReq_5_179;
  assign compressDataVec_hitReq_5_179 = _GEN_1663;
  wire          _GEN_1664 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h33;
  wire          compressDataVec_hitReq_6_51;
  assign compressDataVec_hitReq_6_51 = _GEN_1664;
  wire          compressDataVec_hitReq_6_179;
  assign compressDataVec_hitReq_6_179 = _GEN_1664;
  wire          _GEN_1665 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h33;
  wire          compressDataVec_hitReq_7_51;
  assign compressDataVec_hitReq_7_51 = _GEN_1665;
  wire          compressDataVec_hitReq_7_179;
  assign compressDataVec_hitReq_7_179 = _GEN_1665;
  wire          _GEN_1666 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h33;
  wire          compressDataVec_hitReq_8_51;
  assign compressDataVec_hitReq_8_51 = _GEN_1666;
  wire          compressDataVec_hitReq_8_179;
  assign compressDataVec_hitReq_8_179 = _GEN_1666;
  wire          _GEN_1667 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h33;
  wire          compressDataVec_hitReq_9_51;
  assign compressDataVec_hitReq_9_51 = _GEN_1667;
  wire          compressDataVec_hitReq_9_179;
  assign compressDataVec_hitReq_9_179 = _GEN_1667;
  wire          _GEN_1668 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h33;
  wire          compressDataVec_hitReq_10_51;
  assign compressDataVec_hitReq_10_51 = _GEN_1668;
  wire          compressDataVec_hitReq_10_179;
  assign compressDataVec_hitReq_10_179 = _GEN_1668;
  wire          _GEN_1669 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h33;
  wire          compressDataVec_hitReq_11_51;
  assign compressDataVec_hitReq_11_51 = _GEN_1669;
  wire          compressDataVec_hitReq_11_179;
  assign compressDataVec_hitReq_11_179 = _GEN_1669;
  wire          _GEN_1670 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h33;
  wire          compressDataVec_hitReq_12_51;
  assign compressDataVec_hitReq_12_51 = _GEN_1670;
  wire          compressDataVec_hitReq_12_179;
  assign compressDataVec_hitReq_12_179 = _GEN_1670;
  wire          _GEN_1671 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h33;
  wire          compressDataVec_hitReq_13_51;
  assign compressDataVec_hitReq_13_51 = _GEN_1671;
  wire          compressDataVec_hitReq_13_179;
  assign compressDataVec_hitReq_13_179 = _GEN_1671;
  wire          _GEN_1672 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h33;
  wire          compressDataVec_hitReq_14_51;
  assign compressDataVec_hitReq_14_51 = _GEN_1672;
  wire          compressDataVec_hitReq_14_179;
  assign compressDataVec_hitReq_14_179 = _GEN_1672;
  wire          _GEN_1673 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h33;
  wire          compressDataVec_hitReq_15_51;
  assign compressDataVec_hitReq_15_51 = _GEN_1673;
  wire          compressDataVec_hitReq_15_179;
  assign compressDataVec_hitReq_15_179 = _GEN_1673;
  wire          _GEN_1674 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h33;
  wire          compressDataVec_hitReq_16_51;
  assign compressDataVec_hitReq_16_51 = _GEN_1674;
  wire          compressDataVec_hitReq_16_179;
  assign compressDataVec_hitReq_16_179 = _GEN_1674;
  wire          _GEN_1675 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h33;
  wire          compressDataVec_hitReq_17_51;
  assign compressDataVec_hitReq_17_51 = _GEN_1675;
  wire          compressDataVec_hitReq_17_179;
  assign compressDataVec_hitReq_17_179 = _GEN_1675;
  wire          _GEN_1676 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h33;
  wire          compressDataVec_hitReq_18_51;
  assign compressDataVec_hitReq_18_51 = _GEN_1676;
  wire          compressDataVec_hitReq_18_179;
  assign compressDataVec_hitReq_18_179 = _GEN_1676;
  wire          _GEN_1677 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h33;
  wire          compressDataVec_hitReq_19_51;
  assign compressDataVec_hitReq_19_51 = _GEN_1677;
  wire          compressDataVec_hitReq_19_179;
  assign compressDataVec_hitReq_19_179 = _GEN_1677;
  wire          _GEN_1678 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h33;
  wire          compressDataVec_hitReq_20_51;
  assign compressDataVec_hitReq_20_51 = _GEN_1678;
  wire          compressDataVec_hitReq_20_179;
  assign compressDataVec_hitReq_20_179 = _GEN_1678;
  wire          _GEN_1679 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h33;
  wire          compressDataVec_hitReq_21_51;
  assign compressDataVec_hitReq_21_51 = _GEN_1679;
  wire          compressDataVec_hitReq_21_179;
  assign compressDataVec_hitReq_21_179 = _GEN_1679;
  wire          _GEN_1680 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h33;
  wire          compressDataVec_hitReq_22_51;
  assign compressDataVec_hitReq_22_51 = _GEN_1680;
  wire          compressDataVec_hitReq_22_179;
  assign compressDataVec_hitReq_22_179 = _GEN_1680;
  wire          _GEN_1681 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h33;
  wire          compressDataVec_hitReq_23_51;
  assign compressDataVec_hitReq_23_51 = _GEN_1681;
  wire          compressDataVec_hitReq_23_179;
  assign compressDataVec_hitReq_23_179 = _GEN_1681;
  wire          _GEN_1682 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h33;
  wire          compressDataVec_hitReq_24_51;
  assign compressDataVec_hitReq_24_51 = _GEN_1682;
  wire          compressDataVec_hitReq_24_179;
  assign compressDataVec_hitReq_24_179 = _GEN_1682;
  wire          _GEN_1683 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h33;
  wire          compressDataVec_hitReq_25_51;
  assign compressDataVec_hitReq_25_51 = _GEN_1683;
  wire          compressDataVec_hitReq_25_179;
  assign compressDataVec_hitReq_25_179 = _GEN_1683;
  wire          _GEN_1684 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h33;
  wire          compressDataVec_hitReq_26_51;
  assign compressDataVec_hitReq_26_51 = _GEN_1684;
  wire          compressDataVec_hitReq_26_179;
  assign compressDataVec_hitReq_26_179 = _GEN_1684;
  wire          _GEN_1685 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h33;
  wire          compressDataVec_hitReq_27_51;
  assign compressDataVec_hitReq_27_51 = _GEN_1685;
  wire          compressDataVec_hitReq_27_179;
  assign compressDataVec_hitReq_27_179 = _GEN_1685;
  wire          _GEN_1686 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h33;
  wire          compressDataVec_hitReq_28_51;
  assign compressDataVec_hitReq_28_51 = _GEN_1686;
  wire          compressDataVec_hitReq_28_179;
  assign compressDataVec_hitReq_28_179 = _GEN_1686;
  wire          _GEN_1687 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h33;
  wire          compressDataVec_hitReq_29_51;
  assign compressDataVec_hitReq_29_51 = _GEN_1687;
  wire          compressDataVec_hitReq_29_179;
  assign compressDataVec_hitReq_29_179 = _GEN_1687;
  wire          _GEN_1688 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h33;
  wire          compressDataVec_hitReq_30_51;
  assign compressDataVec_hitReq_30_51 = _GEN_1688;
  wire          compressDataVec_hitReq_30_179;
  assign compressDataVec_hitReq_30_179 = _GEN_1688;
  wire          _GEN_1689 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h33;
  wire          compressDataVec_hitReq_31_51;
  assign compressDataVec_hitReq_31_51 = _GEN_1689;
  wire          compressDataVec_hitReq_31_179;
  assign compressDataVec_hitReq_31_179 = _GEN_1689;
  wire          compressDataVec_hitReq_32_51 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h33;
  wire          compressDataVec_hitReq_33_51 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h33;
  wire          compressDataVec_hitReq_34_51 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h33;
  wire          compressDataVec_hitReq_35_51 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h33;
  wire          compressDataVec_hitReq_36_51 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h33;
  wire          compressDataVec_hitReq_37_51 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h33;
  wire          compressDataVec_hitReq_38_51 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h33;
  wire          compressDataVec_hitReq_39_51 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h33;
  wire          compressDataVec_hitReq_40_51 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h33;
  wire          compressDataVec_hitReq_41_51 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h33;
  wire          compressDataVec_hitReq_42_51 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h33;
  wire          compressDataVec_hitReq_43_51 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h33;
  wire          compressDataVec_hitReq_44_51 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h33;
  wire          compressDataVec_hitReq_45_51 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h33;
  wire          compressDataVec_hitReq_46_51 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h33;
  wire          compressDataVec_hitReq_47_51 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h33;
  wire          compressDataVec_hitReq_48_51 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h33;
  wire          compressDataVec_hitReq_49_51 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h33;
  wire          compressDataVec_hitReq_50_51 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h33;
  wire          compressDataVec_hitReq_51_51 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h33;
  wire          compressDataVec_hitReq_52_51 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h33;
  wire          compressDataVec_hitReq_53_51 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h33;
  wire          compressDataVec_hitReq_54_51 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h33;
  wire          compressDataVec_hitReq_55_51 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h33;
  wire          compressDataVec_hitReq_56_51 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h33;
  wire          compressDataVec_hitReq_57_51 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h33;
  wire          compressDataVec_hitReq_58_51 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h33;
  wire          compressDataVec_hitReq_59_51 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h33;
  wire          compressDataVec_hitReq_60_51 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h33;
  wire          compressDataVec_hitReq_61_51 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h33;
  wire          compressDataVec_hitReq_62_51 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h33;
  wire          compressDataVec_hitReq_63_51 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h33;
  wire [7:0]    compressDataVec_selectReqData_51 =
    (compressDataVec_hitReq_0_51 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_51 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_51 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_51 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_51 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_51 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_51 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_51 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_51 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_51 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_51 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_51 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_51 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_51 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_51 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_51 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_51 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_51 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_51 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_51 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_51 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_51 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_51 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_51 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_51 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_51 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_51 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_51 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_51 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_51 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_51 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_51 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_51 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_51 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_51 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_51 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_51 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_51 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_51 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_51 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_51 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_51 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_51 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_51 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_51 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_51 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_51 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_51 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_51 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_51 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_51 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_51 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_51 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_51 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_51 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_51 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_51 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_51 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_51 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_51 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_51 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_51 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_51 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_51 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_51 = tailCount > 6'h33;
  wire          _GEN_1690 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h34;
  wire          compressDataVec_hitReq_0_52;
  assign compressDataVec_hitReq_0_52 = _GEN_1690;
  wire          compressDataVec_hitReq_0_180;
  assign compressDataVec_hitReq_0_180 = _GEN_1690;
  wire          _GEN_1691 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h34;
  wire          compressDataVec_hitReq_1_52;
  assign compressDataVec_hitReq_1_52 = _GEN_1691;
  wire          compressDataVec_hitReq_1_180;
  assign compressDataVec_hitReq_1_180 = _GEN_1691;
  wire          _GEN_1692 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h34;
  wire          compressDataVec_hitReq_2_52;
  assign compressDataVec_hitReq_2_52 = _GEN_1692;
  wire          compressDataVec_hitReq_2_180;
  assign compressDataVec_hitReq_2_180 = _GEN_1692;
  wire          _GEN_1693 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h34;
  wire          compressDataVec_hitReq_3_52;
  assign compressDataVec_hitReq_3_52 = _GEN_1693;
  wire          compressDataVec_hitReq_3_180;
  assign compressDataVec_hitReq_3_180 = _GEN_1693;
  wire          _GEN_1694 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h34;
  wire          compressDataVec_hitReq_4_52;
  assign compressDataVec_hitReq_4_52 = _GEN_1694;
  wire          compressDataVec_hitReq_4_180;
  assign compressDataVec_hitReq_4_180 = _GEN_1694;
  wire          _GEN_1695 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h34;
  wire          compressDataVec_hitReq_5_52;
  assign compressDataVec_hitReq_5_52 = _GEN_1695;
  wire          compressDataVec_hitReq_5_180;
  assign compressDataVec_hitReq_5_180 = _GEN_1695;
  wire          _GEN_1696 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h34;
  wire          compressDataVec_hitReq_6_52;
  assign compressDataVec_hitReq_6_52 = _GEN_1696;
  wire          compressDataVec_hitReq_6_180;
  assign compressDataVec_hitReq_6_180 = _GEN_1696;
  wire          _GEN_1697 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h34;
  wire          compressDataVec_hitReq_7_52;
  assign compressDataVec_hitReq_7_52 = _GEN_1697;
  wire          compressDataVec_hitReq_7_180;
  assign compressDataVec_hitReq_7_180 = _GEN_1697;
  wire          _GEN_1698 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h34;
  wire          compressDataVec_hitReq_8_52;
  assign compressDataVec_hitReq_8_52 = _GEN_1698;
  wire          compressDataVec_hitReq_8_180;
  assign compressDataVec_hitReq_8_180 = _GEN_1698;
  wire          _GEN_1699 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h34;
  wire          compressDataVec_hitReq_9_52;
  assign compressDataVec_hitReq_9_52 = _GEN_1699;
  wire          compressDataVec_hitReq_9_180;
  assign compressDataVec_hitReq_9_180 = _GEN_1699;
  wire          _GEN_1700 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h34;
  wire          compressDataVec_hitReq_10_52;
  assign compressDataVec_hitReq_10_52 = _GEN_1700;
  wire          compressDataVec_hitReq_10_180;
  assign compressDataVec_hitReq_10_180 = _GEN_1700;
  wire          _GEN_1701 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h34;
  wire          compressDataVec_hitReq_11_52;
  assign compressDataVec_hitReq_11_52 = _GEN_1701;
  wire          compressDataVec_hitReq_11_180;
  assign compressDataVec_hitReq_11_180 = _GEN_1701;
  wire          _GEN_1702 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h34;
  wire          compressDataVec_hitReq_12_52;
  assign compressDataVec_hitReq_12_52 = _GEN_1702;
  wire          compressDataVec_hitReq_12_180;
  assign compressDataVec_hitReq_12_180 = _GEN_1702;
  wire          _GEN_1703 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h34;
  wire          compressDataVec_hitReq_13_52;
  assign compressDataVec_hitReq_13_52 = _GEN_1703;
  wire          compressDataVec_hitReq_13_180;
  assign compressDataVec_hitReq_13_180 = _GEN_1703;
  wire          _GEN_1704 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h34;
  wire          compressDataVec_hitReq_14_52;
  assign compressDataVec_hitReq_14_52 = _GEN_1704;
  wire          compressDataVec_hitReq_14_180;
  assign compressDataVec_hitReq_14_180 = _GEN_1704;
  wire          _GEN_1705 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h34;
  wire          compressDataVec_hitReq_15_52;
  assign compressDataVec_hitReq_15_52 = _GEN_1705;
  wire          compressDataVec_hitReq_15_180;
  assign compressDataVec_hitReq_15_180 = _GEN_1705;
  wire          _GEN_1706 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h34;
  wire          compressDataVec_hitReq_16_52;
  assign compressDataVec_hitReq_16_52 = _GEN_1706;
  wire          compressDataVec_hitReq_16_180;
  assign compressDataVec_hitReq_16_180 = _GEN_1706;
  wire          _GEN_1707 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h34;
  wire          compressDataVec_hitReq_17_52;
  assign compressDataVec_hitReq_17_52 = _GEN_1707;
  wire          compressDataVec_hitReq_17_180;
  assign compressDataVec_hitReq_17_180 = _GEN_1707;
  wire          _GEN_1708 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h34;
  wire          compressDataVec_hitReq_18_52;
  assign compressDataVec_hitReq_18_52 = _GEN_1708;
  wire          compressDataVec_hitReq_18_180;
  assign compressDataVec_hitReq_18_180 = _GEN_1708;
  wire          _GEN_1709 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h34;
  wire          compressDataVec_hitReq_19_52;
  assign compressDataVec_hitReq_19_52 = _GEN_1709;
  wire          compressDataVec_hitReq_19_180;
  assign compressDataVec_hitReq_19_180 = _GEN_1709;
  wire          _GEN_1710 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h34;
  wire          compressDataVec_hitReq_20_52;
  assign compressDataVec_hitReq_20_52 = _GEN_1710;
  wire          compressDataVec_hitReq_20_180;
  assign compressDataVec_hitReq_20_180 = _GEN_1710;
  wire          _GEN_1711 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h34;
  wire          compressDataVec_hitReq_21_52;
  assign compressDataVec_hitReq_21_52 = _GEN_1711;
  wire          compressDataVec_hitReq_21_180;
  assign compressDataVec_hitReq_21_180 = _GEN_1711;
  wire          _GEN_1712 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h34;
  wire          compressDataVec_hitReq_22_52;
  assign compressDataVec_hitReq_22_52 = _GEN_1712;
  wire          compressDataVec_hitReq_22_180;
  assign compressDataVec_hitReq_22_180 = _GEN_1712;
  wire          _GEN_1713 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h34;
  wire          compressDataVec_hitReq_23_52;
  assign compressDataVec_hitReq_23_52 = _GEN_1713;
  wire          compressDataVec_hitReq_23_180;
  assign compressDataVec_hitReq_23_180 = _GEN_1713;
  wire          _GEN_1714 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h34;
  wire          compressDataVec_hitReq_24_52;
  assign compressDataVec_hitReq_24_52 = _GEN_1714;
  wire          compressDataVec_hitReq_24_180;
  assign compressDataVec_hitReq_24_180 = _GEN_1714;
  wire          _GEN_1715 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h34;
  wire          compressDataVec_hitReq_25_52;
  assign compressDataVec_hitReq_25_52 = _GEN_1715;
  wire          compressDataVec_hitReq_25_180;
  assign compressDataVec_hitReq_25_180 = _GEN_1715;
  wire          _GEN_1716 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h34;
  wire          compressDataVec_hitReq_26_52;
  assign compressDataVec_hitReq_26_52 = _GEN_1716;
  wire          compressDataVec_hitReq_26_180;
  assign compressDataVec_hitReq_26_180 = _GEN_1716;
  wire          _GEN_1717 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h34;
  wire          compressDataVec_hitReq_27_52;
  assign compressDataVec_hitReq_27_52 = _GEN_1717;
  wire          compressDataVec_hitReq_27_180;
  assign compressDataVec_hitReq_27_180 = _GEN_1717;
  wire          _GEN_1718 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h34;
  wire          compressDataVec_hitReq_28_52;
  assign compressDataVec_hitReq_28_52 = _GEN_1718;
  wire          compressDataVec_hitReq_28_180;
  assign compressDataVec_hitReq_28_180 = _GEN_1718;
  wire          _GEN_1719 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h34;
  wire          compressDataVec_hitReq_29_52;
  assign compressDataVec_hitReq_29_52 = _GEN_1719;
  wire          compressDataVec_hitReq_29_180;
  assign compressDataVec_hitReq_29_180 = _GEN_1719;
  wire          _GEN_1720 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h34;
  wire          compressDataVec_hitReq_30_52;
  assign compressDataVec_hitReq_30_52 = _GEN_1720;
  wire          compressDataVec_hitReq_30_180;
  assign compressDataVec_hitReq_30_180 = _GEN_1720;
  wire          _GEN_1721 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h34;
  wire          compressDataVec_hitReq_31_52;
  assign compressDataVec_hitReq_31_52 = _GEN_1721;
  wire          compressDataVec_hitReq_31_180;
  assign compressDataVec_hitReq_31_180 = _GEN_1721;
  wire          compressDataVec_hitReq_32_52 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h34;
  wire          compressDataVec_hitReq_33_52 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h34;
  wire          compressDataVec_hitReq_34_52 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h34;
  wire          compressDataVec_hitReq_35_52 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h34;
  wire          compressDataVec_hitReq_36_52 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h34;
  wire          compressDataVec_hitReq_37_52 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h34;
  wire          compressDataVec_hitReq_38_52 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h34;
  wire          compressDataVec_hitReq_39_52 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h34;
  wire          compressDataVec_hitReq_40_52 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h34;
  wire          compressDataVec_hitReq_41_52 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h34;
  wire          compressDataVec_hitReq_42_52 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h34;
  wire          compressDataVec_hitReq_43_52 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h34;
  wire          compressDataVec_hitReq_44_52 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h34;
  wire          compressDataVec_hitReq_45_52 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h34;
  wire          compressDataVec_hitReq_46_52 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h34;
  wire          compressDataVec_hitReq_47_52 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h34;
  wire          compressDataVec_hitReq_48_52 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h34;
  wire          compressDataVec_hitReq_49_52 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h34;
  wire          compressDataVec_hitReq_50_52 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h34;
  wire          compressDataVec_hitReq_51_52 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h34;
  wire          compressDataVec_hitReq_52_52 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h34;
  wire          compressDataVec_hitReq_53_52 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h34;
  wire          compressDataVec_hitReq_54_52 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h34;
  wire          compressDataVec_hitReq_55_52 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h34;
  wire          compressDataVec_hitReq_56_52 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h34;
  wire          compressDataVec_hitReq_57_52 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h34;
  wire          compressDataVec_hitReq_58_52 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h34;
  wire          compressDataVec_hitReq_59_52 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h34;
  wire          compressDataVec_hitReq_60_52 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h34;
  wire          compressDataVec_hitReq_61_52 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h34;
  wire          compressDataVec_hitReq_62_52 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h34;
  wire          compressDataVec_hitReq_63_52 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h34;
  wire [7:0]    compressDataVec_selectReqData_52 =
    (compressDataVec_hitReq_0_52 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_52 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_52 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_52 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_52 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_52 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_52 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_52 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_52 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_52 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_52 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_52 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_52 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_52 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_52 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_52 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_52 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_52 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_52 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_52 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_52 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_52 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_52 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_52 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_52 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_52 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_52 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_52 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_52 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_52 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_52 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_52 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_52 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_52 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_52 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_52 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_52 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_52 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_52 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_52 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_52 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_52 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_52 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_52 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_52 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_52 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_52 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_52 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_52 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_52 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_52 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_52 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_52 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_52 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_52 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_52 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_52 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_52 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_52 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_52 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_52 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_52 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_52 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_52 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_52 = tailCount > 6'h34;
  wire          _GEN_1722 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h35;
  wire          compressDataVec_hitReq_0_53;
  assign compressDataVec_hitReq_0_53 = _GEN_1722;
  wire          compressDataVec_hitReq_0_181;
  assign compressDataVec_hitReq_0_181 = _GEN_1722;
  wire          _GEN_1723 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h35;
  wire          compressDataVec_hitReq_1_53;
  assign compressDataVec_hitReq_1_53 = _GEN_1723;
  wire          compressDataVec_hitReq_1_181;
  assign compressDataVec_hitReq_1_181 = _GEN_1723;
  wire          _GEN_1724 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h35;
  wire          compressDataVec_hitReq_2_53;
  assign compressDataVec_hitReq_2_53 = _GEN_1724;
  wire          compressDataVec_hitReq_2_181;
  assign compressDataVec_hitReq_2_181 = _GEN_1724;
  wire          _GEN_1725 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h35;
  wire          compressDataVec_hitReq_3_53;
  assign compressDataVec_hitReq_3_53 = _GEN_1725;
  wire          compressDataVec_hitReq_3_181;
  assign compressDataVec_hitReq_3_181 = _GEN_1725;
  wire          _GEN_1726 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h35;
  wire          compressDataVec_hitReq_4_53;
  assign compressDataVec_hitReq_4_53 = _GEN_1726;
  wire          compressDataVec_hitReq_4_181;
  assign compressDataVec_hitReq_4_181 = _GEN_1726;
  wire          _GEN_1727 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h35;
  wire          compressDataVec_hitReq_5_53;
  assign compressDataVec_hitReq_5_53 = _GEN_1727;
  wire          compressDataVec_hitReq_5_181;
  assign compressDataVec_hitReq_5_181 = _GEN_1727;
  wire          _GEN_1728 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h35;
  wire          compressDataVec_hitReq_6_53;
  assign compressDataVec_hitReq_6_53 = _GEN_1728;
  wire          compressDataVec_hitReq_6_181;
  assign compressDataVec_hitReq_6_181 = _GEN_1728;
  wire          _GEN_1729 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h35;
  wire          compressDataVec_hitReq_7_53;
  assign compressDataVec_hitReq_7_53 = _GEN_1729;
  wire          compressDataVec_hitReq_7_181;
  assign compressDataVec_hitReq_7_181 = _GEN_1729;
  wire          _GEN_1730 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h35;
  wire          compressDataVec_hitReq_8_53;
  assign compressDataVec_hitReq_8_53 = _GEN_1730;
  wire          compressDataVec_hitReq_8_181;
  assign compressDataVec_hitReq_8_181 = _GEN_1730;
  wire          _GEN_1731 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h35;
  wire          compressDataVec_hitReq_9_53;
  assign compressDataVec_hitReq_9_53 = _GEN_1731;
  wire          compressDataVec_hitReq_9_181;
  assign compressDataVec_hitReq_9_181 = _GEN_1731;
  wire          _GEN_1732 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h35;
  wire          compressDataVec_hitReq_10_53;
  assign compressDataVec_hitReq_10_53 = _GEN_1732;
  wire          compressDataVec_hitReq_10_181;
  assign compressDataVec_hitReq_10_181 = _GEN_1732;
  wire          _GEN_1733 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h35;
  wire          compressDataVec_hitReq_11_53;
  assign compressDataVec_hitReq_11_53 = _GEN_1733;
  wire          compressDataVec_hitReq_11_181;
  assign compressDataVec_hitReq_11_181 = _GEN_1733;
  wire          _GEN_1734 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h35;
  wire          compressDataVec_hitReq_12_53;
  assign compressDataVec_hitReq_12_53 = _GEN_1734;
  wire          compressDataVec_hitReq_12_181;
  assign compressDataVec_hitReq_12_181 = _GEN_1734;
  wire          _GEN_1735 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h35;
  wire          compressDataVec_hitReq_13_53;
  assign compressDataVec_hitReq_13_53 = _GEN_1735;
  wire          compressDataVec_hitReq_13_181;
  assign compressDataVec_hitReq_13_181 = _GEN_1735;
  wire          _GEN_1736 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h35;
  wire          compressDataVec_hitReq_14_53;
  assign compressDataVec_hitReq_14_53 = _GEN_1736;
  wire          compressDataVec_hitReq_14_181;
  assign compressDataVec_hitReq_14_181 = _GEN_1736;
  wire          _GEN_1737 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h35;
  wire          compressDataVec_hitReq_15_53;
  assign compressDataVec_hitReq_15_53 = _GEN_1737;
  wire          compressDataVec_hitReq_15_181;
  assign compressDataVec_hitReq_15_181 = _GEN_1737;
  wire          _GEN_1738 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h35;
  wire          compressDataVec_hitReq_16_53;
  assign compressDataVec_hitReq_16_53 = _GEN_1738;
  wire          compressDataVec_hitReq_16_181;
  assign compressDataVec_hitReq_16_181 = _GEN_1738;
  wire          _GEN_1739 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h35;
  wire          compressDataVec_hitReq_17_53;
  assign compressDataVec_hitReq_17_53 = _GEN_1739;
  wire          compressDataVec_hitReq_17_181;
  assign compressDataVec_hitReq_17_181 = _GEN_1739;
  wire          _GEN_1740 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h35;
  wire          compressDataVec_hitReq_18_53;
  assign compressDataVec_hitReq_18_53 = _GEN_1740;
  wire          compressDataVec_hitReq_18_181;
  assign compressDataVec_hitReq_18_181 = _GEN_1740;
  wire          _GEN_1741 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h35;
  wire          compressDataVec_hitReq_19_53;
  assign compressDataVec_hitReq_19_53 = _GEN_1741;
  wire          compressDataVec_hitReq_19_181;
  assign compressDataVec_hitReq_19_181 = _GEN_1741;
  wire          _GEN_1742 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h35;
  wire          compressDataVec_hitReq_20_53;
  assign compressDataVec_hitReq_20_53 = _GEN_1742;
  wire          compressDataVec_hitReq_20_181;
  assign compressDataVec_hitReq_20_181 = _GEN_1742;
  wire          _GEN_1743 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h35;
  wire          compressDataVec_hitReq_21_53;
  assign compressDataVec_hitReq_21_53 = _GEN_1743;
  wire          compressDataVec_hitReq_21_181;
  assign compressDataVec_hitReq_21_181 = _GEN_1743;
  wire          _GEN_1744 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h35;
  wire          compressDataVec_hitReq_22_53;
  assign compressDataVec_hitReq_22_53 = _GEN_1744;
  wire          compressDataVec_hitReq_22_181;
  assign compressDataVec_hitReq_22_181 = _GEN_1744;
  wire          _GEN_1745 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h35;
  wire          compressDataVec_hitReq_23_53;
  assign compressDataVec_hitReq_23_53 = _GEN_1745;
  wire          compressDataVec_hitReq_23_181;
  assign compressDataVec_hitReq_23_181 = _GEN_1745;
  wire          _GEN_1746 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h35;
  wire          compressDataVec_hitReq_24_53;
  assign compressDataVec_hitReq_24_53 = _GEN_1746;
  wire          compressDataVec_hitReq_24_181;
  assign compressDataVec_hitReq_24_181 = _GEN_1746;
  wire          _GEN_1747 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h35;
  wire          compressDataVec_hitReq_25_53;
  assign compressDataVec_hitReq_25_53 = _GEN_1747;
  wire          compressDataVec_hitReq_25_181;
  assign compressDataVec_hitReq_25_181 = _GEN_1747;
  wire          _GEN_1748 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h35;
  wire          compressDataVec_hitReq_26_53;
  assign compressDataVec_hitReq_26_53 = _GEN_1748;
  wire          compressDataVec_hitReq_26_181;
  assign compressDataVec_hitReq_26_181 = _GEN_1748;
  wire          _GEN_1749 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h35;
  wire          compressDataVec_hitReq_27_53;
  assign compressDataVec_hitReq_27_53 = _GEN_1749;
  wire          compressDataVec_hitReq_27_181;
  assign compressDataVec_hitReq_27_181 = _GEN_1749;
  wire          _GEN_1750 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h35;
  wire          compressDataVec_hitReq_28_53;
  assign compressDataVec_hitReq_28_53 = _GEN_1750;
  wire          compressDataVec_hitReq_28_181;
  assign compressDataVec_hitReq_28_181 = _GEN_1750;
  wire          _GEN_1751 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h35;
  wire          compressDataVec_hitReq_29_53;
  assign compressDataVec_hitReq_29_53 = _GEN_1751;
  wire          compressDataVec_hitReq_29_181;
  assign compressDataVec_hitReq_29_181 = _GEN_1751;
  wire          _GEN_1752 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h35;
  wire          compressDataVec_hitReq_30_53;
  assign compressDataVec_hitReq_30_53 = _GEN_1752;
  wire          compressDataVec_hitReq_30_181;
  assign compressDataVec_hitReq_30_181 = _GEN_1752;
  wire          _GEN_1753 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h35;
  wire          compressDataVec_hitReq_31_53;
  assign compressDataVec_hitReq_31_53 = _GEN_1753;
  wire          compressDataVec_hitReq_31_181;
  assign compressDataVec_hitReq_31_181 = _GEN_1753;
  wire          compressDataVec_hitReq_32_53 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h35;
  wire          compressDataVec_hitReq_33_53 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h35;
  wire          compressDataVec_hitReq_34_53 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h35;
  wire          compressDataVec_hitReq_35_53 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h35;
  wire          compressDataVec_hitReq_36_53 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h35;
  wire          compressDataVec_hitReq_37_53 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h35;
  wire          compressDataVec_hitReq_38_53 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h35;
  wire          compressDataVec_hitReq_39_53 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h35;
  wire          compressDataVec_hitReq_40_53 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h35;
  wire          compressDataVec_hitReq_41_53 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h35;
  wire          compressDataVec_hitReq_42_53 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h35;
  wire          compressDataVec_hitReq_43_53 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h35;
  wire          compressDataVec_hitReq_44_53 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h35;
  wire          compressDataVec_hitReq_45_53 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h35;
  wire          compressDataVec_hitReq_46_53 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h35;
  wire          compressDataVec_hitReq_47_53 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h35;
  wire          compressDataVec_hitReq_48_53 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h35;
  wire          compressDataVec_hitReq_49_53 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h35;
  wire          compressDataVec_hitReq_50_53 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h35;
  wire          compressDataVec_hitReq_51_53 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h35;
  wire          compressDataVec_hitReq_52_53 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h35;
  wire          compressDataVec_hitReq_53_53 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h35;
  wire          compressDataVec_hitReq_54_53 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h35;
  wire          compressDataVec_hitReq_55_53 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h35;
  wire          compressDataVec_hitReq_56_53 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h35;
  wire          compressDataVec_hitReq_57_53 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h35;
  wire          compressDataVec_hitReq_58_53 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h35;
  wire          compressDataVec_hitReq_59_53 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h35;
  wire          compressDataVec_hitReq_60_53 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h35;
  wire          compressDataVec_hitReq_61_53 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h35;
  wire          compressDataVec_hitReq_62_53 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h35;
  wire          compressDataVec_hitReq_63_53 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h35;
  wire [7:0]    compressDataVec_selectReqData_53 =
    (compressDataVec_hitReq_0_53 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_53 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_53 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_53 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_53 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_53 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_53 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_53 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_53 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_53 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_53 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_53 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_53 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_53 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_53 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_53 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_53 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_53 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_53 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_53 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_53 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_53 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_53 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_53 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_53 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_53 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_53 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_53 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_53 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_53 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_53 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_53 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_53 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_53 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_53 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_53 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_53 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_53 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_53 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_53 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_53 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_53 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_53 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_53 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_53 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_53 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_53 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_53 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_53 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_53 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_53 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_53 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_53 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_53 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_53 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_53 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_53 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_53 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_53 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_53 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_53 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_53 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_53 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_53 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_53 = tailCount > 6'h35;
  wire          _GEN_1754 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h36;
  wire          compressDataVec_hitReq_0_54;
  assign compressDataVec_hitReq_0_54 = _GEN_1754;
  wire          compressDataVec_hitReq_0_182;
  assign compressDataVec_hitReq_0_182 = _GEN_1754;
  wire          _GEN_1755 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h36;
  wire          compressDataVec_hitReq_1_54;
  assign compressDataVec_hitReq_1_54 = _GEN_1755;
  wire          compressDataVec_hitReq_1_182;
  assign compressDataVec_hitReq_1_182 = _GEN_1755;
  wire          _GEN_1756 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h36;
  wire          compressDataVec_hitReq_2_54;
  assign compressDataVec_hitReq_2_54 = _GEN_1756;
  wire          compressDataVec_hitReq_2_182;
  assign compressDataVec_hitReq_2_182 = _GEN_1756;
  wire          _GEN_1757 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h36;
  wire          compressDataVec_hitReq_3_54;
  assign compressDataVec_hitReq_3_54 = _GEN_1757;
  wire          compressDataVec_hitReq_3_182;
  assign compressDataVec_hitReq_3_182 = _GEN_1757;
  wire          _GEN_1758 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h36;
  wire          compressDataVec_hitReq_4_54;
  assign compressDataVec_hitReq_4_54 = _GEN_1758;
  wire          compressDataVec_hitReq_4_182;
  assign compressDataVec_hitReq_4_182 = _GEN_1758;
  wire          _GEN_1759 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h36;
  wire          compressDataVec_hitReq_5_54;
  assign compressDataVec_hitReq_5_54 = _GEN_1759;
  wire          compressDataVec_hitReq_5_182;
  assign compressDataVec_hitReq_5_182 = _GEN_1759;
  wire          _GEN_1760 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h36;
  wire          compressDataVec_hitReq_6_54;
  assign compressDataVec_hitReq_6_54 = _GEN_1760;
  wire          compressDataVec_hitReq_6_182;
  assign compressDataVec_hitReq_6_182 = _GEN_1760;
  wire          _GEN_1761 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h36;
  wire          compressDataVec_hitReq_7_54;
  assign compressDataVec_hitReq_7_54 = _GEN_1761;
  wire          compressDataVec_hitReq_7_182;
  assign compressDataVec_hitReq_7_182 = _GEN_1761;
  wire          _GEN_1762 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h36;
  wire          compressDataVec_hitReq_8_54;
  assign compressDataVec_hitReq_8_54 = _GEN_1762;
  wire          compressDataVec_hitReq_8_182;
  assign compressDataVec_hitReq_8_182 = _GEN_1762;
  wire          _GEN_1763 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h36;
  wire          compressDataVec_hitReq_9_54;
  assign compressDataVec_hitReq_9_54 = _GEN_1763;
  wire          compressDataVec_hitReq_9_182;
  assign compressDataVec_hitReq_9_182 = _GEN_1763;
  wire          _GEN_1764 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h36;
  wire          compressDataVec_hitReq_10_54;
  assign compressDataVec_hitReq_10_54 = _GEN_1764;
  wire          compressDataVec_hitReq_10_182;
  assign compressDataVec_hitReq_10_182 = _GEN_1764;
  wire          _GEN_1765 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h36;
  wire          compressDataVec_hitReq_11_54;
  assign compressDataVec_hitReq_11_54 = _GEN_1765;
  wire          compressDataVec_hitReq_11_182;
  assign compressDataVec_hitReq_11_182 = _GEN_1765;
  wire          _GEN_1766 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h36;
  wire          compressDataVec_hitReq_12_54;
  assign compressDataVec_hitReq_12_54 = _GEN_1766;
  wire          compressDataVec_hitReq_12_182;
  assign compressDataVec_hitReq_12_182 = _GEN_1766;
  wire          _GEN_1767 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h36;
  wire          compressDataVec_hitReq_13_54;
  assign compressDataVec_hitReq_13_54 = _GEN_1767;
  wire          compressDataVec_hitReq_13_182;
  assign compressDataVec_hitReq_13_182 = _GEN_1767;
  wire          _GEN_1768 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h36;
  wire          compressDataVec_hitReq_14_54;
  assign compressDataVec_hitReq_14_54 = _GEN_1768;
  wire          compressDataVec_hitReq_14_182;
  assign compressDataVec_hitReq_14_182 = _GEN_1768;
  wire          _GEN_1769 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h36;
  wire          compressDataVec_hitReq_15_54;
  assign compressDataVec_hitReq_15_54 = _GEN_1769;
  wire          compressDataVec_hitReq_15_182;
  assign compressDataVec_hitReq_15_182 = _GEN_1769;
  wire          _GEN_1770 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h36;
  wire          compressDataVec_hitReq_16_54;
  assign compressDataVec_hitReq_16_54 = _GEN_1770;
  wire          compressDataVec_hitReq_16_182;
  assign compressDataVec_hitReq_16_182 = _GEN_1770;
  wire          _GEN_1771 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h36;
  wire          compressDataVec_hitReq_17_54;
  assign compressDataVec_hitReq_17_54 = _GEN_1771;
  wire          compressDataVec_hitReq_17_182;
  assign compressDataVec_hitReq_17_182 = _GEN_1771;
  wire          _GEN_1772 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h36;
  wire          compressDataVec_hitReq_18_54;
  assign compressDataVec_hitReq_18_54 = _GEN_1772;
  wire          compressDataVec_hitReq_18_182;
  assign compressDataVec_hitReq_18_182 = _GEN_1772;
  wire          _GEN_1773 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h36;
  wire          compressDataVec_hitReq_19_54;
  assign compressDataVec_hitReq_19_54 = _GEN_1773;
  wire          compressDataVec_hitReq_19_182;
  assign compressDataVec_hitReq_19_182 = _GEN_1773;
  wire          _GEN_1774 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h36;
  wire          compressDataVec_hitReq_20_54;
  assign compressDataVec_hitReq_20_54 = _GEN_1774;
  wire          compressDataVec_hitReq_20_182;
  assign compressDataVec_hitReq_20_182 = _GEN_1774;
  wire          _GEN_1775 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h36;
  wire          compressDataVec_hitReq_21_54;
  assign compressDataVec_hitReq_21_54 = _GEN_1775;
  wire          compressDataVec_hitReq_21_182;
  assign compressDataVec_hitReq_21_182 = _GEN_1775;
  wire          _GEN_1776 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h36;
  wire          compressDataVec_hitReq_22_54;
  assign compressDataVec_hitReq_22_54 = _GEN_1776;
  wire          compressDataVec_hitReq_22_182;
  assign compressDataVec_hitReq_22_182 = _GEN_1776;
  wire          _GEN_1777 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h36;
  wire          compressDataVec_hitReq_23_54;
  assign compressDataVec_hitReq_23_54 = _GEN_1777;
  wire          compressDataVec_hitReq_23_182;
  assign compressDataVec_hitReq_23_182 = _GEN_1777;
  wire          _GEN_1778 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h36;
  wire          compressDataVec_hitReq_24_54;
  assign compressDataVec_hitReq_24_54 = _GEN_1778;
  wire          compressDataVec_hitReq_24_182;
  assign compressDataVec_hitReq_24_182 = _GEN_1778;
  wire          _GEN_1779 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h36;
  wire          compressDataVec_hitReq_25_54;
  assign compressDataVec_hitReq_25_54 = _GEN_1779;
  wire          compressDataVec_hitReq_25_182;
  assign compressDataVec_hitReq_25_182 = _GEN_1779;
  wire          _GEN_1780 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h36;
  wire          compressDataVec_hitReq_26_54;
  assign compressDataVec_hitReq_26_54 = _GEN_1780;
  wire          compressDataVec_hitReq_26_182;
  assign compressDataVec_hitReq_26_182 = _GEN_1780;
  wire          _GEN_1781 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h36;
  wire          compressDataVec_hitReq_27_54;
  assign compressDataVec_hitReq_27_54 = _GEN_1781;
  wire          compressDataVec_hitReq_27_182;
  assign compressDataVec_hitReq_27_182 = _GEN_1781;
  wire          _GEN_1782 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h36;
  wire          compressDataVec_hitReq_28_54;
  assign compressDataVec_hitReq_28_54 = _GEN_1782;
  wire          compressDataVec_hitReq_28_182;
  assign compressDataVec_hitReq_28_182 = _GEN_1782;
  wire          _GEN_1783 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h36;
  wire          compressDataVec_hitReq_29_54;
  assign compressDataVec_hitReq_29_54 = _GEN_1783;
  wire          compressDataVec_hitReq_29_182;
  assign compressDataVec_hitReq_29_182 = _GEN_1783;
  wire          _GEN_1784 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h36;
  wire          compressDataVec_hitReq_30_54;
  assign compressDataVec_hitReq_30_54 = _GEN_1784;
  wire          compressDataVec_hitReq_30_182;
  assign compressDataVec_hitReq_30_182 = _GEN_1784;
  wire          _GEN_1785 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h36;
  wire          compressDataVec_hitReq_31_54;
  assign compressDataVec_hitReq_31_54 = _GEN_1785;
  wire          compressDataVec_hitReq_31_182;
  assign compressDataVec_hitReq_31_182 = _GEN_1785;
  wire          compressDataVec_hitReq_32_54 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h36;
  wire          compressDataVec_hitReq_33_54 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h36;
  wire          compressDataVec_hitReq_34_54 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h36;
  wire          compressDataVec_hitReq_35_54 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h36;
  wire          compressDataVec_hitReq_36_54 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h36;
  wire          compressDataVec_hitReq_37_54 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h36;
  wire          compressDataVec_hitReq_38_54 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h36;
  wire          compressDataVec_hitReq_39_54 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h36;
  wire          compressDataVec_hitReq_40_54 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h36;
  wire          compressDataVec_hitReq_41_54 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h36;
  wire          compressDataVec_hitReq_42_54 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h36;
  wire          compressDataVec_hitReq_43_54 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h36;
  wire          compressDataVec_hitReq_44_54 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h36;
  wire          compressDataVec_hitReq_45_54 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h36;
  wire          compressDataVec_hitReq_46_54 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h36;
  wire          compressDataVec_hitReq_47_54 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h36;
  wire          compressDataVec_hitReq_48_54 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h36;
  wire          compressDataVec_hitReq_49_54 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h36;
  wire          compressDataVec_hitReq_50_54 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h36;
  wire          compressDataVec_hitReq_51_54 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h36;
  wire          compressDataVec_hitReq_52_54 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h36;
  wire          compressDataVec_hitReq_53_54 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h36;
  wire          compressDataVec_hitReq_54_54 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h36;
  wire          compressDataVec_hitReq_55_54 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h36;
  wire          compressDataVec_hitReq_56_54 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h36;
  wire          compressDataVec_hitReq_57_54 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h36;
  wire          compressDataVec_hitReq_58_54 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h36;
  wire          compressDataVec_hitReq_59_54 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h36;
  wire          compressDataVec_hitReq_60_54 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h36;
  wire          compressDataVec_hitReq_61_54 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h36;
  wire          compressDataVec_hitReq_62_54 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h36;
  wire          compressDataVec_hitReq_63_54 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h36;
  wire [7:0]    compressDataVec_selectReqData_54 =
    (compressDataVec_hitReq_0_54 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_54 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_54 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_54 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_54 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_54 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_54 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_54 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_54 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_54 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_54 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_54 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_54 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_54 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_54 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_54 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_54 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_54 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_54 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_54 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_54 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_54 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_54 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_54 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_54 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_54 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_54 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_54 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_54 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_54 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_54 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_54 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_54 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_54 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_54 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_54 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_54 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_54 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_54 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_54 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_54 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_54 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_54 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_54 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_54 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_54 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_54 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_54 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_54 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_54 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_54 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_54 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_54 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_54 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_54 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_54 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_54 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_54 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_54 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_54 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_54 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_54 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_54 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_54 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_54 = tailCount > 6'h36;
  wire          _GEN_1786 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h37;
  wire          compressDataVec_hitReq_0_55;
  assign compressDataVec_hitReq_0_55 = _GEN_1786;
  wire          compressDataVec_hitReq_0_183;
  assign compressDataVec_hitReq_0_183 = _GEN_1786;
  wire          _GEN_1787 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h37;
  wire          compressDataVec_hitReq_1_55;
  assign compressDataVec_hitReq_1_55 = _GEN_1787;
  wire          compressDataVec_hitReq_1_183;
  assign compressDataVec_hitReq_1_183 = _GEN_1787;
  wire          _GEN_1788 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h37;
  wire          compressDataVec_hitReq_2_55;
  assign compressDataVec_hitReq_2_55 = _GEN_1788;
  wire          compressDataVec_hitReq_2_183;
  assign compressDataVec_hitReq_2_183 = _GEN_1788;
  wire          _GEN_1789 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h37;
  wire          compressDataVec_hitReq_3_55;
  assign compressDataVec_hitReq_3_55 = _GEN_1789;
  wire          compressDataVec_hitReq_3_183;
  assign compressDataVec_hitReq_3_183 = _GEN_1789;
  wire          _GEN_1790 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h37;
  wire          compressDataVec_hitReq_4_55;
  assign compressDataVec_hitReq_4_55 = _GEN_1790;
  wire          compressDataVec_hitReq_4_183;
  assign compressDataVec_hitReq_4_183 = _GEN_1790;
  wire          _GEN_1791 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h37;
  wire          compressDataVec_hitReq_5_55;
  assign compressDataVec_hitReq_5_55 = _GEN_1791;
  wire          compressDataVec_hitReq_5_183;
  assign compressDataVec_hitReq_5_183 = _GEN_1791;
  wire          _GEN_1792 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h37;
  wire          compressDataVec_hitReq_6_55;
  assign compressDataVec_hitReq_6_55 = _GEN_1792;
  wire          compressDataVec_hitReq_6_183;
  assign compressDataVec_hitReq_6_183 = _GEN_1792;
  wire          _GEN_1793 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h37;
  wire          compressDataVec_hitReq_7_55;
  assign compressDataVec_hitReq_7_55 = _GEN_1793;
  wire          compressDataVec_hitReq_7_183;
  assign compressDataVec_hitReq_7_183 = _GEN_1793;
  wire          _GEN_1794 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h37;
  wire          compressDataVec_hitReq_8_55;
  assign compressDataVec_hitReq_8_55 = _GEN_1794;
  wire          compressDataVec_hitReq_8_183;
  assign compressDataVec_hitReq_8_183 = _GEN_1794;
  wire          _GEN_1795 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h37;
  wire          compressDataVec_hitReq_9_55;
  assign compressDataVec_hitReq_9_55 = _GEN_1795;
  wire          compressDataVec_hitReq_9_183;
  assign compressDataVec_hitReq_9_183 = _GEN_1795;
  wire          _GEN_1796 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h37;
  wire          compressDataVec_hitReq_10_55;
  assign compressDataVec_hitReq_10_55 = _GEN_1796;
  wire          compressDataVec_hitReq_10_183;
  assign compressDataVec_hitReq_10_183 = _GEN_1796;
  wire          _GEN_1797 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h37;
  wire          compressDataVec_hitReq_11_55;
  assign compressDataVec_hitReq_11_55 = _GEN_1797;
  wire          compressDataVec_hitReq_11_183;
  assign compressDataVec_hitReq_11_183 = _GEN_1797;
  wire          _GEN_1798 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h37;
  wire          compressDataVec_hitReq_12_55;
  assign compressDataVec_hitReq_12_55 = _GEN_1798;
  wire          compressDataVec_hitReq_12_183;
  assign compressDataVec_hitReq_12_183 = _GEN_1798;
  wire          _GEN_1799 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h37;
  wire          compressDataVec_hitReq_13_55;
  assign compressDataVec_hitReq_13_55 = _GEN_1799;
  wire          compressDataVec_hitReq_13_183;
  assign compressDataVec_hitReq_13_183 = _GEN_1799;
  wire          _GEN_1800 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h37;
  wire          compressDataVec_hitReq_14_55;
  assign compressDataVec_hitReq_14_55 = _GEN_1800;
  wire          compressDataVec_hitReq_14_183;
  assign compressDataVec_hitReq_14_183 = _GEN_1800;
  wire          _GEN_1801 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h37;
  wire          compressDataVec_hitReq_15_55;
  assign compressDataVec_hitReq_15_55 = _GEN_1801;
  wire          compressDataVec_hitReq_15_183;
  assign compressDataVec_hitReq_15_183 = _GEN_1801;
  wire          _GEN_1802 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h37;
  wire          compressDataVec_hitReq_16_55;
  assign compressDataVec_hitReq_16_55 = _GEN_1802;
  wire          compressDataVec_hitReq_16_183;
  assign compressDataVec_hitReq_16_183 = _GEN_1802;
  wire          _GEN_1803 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h37;
  wire          compressDataVec_hitReq_17_55;
  assign compressDataVec_hitReq_17_55 = _GEN_1803;
  wire          compressDataVec_hitReq_17_183;
  assign compressDataVec_hitReq_17_183 = _GEN_1803;
  wire          _GEN_1804 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h37;
  wire          compressDataVec_hitReq_18_55;
  assign compressDataVec_hitReq_18_55 = _GEN_1804;
  wire          compressDataVec_hitReq_18_183;
  assign compressDataVec_hitReq_18_183 = _GEN_1804;
  wire          _GEN_1805 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h37;
  wire          compressDataVec_hitReq_19_55;
  assign compressDataVec_hitReq_19_55 = _GEN_1805;
  wire          compressDataVec_hitReq_19_183;
  assign compressDataVec_hitReq_19_183 = _GEN_1805;
  wire          _GEN_1806 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h37;
  wire          compressDataVec_hitReq_20_55;
  assign compressDataVec_hitReq_20_55 = _GEN_1806;
  wire          compressDataVec_hitReq_20_183;
  assign compressDataVec_hitReq_20_183 = _GEN_1806;
  wire          _GEN_1807 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h37;
  wire          compressDataVec_hitReq_21_55;
  assign compressDataVec_hitReq_21_55 = _GEN_1807;
  wire          compressDataVec_hitReq_21_183;
  assign compressDataVec_hitReq_21_183 = _GEN_1807;
  wire          _GEN_1808 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h37;
  wire          compressDataVec_hitReq_22_55;
  assign compressDataVec_hitReq_22_55 = _GEN_1808;
  wire          compressDataVec_hitReq_22_183;
  assign compressDataVec_hitReq_22_183 = _GEN_1808;
  wire          _GEN_1809 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h37;
  wire          compressDataVec_hitReq_23_55;
  assign compressDataVec_hitReq_23_55 = _GEN_1809;
  wire          compressDataVec_hitReq_23_183;
  assign compressDataVec_hitReq_23_183 = _GEN_1809;
  wire          _GEN_1810 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h37;
  wire          compressDataVec_hitReq_24_55;
  assign compressDataVec_hitReq_24_55 = _GEN_1810;
  wire          compressDataVec_hitReq_24_183;
  assign compressDataVec_hitReq_24_183 = _GEN_1810;
  wire          _GEN_1811 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h37;
  wire          compressDataVec_hitReq_25_55;
  assign compressDataVec_hitReq_25_55 = _GEN_1811;
  wire          compressDataVec_hitReq_25_183;
  assign compressDataVec_hitReq_25_183 = _GEN_1811;
  wire          _GEN_1812 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h37;
  wire          compressDataVec_hitReq_26_55;
  assign compressDataVec_hitReq_26_55 = _GEN_1812;
  wire          compressDataVec_hitReq_26_183;
  assign compressDataVec_hitReq_26_183 = _GEN_1812;
  wire          _GEN_1813 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h37;
  wire          compressDataVec_hitReq_27_55;
  assign compressDataVec_hitReq_27_55 = _GEN_1813;
  wire          compressDataVec_hitReq_27_183;
  assign compressDataVec_hitReq_27_183 = _GEN_1813;
  wire          _GEN_1814 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h37;
  wire          compressDataVec_hitReq_28_55;
  assign compressDataVec_hitReq_28_55 = _GEN_1814;
  wire          compressDataVec_hitReq_28_183;
  assign compressDataVec_hitReq_28_183 = _GEN_1814;
  wire          _GEN_1815 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h37;
  wire          compressDataVec_hitReq_29_55;
  assign compressDataVec_hitReq_29_55 = _GEN_1815;
  wire          compressDataVec_hitReq_29_183;
  assign compressDataVec_hitReq_29_183 = _GEN_1815;
  wire          _GEN_1816 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h37;
  wire          compressDataVec_hitReq_30_55;
  assign compressDataVec_hitReq_30_55 = _GEN_1816;
  wire          compressDataVec_hitReq_30_183;
  assign compressDataVec_hitReq_30_183 = _GEN_1816;
  wire          _GEN_1817 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h37;
  wire          compressDataVec_hitReq_31_55;
  assign compressDataVec_hitReq_31_55 = _GEN_1817;
  wire          compressDataVec_hitReq_31_183;
  assign compressDataVec_hitReq_31_183 = _GEN_1817;
  wire          compressDataVec_hitReq_32_55 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h37;
  wire          compressDataVec_hitReq_33_55 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h37;
  wire          compressDataVec_hitReq_34_55 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h37;
  wire          compressDataVec_hitReq_35_55 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h37;
  wire          compressDataVec_hitReq_36_55 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h37;
  wire          compressDataVec_hitReq_37_55 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h37;
  wire          compressDataVec_hitReq_38_55 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h37;
  wire          compressDataVec_hitReq_39_55 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h37;
  wire          compressDataVec_hitReq_40_55 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h37;
  wire          compressDataVec_hitReq_41_55 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h37;
  wire          compressDataVec_hitReq_42_55 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h37;
  wire          compressDataVec_hitReq_43_55 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h37;
  wire          compressDataVec_hitReq_44_55 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h37;
  wire          compressDataVec_hitReq_45_55 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h37;
  wire          compressDataVec_hitReq_46_55 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h37;
  wire          compressDataVec_hitReq_47_55 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h37;
  wire          compressDataVec_hitReq_48_55 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h37;
  wire          compressDataVec_hitReq_49_55 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h37;
  wire          compressDataVec_hitReq_50_55 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h37;
  wire          compressDataVec_hitReq_51_55 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h37;
  wire          compressDataVec_hitReq_52_55 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h37;
  wire          compressDataVec_hitReq_53_55 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h37;
  wire          compressDataVec_hitReq_54_55 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h37;
  wire          compressDataVec_hitReq_55_55 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h37;
  wire          compressDataVec_hitReq_56_55 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h37;
  wire          compressDataVec_hitReq_57_55 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h37;
  wire          compressDataVec_hitReq_58_55 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h37;
  wire          compressDataVec_hitReq_59_55 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h37;
  wire          compressDataVec_hitReq_60_55 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h37;
  wire          compressDataVec_hitReq_61_55 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h37;
  wire          compressDataVec_hitReq_62_55 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h37;
  wire          compressDataVec_hitReq_63_55 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h37;
  wire [7:0]    compressDataVec_selectReqData_55 =
    (compressDataVec_hitReq_0_55 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_55 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_55 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_55 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_55 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_55 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_55 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_55 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_55 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_55 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_55 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_55 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_55 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_55 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_55 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_55 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_55 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_55 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_55 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_55 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_55 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_55 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_55 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_55 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_55 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_55 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_55 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_55 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_55 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_55 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_55 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_55 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_55 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_55 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_55 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_55 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_55 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_55 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_55 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_55 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_55 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_55 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_55 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_55 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_55 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_55 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_55 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_55 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_55 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_55 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_55 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_55 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_55 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_55 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_55 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_55 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_55 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_55 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_55 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_55 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_55 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_55 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_55 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_55 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_55 = tailCount > 6'h37;
  wire          _GEN_1818 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h38;
  wire          compressDataVec_hitReq_0_56;
  assign compressDataVec_hitReq_0_56 = _GEN_1818;
  wire          compressDataVec_hitReq_0_184;
  assign compressDataVec_hitReq_0_184 = _GEN_1818;
  wire          _GEN_1819 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h38;
  wire          compressDataVec_hitReq_1_56;
  assign compressDataVec_hitReq_1_56 = _GEN_1819;
  wire          compressDataVec_hitReq_1_184;
  assign compressDataVec_hitReq_1_184 = _GEN_1819;
  wire          _GEN_1820 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h38;
  wire          compressDataVec_hitReq_2_56;
  assign compressDataVec_hitReq_2_56 = _GEN_1820;
  wire          compressDataVec_hitReq_2_184;
  assign compressDataVec_hitReq_2_184 = _GEN_1820;
  wire          _GEN_1821 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h38;
  wire          compressDataVec_hitReq_3_56;
  assign compressDataVec_hitReq_3_56 = _GEN_1821;
  wire          compressDataVec_hitReq_3_184;
  assign compressDataVec_hitReq_3_184 = _GEN_1821;
  wire          _GEN_1822 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h38;
  wire          compressDataVec_hitReq_4_56;
  assign compressDataVec_hitReq_4_56 = _GEN_1822;
  wire          compressDataVec_hitReq_4_184;
  assign compressDataVec_hitReq_4_184 = _GEN_1822;
  wire          _GEN_1823 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h38;
  wire          compressDataVec_hitReq_5_56;
  assign compressDataVec_hitReq_5_56 = _GEN_1823;
  wire          compressDataVec_hitReq_5_184;
  assign compressDataVec_hitReq_5_184 = _GEN_1823;
  wire          _GEN_1824 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h38;
  wire          compressDataVec_hitReq_6_56;
  assign compressDataVec_hitReq_6_56 = _GEN_1824;
  wire          compressDataVec_hitReq_6_184;
  assign compressDataVec_hitReq_6_184 = _GEN_1824;
  wire          _GEN_1825 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h38;
  wire          compressDataVec_hitReq_7_56;
  assign compressDataVec_hitReq_7_56 = _GEN_1825;
  wire          compressDataVec_hitReq_7_184;
  assign compressDataVec_hitReq_7_184 = _GEN_1825;
  wire          _GEN_1826 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h38;
  wire          compressDataVec_hitReq_8_56;
  assign compressDataVec_hitReq_8_56 = _GEN_1826;
  wire          compressDataVec_hitReq_8_184;
  assign compressDataVec_hitReq_8_184 = _GEN_1826;
  wire          _GEN_1827 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h38;
  wire          compressDataVec_hitReq_9_56;
  assign compressDataVec_hitReq_9_56 = _GEN_1827;
  wire          compressDataVec_hitReq_9_184;
  assign compressDataVec_hitReq_9_184 = _GEN_1827;
  wire          _GEN_1828 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h38;
  wire          compressDataVec_hitReq_10_56;
  assign compressDataVec_hitReq_10_56 = _GEN_1828;
  wire          compressDataVec_hitReq_10_184;
  assign compressDataVec_hitReq_10_184 = _GEN_1828;
  wire          _GEN_1829 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h38;
  wire          compressDataVec_hitReq_11_56;
  assign compressDataVec_hitReq_11_56 = _GEN_1829;
  wire          compressDataVec_hitReq_11_184;
  assign compressDataVec_hitReq_11_184 = _GEN_1829;
  wire          _GEN_1830 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h38;
  wire          compressDataVec_hitReq_12_56;
  assign compressDataVec_hitReq_12_56 = _GEN_1830;
  wire          compressDataVec_hitReq_12_184;
  assign compressDataVec_hitReq_12_184 = _GEN_1830;
  wire          _GEN_1831 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h38;
  wire          compressDataVec_hitReq_13_56;
  assign compressDataVec_hitReq_13_56 = _GEN_1831;
  wire          compressDataVec_hitReq_13_184;
  assign compressDataVec_hitReq_13_184 = _GEN_1831;
  wire          _GEN_1832 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h38;
  wire          compressDataVec_hitReq_14_56;
  assign compressDataVec_hitReq_14_56 = _GEN_1832;
  wire          compressDataVec_hitReq_14_184;
  assign compressDataVec_hitReq_14_184 = _GEN_1832;
  wire          _GEN_1833 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h38;
  wire          compressDataVec_hitReq_15_56;
  assign compressDataVec_hitReq_15_56 = _GEN_1833;
  wire          compressDataVec_hitReq_15_184;
  assign compressDataVec_hitReq_15_184 = _GEN_1833;
  wire          _GEN_1834 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h38;
  wire          compressDataVec_hitReq_16_56;
  assign compressDataVec_hitReq_16_56 = _GEN_1834;
  wire          compressDataVec_hitReq_16_184;
  assign compressDataVec_hitReq_16_184 = _GEN_1834;
  wire          _GEN_1835 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h38;
  wire          compressDataVec_hitReq_17_56;
  assign compressDataVec_hitReq_17_56 = _GEN_1835;
  wire          compressDataVec_hitReq_17_184;
  assign compressDataVec_hitReq_17_184 = _GEN_1835;
  wire          _GEN_1836 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h38;
  wire          compressDataVec_hitReq_18_56;
  assign compressDataVec_hitReq_18_56 = _GEN_1836;
  wire          compressDataVec_hitReq_18_184;
  assign compressDataVec_hitReq_18_184 = _GEN_1836;
  wire          _GEN_1837 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h38;
  wire          compressDataVec_hitReq_19_56;
  assign compressDataVec_hitReq_19_56 = _GEN_1837;
  wire          compressDataVec_hitReq_19_184;
  assign compressDataVec_hitReq_19_184 = _GEN_1837;
  wire          _GEN_1838 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h38;
  wire          compressDataVec_hitReq_20_56;
  assign compressDataVec_hitReq_20_56 = _GEN_1838;
  wire          compressDataVec_hitReq_20_184;
  assign compressDataVec_hitReq_20_184 = _GEN_1838;
  wire          _GEN_1839 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h38;
  wire          compressDataVec_hitReq_21_56;
  assign compressDataVec_hitReq_21_56 = _GEN_1839;
  wire          compressDataVec_hitReq_21_184;
  assign compressDataVec_hitReq_21_184 = _GEN_1839;
  wire          _GEN_1840 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h38;
  wire          compressDataVec_hitReq_22_56;
  assign compressDataVec_hitReq_22_56 = _GEN_1840;
  wire          compressDataVec_hitReq_22_184;
  assign compressDataVec_hitReq_22_184 = _GEN_1840;
  wire          _GEN_1841 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h38;
  wire          compressDataVec_hitReq_23_56;
  assign compressDataVec_hitReq_23_56 = _GEN_1841;
  wire          compressDataVec_hitReq_23_184;
  assign compressDataVec_hitReq_23_184 = _GEN_1841;
  wire          _GEN_1842 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h38;
  wire          compressDataVec_hitReq_24_56;
  assign compressDataVec_hitReq_24_56 = _GEN_1842;
  wire          compressDataVec_hitReq_24_184;
  assign compressDataVec_hitReq_24_184 = _GEN_1842;
  wire          _GEN_1843 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h38;
  wire          compressDataVec_hitReq_25_56;
  assign compressDataVec_hitReq_25_56 = _GEN_1843;
  wire          compressDataVec_hitReq_25_184;
  assign compressDataVec_hitReq_25_184 = _GEN_1843;
  wire          _GEN_1844 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h38;
  wire          compressDataVec_hitReq_26_56;
  assign compressDataVec_hitReq_26_56 = _GEN_1844;
  wire          compressDataVec_hitReq_26_184;
  assign compressDataVec_hitReq_26_184 = _GEN_1844;
  wire          _GEN_1845 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h38;
  wire          compressDataVec_hitReq_27_56;
  assign compressDataVec_hitReq_27_56 = _GEN_1845;
  wire          compressDataVec_hitReq_27_184;
  assign compressDataVec_hitReq_27_184 = _GEN_1845;
  wire          _GEN_1846 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h38;
  wire          compressDataVec_hitReq_28_56;
  assign compressDataVec_hitReq_28_56 = _GEN_1846;
  wire          compressDataVec_hitReq_28_184;
  assign compressDataVec_hitReq_28_184 = _GEN_1846;
  wire          _GEN_1847 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h38;
  wire          compressDataVec_hitReq_29_56;
  assign compressDataVec_hitReq_29_56 = _GEN_1847;
  wire          compressDataVec_hitReq_29_184;
  assign compressDataVec_hitReq_29_184 = _GEN_1847;
  wire          _GEN_1848 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h38;
  wire          compressDataVec_hitReq_30_56;
  assign compressDataVec_hitReq_30_56 = _GEN_1848;
  wire          compressDataVec_hitReq_30_184;
  assign compressDataVec_hitReq_30_184 = _GEN_1848;
  wire          _GEN_1849 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h38;
  wire          compressDataVec_hitReq_31_56;
  assign compressDataVec_hitReq_31_56 = _GEN_1849;
  wire          compressDataVec_hitReq_31_184;
  assign compressDataVec_hitReq_31_184 = _GEN_1849;
  wire          compressDataVec_hitReq_32_56 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h38;
  wire          compressDataVec_hitReq_33_56 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h38;
  wire          compressDataVec_hitReq_34_56 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h38;
  wire          compressDataVec_hitReq_35_56 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h38;
  wire          compressDataVec_hitReq_36_56 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h38;
  wire          compressDataVec_hitReq_37_56 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h38;
  wire          compressDataVec_hitReq_38_56 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h38;
  wire          compressDataVec_hitReq_39_56 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h38;
  wire          compressDataVec_hitReq_40_56 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h38;
  wire          compressDataVec_hitReq_41_56 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h38;
  wire          compressDataVec_hitReq_42_56 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h38;
  wire          compressDataVec_hitReq_43_56 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h38;
  wire          compressDataVec_hitReq_44_56 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h38;
  wire          compressDataVec_hitReq_45_56 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h38;
  wire          compressDataVec_hitReq_46_56 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h38;
  wire          compressDataVec_hitReq_47_56 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h38;
  wire          compressDataVec_hitReq_48_56 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h38;
  wire          compressDataVec_hitReq_49_56 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h38;
  wire          compressDataVec_hitReq_50_56 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h38;
  wire          compressDataVec_hitReq_51_56 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h38;
  wire          compressDataVec_hitReq_52_56 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h38;
  wire          compressDataVec_hitReq_53_56 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h38;
  wire          compressDataVec_hitReq_54_56 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h38;
  wire          compressDataVec_hitReq_55_56 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h38;
  wire          compressDataVec_hitReq_56_56 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h38;
  wire          compressDataVec_hitReq_57_56 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h38;
  wire          compressDataVec_hitReq_58_56 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h38;
  wire          compressDataVec_hitReq_59_56 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h38;
  wire          compressDataVec_hitReq_60_56 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h38;
  wire          compressDataVec_hitReq_61_56 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h38;
  wire          compressDataVec_hitReq_62_56 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h38;
  wire          compressDataVec_hitReq_63_56 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h38;
  wire [7:0]    compressDataVec_selectReqData_56 =
    (compressDataVec_hitReq_0_56 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_56 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_56 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_56 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_56 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_56 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_56 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_56 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_56 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_56 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_56 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_56 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_56 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_56 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_56 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_56 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_56 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_56 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_56 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_56 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_56 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_56 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_56 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_56 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_56 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_56 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_56 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_56 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_56 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_56 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_56 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_56 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_56 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_56 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_56 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_56 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_56 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_56 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_56 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_56 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_56 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_56 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_56 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_56 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_56 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_56 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_56 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_56 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_56 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_56 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_56 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_56 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_56 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_56 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_56 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_56 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_56 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_56 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_56 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_56 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_56 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_56 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_56 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_56 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_56 = tailCount > 6'h38;
  wire          _GEN_1850 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h39;
  wire          compressDataVec_hitReq_0_57;
  assign compressDataVec_hitReq_0_57 = _GEN_1850;
  wire          compressDataVec_hitReq_0_185;
  assign compressDataVec_hitReq_0_185 = _GEN_1850;
  wire          _GEN_1851 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h39;
  wire          compressDataVec_hitReq_1_57;
  assign compressDataVec_hitReq_1_57 = _GEN_1851;
  wire          compressDataVec_hitReq_1_185;
  assign compressDataVec_hitReq_1_185 = _GEN_1851;
  wire          _GEN_1852 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h39;
  wire          compressDataVec_hitReq_2_57;
  assign compressDataVec_hitReq_2_57 = _GEN_1852;
  wire          compressDataVec_hitReq_2_185;
  assign compressDataVec_hitReq_2_185 = _GEN_1852;
  wire          _GEN_1853 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h39;
  wire          compressDataVec_hitReq_3_57;
  assign compressDataVec_hitReq_3_57 = _GEN_1853;
  wire          compressDataVec_hitReq_3_185;
  assign compressDataVec_hitReq_3_185 = _GEN_1853;
  wire          _GEN_1854 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h39;
  wire          compressDataVec_hitReq_4_57;
  assign compressDataVec_hitReq_4_57 = _GEN_1854;
  wire          compressDataVec_hitReq_4_185;
  assign compressDataVec_hitReq_4_185 = _GEN_1854;
  wire          _GEN_1855 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h39;
  wire          compressDataVec_hitReq_5_57;
  assign compressDataVec_hitReq_5_57 = _GEN_1855;
  wire          compressDataVec_hitReq_5_185;
  assign compressDataVec_hitReq_5_185 = _GEN_1855;
  wire          _GEN_1856 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h39;
  wire          compressDataVec_hitReq_6_57;
  assign compressDataVec_hitReq_6_57 = _GEN_1856;
  wire          compressDataVec_hitReq_6_185;
  assign compressDataVec_hitReq_6_185 = _GEN_1856;
  wire          _GEN_1857 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h39;
  wire          compressDataVec_hitReq_7_57;
  assign compressDataVec_hitReq_7_57 = _GEN_1857;
  wire          compressDataVec_hitReq_7_185;
  assign compressDataVec_hitReq_7_185 = _GEN_1857;
  wire          _GEN_1858 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h39;
  wire          compressDataVec_hitReq_8_57;
  assign compressDataVec_hitReq_8_57 = _GEN_1858;
  wire          compressDataVec_hitReq_8_185;
  assign compressDataVec_hitReq_8_185 = _GEN_1858;
  wire          _GEN_1859 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h39;
  wire          compressDataVec_hitReq_9_57;
  assign compressDataVec_hitReq_9_57 = _GEN_1859;
  wire          compressDataVec_hitReq_9_185;
  assign compressDataVec_hitReq_9_185 = _GEN_1859;
  wire          _GEN_1860 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h39;
  wire          compressDataVec_hitReq_10_57;
  assign compressDataVec_hitReq_10_57 = _GEN_1860;
  wire          compressDataVec_hitReq_10_185;
  assign compressDataVec_hitReq_10_185 = _GEN_1860;
  wire          _GEN_1861 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h39;
  wire          compressDataVec_hitReq_11_57;
  assign compressDataVec_hitReq_11_57 = _GEN_1861;
  wire          compressDataVec_hitReq_11_185;
  assign compressDataVec_hitReq_11_185 = _GEN_1861;
  wire          _GEN_1862 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h39;
  wire          compressDataVec_hitReq_12_57;
  assign compressDataVec_hitReq_12_57 = _GEN_1862;
  wire          compressDataVec_hitReq_12_185;
  assign compressDataVec_hitReq_12_185 = _GEN_1862;
  wire          _GEN_1863 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h39;
  wire          compressDataVec_hitReq_13_57;
  assign compressDataVec_hitReq_13_57 = _GEN_1863;
  wire          compressDataVec_hitReq_13_185;
  assign compressDataVec_hitReq_13_185 = _GEN_1863;
  wire          _GEN_1864 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h39;
  wire          compressDataVec_hitReq_14_57;
  assign compressDataVec_hitReq_14_57 = _GEN_1864;
  wire          compressDataVec_hitReq_14_185;
  assign compressDataVec_hitReq_14_185 = _GEN_1864;
  wire          _GEN_1865 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h39;
  wire          compressDataVec_hitReq_15_57;
  assign compressDataVec_hitReq_15_57 = _GEN_1865;
  wire          compressDataVec_hitReq_15_185;
  assign compressDataVec_hitReq_15_185 = _GEN_1865;
  wire          _GEN_1866 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h39;
  wire          compressDataVec_hitReq_16_57;
  assign compressDataVec_hitReq_16_57 = _GEN_1866;
  wire          compressDataVec_hitReq_16_185;
  assign compressDataVec_hitReq_16_185 = _GEN_1866;
  wire          _GEN_1867 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h39;
  wire          compressDataVec_hitReq_17_57;
  assign compressDataVec_hitReq_17_57 = _GEN_1867;
  wire          compressDataVec_hitReq_17_185;
  assign compressDataVec_hitReq_17_185 = _GEN_1867;
  wire          _GEN_1868 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h39;
  wire          compressDataVec_hitReq_18_57;
  assign compressDataVec_hitReq_18_57 = _GEN_1868;
  wire          compressDataVec_hitReq_18_185;
  assign compressDataVec_hitReq_18_185 = _GEN_1868;
  wire          _GEN_1869 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h39;
  wire          compressDataVec_hitReq_19_57;
  assign compressDataVec_hitReq_19_57 = _GEN_1869;
  wire          compressDataVec_hitReq_19_185;
  assign compressDataVec_hitReq_19_185 = _GEN_1869;
  wire          _GEN_1870 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h39;
  wire          compressDataVec_hitReq_20_57;
  assign compressDataVec_hitReq_20_57 = _GEN_1870;
  wire          compressDataVec_hitReq_20_185;
  assign compressDataVec_hitReq_20_185 = _GEN_1870;
  wire          _GEN_1871 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h39;
  wire          compressDataVec_hitReq_21_57;
  assign compressDataVec_hitReq_21_57 = _GEN_1871;
  wire          compressDataVec_hitReq_21_185;
  assign compressDataVec_hitReq_21_185 = _GEN_1871;
  wire          _GEN_1872 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h39;
  wire          compressDataVec_hitReq_22_57;
  assign compressDataVec_hitReq_22_57 = _GEN_1872;
  wire          compressDataVec_hitReq_22_185;
  assign compressDataVec_hitReq_22_185 = _GEN_1872;
  wire          _GEN_1873 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h39;
  wire          compressDataVec_hitReq_23_57;
  assign compressDataVec_hitReq_23_57 = _GEN_1873;
  wire          compressDataVec_hitReq_23_185;
  assign compressDataVec_hitReq_23_185 = _GEN_1873;
  wire          _GEN_1874 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h39;
  wire          compressDataVec_hitReq_24_57;
  assign compressDataVec_hitReq_24_57 = _GEN_1874;
  wire          compressDataVec_hitReq_24_185;
  assign compressDataVec_hitReq_24_185 = _GEN_1874;
  wire          _GEN_1875 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h39;
  wire          compressDataVec_hitReq_25_57;
  assign compressDataVec_hitReq_25_57 = _GEN_1875;
  wire          compressDataVec_hitReq_25_185;
  assign compressDataVec_hitReq_25_185 = _GEN_1875;
  wire          _GEN_1876 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h39;
  wire          compressDataVec_hitReq_26_57;
  assign compressDataVec_hitReq_26_57 = _GEN_1876;
  wire          compressDataVec_hitReq_26_185;
  assign compressDataVec_hitReq_26_185 = _GEN_1876;
  wire          _GEN_1877 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h39;
  wire          compressDataVec_hitReq_27_57;
  assign compressDataVec_hitReq_27_57 = _GEN_1877;
  wire          compressDataVec_hitReq_27_185;
  assign compressDataVec_hitReq_27_185 = _GEN_1877;
  wire          _GEN_1878 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h39;
  wire          compressDataVec_hitReq_28_57;
  assign compressDataVec_hitReq_28_57 = _GEN_1878;
  wire          compressDataVec_hitReq_28_185;
  assign compressDataVec_hitReq_28_185 = _GEN_1878;
  wire          _GEN_1879 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h39;
  wire          compressDataVec_hitReq_29_57;
  assign compressDataVec_hitReq_29_57 = _GEN_1879;
  wire          compressDataVec_hitReq_29_185;
  assign compressDataVec_hitReq_29_185 = _GEN_1879;
  wire          _GEN_1880 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h39;
  wire          compressDataVec_hitReq_30_57;
  assign compressDataVec_hitReq_30_57 = _GEN_1880;
  wire          compressDataVec_hitReq_30_185;
  assign compressDataVec_hitReq_30_185 = _GEN_1880;
  wire          _GEN_1881 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h39;
  wire          compressDataVec_hitReq_31_57;
  assign compressDataVec_hitReq_31_57 = _GEN_1881;
  wire          compressDataVec_hitReq_31_185;
  assign compressDataVec_hitReq_31_185 = _GEN_1881;
  wire          compressDataVec_hitReq_32_57 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h39;
  wire          compressDataVec_hitReq_33_57 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h39;
  wire          compressDataVec_hitReq_34_57 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h39;
  wire          compressDataVec_hitReq_35_57 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h39;
  wire          compressDataVec_hitReq_36_57 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h39;
  wire          compressDataVec_hitReq_37_57 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h39;
  wire          compressDataVec_hitReq_38_57 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h39;
  wire          compressDataVec_hitReq_39_57 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h39;
  wire          compressDataVec_hitReq_40_57 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h39;
  wire          compressDataVec_hitReq_41_57 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h39;
  wire          compressDataVec_hitReq_42_57 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h39;
  wire          compressDataVec_hitReq_43_57 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h39;
  wire          compressDataVec_hitReq_44_57 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h39;
  wire          compressDataVec_hitReq_45_57 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h39;
  wire          compressDataVec_hitReq_46_57 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h39;
  wire          compressDataVec_hitReq_47_57 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h39;
  wire          compressDataVec_hitReq_48_57 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h39;
  wire          compressDataVec_hitReq_49_57 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h39;
  wire          compressDataVec_hitReq_50_57 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h39;
  wire          compressDataVec_hitReq_51_57 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h39;
  wire          compressDataVec_hitReq_52_57 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h39;
  wire          compressDataVec_hitReq_53_57 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h39;
  wire          compressDataVec_hitReq_54_57 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h39;
  wire          compressDataVec_hitReq_55_57 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h39;
  wire          compressDataVec_hitReq_56_57 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h39;
  wire          compressDataVec_hitReq_57_57 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h39;
  wire          compressDataVec_hitReq_58_57 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h39;
  wire          compressDataVec_hitReq_59_57 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h39;
  wire          compressDataVec_hitReq_60_57 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h39;
  wire          compressDataVec_hitReq_61_57 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h39;
  wire          compressDataVec_hitReq_62_57 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h39;
  wire          compressDataVec_hitReq_63_57 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h39;
  wire [7:0]    compressDataVec_selectReqData_57 =
    (compressDataVec_hitReq_0_57 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_57 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_57 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_57 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_57 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_57 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_57 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_57 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_57 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_57 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_57 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_57 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_57 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_57 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_57 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_57 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_57 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_57 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_57 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_57 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_57 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_57 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_57 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_57 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_57 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_57 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_57 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_57 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_57 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_57 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_57 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_57 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_57 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_57 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_57 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_57 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_57 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_57 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_57 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_57 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_57 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_57 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_57 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_57 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_57 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_57 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_57 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_57 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_57 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_57 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_57 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_57 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_57 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_57 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_57 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_57 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_57 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_57 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_57 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_57 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_57 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_57 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_57 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_57 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_57 = tailCount > 6'h39;
  wire          _GEN_1882 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h3A;
  wire          compressDataVec_hitReq_0_58;
  assign compressDataVec_hitReq_0_58 = _GEN_1882;
  wire          compressDataVec_hitReq_0_186;
  assign compressDataVec_hitReq_0_186 = _GEN_1882;
  wire          _GEN_1883 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h3A;
  wire          compressDataVec_hitReq_1_58;
  assign compressDataVec_hitReq_1_58 = _GEN_1883;
  wire          compressDataVec_hitReq_1_186;
  assign compressDataVec_hitReq_1_186 = _GEN_1883;
  wire          _GEN_1884 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h3A;
  wire          compressDataVec_hitReq_2_58;
  assign compressDataVec_hitReq_2_58 = _GEN_1884;
  wire          compressDataVec_hitReq_2_186;
  assign compressDataVec_hitReq_2_186 = _GEN_1884;
  wire          _GEN_1885 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h3A;
  wire          compressDataVec_hitReq_3_58;
  assign compressDataVec_hitReq_3_58 = _GEN_1885;
  wire          compressDataVec_hitReq_3_186;
  assign compressDataVec_hitReq_3_186 = _GEN_1885;
  wire          _GEN_1886 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h3A;
  wire          compressDataVec_hitReq_4_58;
  assign compressDataVec_hitReq_4_58 = _GEN_1886;
  wire          compressDataVec_hitReq_4_186;
  assign compressDataVec_hitReq_4_186 = _GEN_1886;
  wire          _GEN_1887 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h3A;
  wire          compressDataVec_hitReq_5_58;
  assign compressDataVec_hitReq_5_58 = _GEN_1887;
  wire          compressDataVec_hitReq_5_186;
  assign compressDataVec_hitReq_5_186 = _GEN_1887;
  wire          _GEN_1888 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h3A;
  wire          compressDataVec_hitReq_6_58;
  assign compressDataVec_hitReq_6_58 = _GEN_1888;
  wire          compressDataVec_hitReq_6_186;
  assign compressDataVec_hitReq_6_186 = _GEN_1888;
  wire          _GEN_1889 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h3A;
  wire          compressDataVec_hitReq_7_58;
  assign compressDataVec_hitReq_7_58 = _GEN_1889;
  wire          compressDataVec_hitReq_7_186;
  assign compressDataVec_hitReq_7_186 = _GEN_1889;
  wire          _GEN_1890 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h3A;
  wire          compressDataVec_hitReq_8_58;
  assign compressDataVec_hitReq_8_58 = _GEN_1890;
  wire          compressDataVec_hitReq_8_186;
  assign compressDataVec_hitReq_8_186 = _GEN_1890;
  wire          _GEN_1891 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h3A;
  wire          compressDataVec_hitReq_9_58;
  assign compressDataVec_hitReq_9_58 = _GEN_1891;
  wire          compressDataVec_hitReq_9_186;
  assign compressDataVec_hitReq_9_186 = _GEN_1891;
  wire          _GEN_1892 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h3A;
  wire          compressDataVec_hitReq_10_58;
  assign compressDataVec_hitReq_10_58 = _GEN_1892;
  wire          compressDataVec_hitReq_10_186;
  assign compressDataVec_hitReq_10_186 = _GEN_1892;
  wire          _GEN_1893 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h3A;
  wire          compressDataVec_hitReq_11_58;
  assign compressDataVec_hitReq_11_58 = _GEN_1893;
  wire          compressDataVec_hitReq_11_186;
  assign compressDataVec_hitReq_11_186 = _GEN_1893;
  wire          _GEN_1894 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h3A;
  wire          compressDataVec_hitReq_12_58;
  assign compressDataVec_hitReq_12_58 = _GEN_1894;
  wire          compressDataVec_hitReq_12_186;
  assign compressDataVec_hitReq_12_186 = _GEN_1894;
  wire          _GEN_1895 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h3A;
  wire          compressDataVec_hitReq_13_58;
  assign compressDataVec_hitReq_13_58 = _GEN_1895;
  wire          compressDataVec_hitReq_13_186;
  assign compressDataVec_hitReq_13_186 = _GEN_1895;
  wire          _GEN_1896 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h3A;
  wire          compressDataVec_hitReq_14_58;
  assign compressDataVec_hitReq_14_58 = _GEN_1896;
  wire          compressDataVec_hitReq_14_186;
  assign compressDataVec_hitReq_14_186 = _GEN_1896;
  wire          _GEN_1897 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h3A;
  wire          compressDataVec_hitReq_15_58;
  assign compressDataVec_hitReq_15_58 = _GEN_1897;
  wire          compressDataVec_hitReq_15_186;
  assign compressDataVec_hitReq_15_186 = _GEN_1897;
  wire          _GEN_1898 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h3A;
  wire          compressDataVec_hitReq_16_58;
  assign compressDataVec_hitReq_16_58 = _GEN_1898;
  wire          compressDataVec_hitReq_16_186;
  assign compressDataVec_hitReq_16_186 = _GEN_1898;
  wire          _GEN_1899 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h3A;
  wire          compressDataVec_hitReq_17_58;
  assign compressDataVec_hitReq_17_58 = _GEN_1899;
  wire          compressDataVec_hitReq_17_186;
  assign compressDataVec_hitReq_17_186 = _GEN_1899;
  wire          _GEN_1900 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h3A;
  wire          compressDataVec_hitReq_18_58;
  assign compressDataVec_hitReq_18_58 = _GEN_1900;
  wire          compressDataVec_hitReq_18_186;
  assign compressDataVec_hitReq_18_186 = _GEN_1900;
  wire          _GEN_1901 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h3A;
  wire          compressDataVec_hitReq_19_58;
  assign compressDataVec_hitReq_19_58 = _GEN_1901;
  wire          compressDataVec_hitReq_19_186;
  assign compressDataVec_hitReq_19_186 = _GEN_1901;
  wire          _GEN_1902 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h3A;
  wire          compressDataVec_hitReq_20_58;
  assign compressDataVec_hitReq_20_58 = _GEN_1902;
  wire          compressDataVec_hitReq_20_186;
  assign compressDataVec_hitReq_20_186 = _GEN_1902;
  wire          _GEN_1903 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h3A;
  wire          compressDataVec_hitReq_21_58;
  assign compressDataVec_hitReq_21_58 = _GEN_1903;
  wire          compressDataVec_hitReq_21_186;
  assign compressDataVec_hitReq_21_186 = _GEN_1903;
  wire          _GEN_1904 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h3A;
  wire          compressDataVec_hitReq_22_58;
  assign compressDataVec_hitReq_22_58 = _GEN_1904;
  wire          compressDataVec_hitReq_22_186;
  assign compressDataVec_hitReq_22_186 = _GEN_1904;
  wire          _GEN_1905 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h3A;
  wire          compressDataVec_hitReq_23_58;
  assign compressDataVec_hitReq_23_58 = _GEN_1905;
  wire          compressDataVec_hitReq_23_186;
  assign compressDataVec_hitReq_23_186 = _GEN_1905;
  wire          _GEN_1906 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h3A;
  wire          compressDataVec_hitReq_24_58;
  assign compressDataVec_hitReq_24_58 = _GEN_1906;
  wire          compressDataVec_hitReq_24_186;
  assign compressDataVec_hitReq_24_186 = _GEN_1906;
  wire          _GEN_1907 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h3A;
  wire          compressDataVec_hitReq_25_58;
  assign compressDataVec_hitReq_25_58 = _GEN_1907;
  wire          compressDataVec_hitReq_25_186;
  assign compressDataVec_hitReq_25_186 = _GEN_1907;
  wire          _GEN_1908 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h3A;
  wire          compressDataVec_hitReq_26_58;
  assign compressDataVec_hitReq_26_58 = _GEN_1908;
  wire          compressDataVec_hitReq_26_186;
  assign compressDataVec_hitReq_26_186 = _GEN_1908;
  wire          _GEN_1909 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h3A;
  wire          compressDataVec_hitReq_27_58;
  assign compressDataVec_hitReq_27_58 = _GEN_1909;
  wire          compressDataVec_hitReq_27_186;
  assign compressDataVec_hitReq_27_186 = _GEN_1909;
  wire          _GEN_1910 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h3A;
  wire          compressDataVec_hitReq_28_58;
  assign compressDataVec_hitReq_28_58 = _GEN_1910;
  wire          compressDataVec_hitReq_28_186;
  assign compressDataVec_hitReq_28_186 = _GEN_1910;
  wire          _GEN_1911 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h3A;
  wire          compressDataVec_hitReq_29_58;
  assign compressDataVec_hitReq_29_58 = _GEN_1911;
  wire          compressDataVec_hitReq_29_186;
  assign compressDataVec_hitReq_29_186 = _GEN_1911;
  wire          _GEN_1912 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h3A;
  wire          compressDataVec_hitReq_30_58;
  assign compressDataVec_hitReq_30_58 = _GEN_1912;
  wire          compressDataVec_hitReq_30_186;
  assign compressDataVec_hitReq_30_186 = _GEN_1912;
  wire          _GEN_1913 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h3A;
  wire          compressDataVec_hitReq_31_58;
  assign compressDataVec_hitReq_31_58 = _GEN_1913;
  wire          compressDataVec_hitReq_31_186;
  assign compressDataVec_hitReq_31_186 = _GEN_1913;
  wire          compressDataVec_hitReq_32_58 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h3A;
  wire          compressDataVec_hitReq_33_58 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h3A;
  wire          compressDataVec_hitReq_34_58 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h3A;
  wire          compressDataVec_hitReq_35_58 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h3A;
  wire          compressDataVec_hitReq_36_58 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h3A;
  wire          compressDataVec_hitReq_37_58 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h3A;
  wire          compressDataVec_hitReq_38_58 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h3A;
  wire          compressDataVec_hitReq_39_58 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h3A;
  wire          compressDataVec_hitReq_40_58 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h3A;
  wire          compressDataVec_hitReq_41_58 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h3A;
  wire          compressDataVec_hitReq_42_58 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h3A;
  wire          compressDataVec_hitReq_43_58 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h3A;
  wire          compressDataVec_hitReq_44_58 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h3A;
  wire          compressDataVec_hitReq_45_58 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h3A;
  wire          compressDataVec_hitReq_46_58 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h3A;
  wire          compressDataVec_hitReq_47_58 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h3A;
  wire          compressDataVec_hitReq_48_58 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h3A;
  wire          compressDataVec_hitReq_49_58 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h3A;
  wire          compressDataVec_hitReq_50_58 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h3A;
  wire          compressDataVec_hitReq_51_58 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h3A;
  wire          compressDataVec_hitReq_52_58 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h3A;
  wire          compressDataVec_hitReq_53_58 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h3A;
  wire          compressDataVec_hitReq_54_58 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h3A;
  wire          compressDataVec_hitReq_55_58 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h3A;
  wire          compressDataVec_hitReq_56_58 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h3A;
  wire          compressDataVec_hitReq_57_58 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h3A;
  wire          compressDataVec_hitReq_58_58 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h3A;
  wire          compressDataVec_hitReq_59_58 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h3A;
  wire          compressDataVec_hitReq_60_58 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h3A;
  wire          compressDataVec_hitReq_61_58 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h3A;
  wire          compressDataVec_hitReq_62_58 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h3A;
  wire          compressDataVec_hitReq_63_58 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h3A;
  wire [7:0]    compressDataVec_selectReqData_58 =
    (compressDataVec_hitReq_0_58 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_58 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_58 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_58 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_58 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_58 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_58 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_58 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_58 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_58 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_58 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_58 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_58 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_58 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_58 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_58 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_58 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_58 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_58 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_58 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_58 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_58 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_58 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_58 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_58 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_58 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_58 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_58 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_58 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_58 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_58 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_58 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_58 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_58 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_58 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_58 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_58 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_58 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_58 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_58 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_58 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_58 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_58 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_58 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_58 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_58 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_58 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_58 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_58 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_58 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_58 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_58 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_58 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_58 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_58 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_58 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_58 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_58 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_58 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_58 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_58 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_58 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_58 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_58 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_58 = tailCount > 6'h3A;
  wire          _GEN_1914 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h3B;
  wire          compressDataVec_hitReq_0_59;
  assign compressDataVec_hitReq_0_59 = _GEN_1914;
  wire          compressDataVec_hitReq_0_187;
  assign compressDataVec_hitReq_0_187 = _GEN_1914;
  wire          _GEN_1915 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h3B;
  wire          compressDataVec_hitReq_1_59;
  assign compressDataVec_hitReq_1_59 = _GEN_1915;
  wire          compressDataVec_hitReq_1_187;
  assign compressDataVec_hitReq_1_187 = _GEN_1915;
  wire          _GEN_1916 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h3B;
  wire          compressDataVec_hitReq_2_59;
  assign compressDataVec_hitReq_2_59 = _GEN_1916;
  wire          compressDataVec_hitReq_2_187;
  assign compressDataVec_hitReq_2_187 = _GEN_1916;
  wire          _GEN_1917 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h3B;
  wire          compressDataVec_hitReq_3_59;
  assign compressDataVec_hitReq_3_59 = _GEN_1917;
  wire          compressDataVec_hitReq_3_187;
  assign compressDataVec_hitReq_3_187 = _GEN_1917;
  wire          _GEN_1918 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h3B;
  wire          compressDataVec_hitReq_4_59;
  assign compressDataVec_hitReq_4_59 = _GEN_1918;
  wire          compressDataVec_hitReq_4_187;
  assign compressDataVec_hitReq_4_187 = _GEN_1918;
  wire          _GEN_1919 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h3B;
  wire          compressDataVec_hitReq_5_59;
  assign compressDataVec_hitReq_5_59 = _GEN_1919;
  wire          compressDataVec_hitReq_5_187;
  assign compressDataVec_hitReq_5_187 = _GEN_1919;
  wire          _GEN_1920 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h3B;
  wire          compressDataVec_hitReq_6_59;
  assign compressDataVec_hitReq_6_59 = _GEN_1920;
  wire          compressDataVec_hitReq_6_187;
  assign compressDataVec_hitReq_6_187 = _GEN_1920;
  wire          _GEN_1921 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h3B;
  wire          compressDataVec_hitReq_7_59;
  assign compressDataVec_hitReq_7_59 = _GEN_1921;
  wire          compressDataVec_hitReq_7_187;
  assign compressDataVec_hitReq_7_187 = _GEN_1921;
  wire          _GEN_1922 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h3B;
  wire          compressDataVec_hitReq_8_59;
  assign compressDataVec_hitReq_8_59 = _GEN_1922;
  wire          compressDataVec_hitReq_8_187;
  assign compressDataVec_hitReq_8_187 = _GEN_1922;
  wire          _GEN_1923 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h3B;
  wire          compressDataVec_hitReq_9_59;
  assign compressDataVec_hitReq_9_59 = _GEN_1923;
  wire          compressDataVec_hitReq_9_187;
  assign compressDataVec_hitReq_9_187 = _GEN_1923;
  wire          _GEN_1924 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h3B;
  wire          compressDataVec_hitReq_10_59;
  assign compressDataVec_hitReq_10_59 = _GEN_1924;
  wire          compressDataVec_hitReq_10_187;
  assign compressDataVec_hitReq_10_187 = _GEN_1924;
  wire          _GEN_1925 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h3B;
  wire          compressDataVec_hitReq_11_59;
  assign compressDataVec_hitReq_11_59 = _GEN_1925;
  wire          compressDataVec_hitReq_11_187;
  assign compressDataVec_hitReq_11_187 = _GEN_1925;
  wire          _GEN_1926 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h3B;
  wire          compressDataVec_hitReq_12_59;
  assign compressDataVec_hitReq_12_59 = _GEN_1926;
  wire          compressDataVec_hitReq_12_187;
  assign compressDataVec_hitReq_12_187 = _GEN_1926;
  wire          _GEN_1927 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h3B;
  wire          compressDataVec_hitReq_13_59;
  assign compressDataVec_hitReq_13_59 = _GEN_1927;
  wire          compressDataVec_hitReq_13_187;
  assign compressDataVec_hitReq_13_187 = _GEN_1927;
  wire          _GEN_1928 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h3B;
  wire          compressDataVec_hitReq_14_59;
  assign compressDataVec_hitReq_14_59 = _GEN_1928;
  wire          compressDataVec_hitReq_14_187;
  assign compressDataVec_hitReq_14_187 = _GEN_1928;
  wire          _GEN_1929 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h3B;
  wire          compressDataVec_hitReq_15_59;
  assign compressDataVec_hitReq_15_59 = _GEN_1929;
  wire          compressDataVec_hitReq_15_187;
  assign compressDataVec_hitReq_15_187 = _GEN_1929;
  wire          _GEN_1930 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h3B;
  wire          compressDataVec_hitReq_16_59;
  assign compressDataVec_hitReq_16_59 = _GEN_1930;
  wire          compressDataVec_hitReq_16_187;
  assign compressDataVec_hitReq_16_187 = _GEN_1930;
  wire          _GEN_1931 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h3B;
  wire          compressDataVec_hitReq_17_59;
  assign compressDataVec_hitReq_17_59 = _GEN_1931;
  wire          compressDataVec_hitReq_17_187;
  assign compressDataVec_hitReq_17_187 = _GEN_1931;
  wire          _GEN_1932 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h3B;
  wire          compressDataVec_hitReq_18_59;
  assign compressDataVec_hitReq_18_59 = _GEN_1932;
  wire          compressDataVec_hitReq_18_187;
  assign compressDataVec_hitReq_18_187 = _GEN_1932;
  wire          _GEN_1933 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h3B;
  wire          compressDataVec_hitReq_19_59;
  assign compressDataVec_hitReq_19_59 = _GEN_1933;
  wire          compressDataVec_hitReq_19_187;
  assign compressDataVec_hitReq_19_187 = _GEN_1933;
  wire          _GEN_1934 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h3B;
  wire          compressDataVec_hitReq_20_59;
  assign compressDataVec_hitReq_20_59 = _GEN_1934;
  wire          compressDataVec_hitReq_20_187;
  assign compressDataVec_hitReq_20_187 = _GEN_1934;
  wire          _GEN_1935 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h3B;
  wire          compressDataVec_hitReq_21_59;
  assign compressDataVec_hitReq_21_59 = _GEN_1935;
  wire          compressDataVec_hitReq_21_187;
  assign compressDataVec_hitReq_21_187 = _GEN_1935;
  wire          _GEN_1936 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h3B;
  wire          compressDataVec_hitReq_22_59;
  assign compressDataVec_hitReq_22_59 = _GEN_1936;
  wire          compressDataVec_hitReq_22_187;
  assign compressDataVec_hitReq_22_187 = _GEN_1936;
  wire          _GEN_1937 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h3B;
  wire          compressDataVec_hitReq_23_59;
  assign compressDataVec_hitReq_23_59 = _GEN_1937;
  wire          compressDataVec_hitReq_23_187;
  assign compressDataVec_hitReq_23_187 = _GEN_1937;
  wire          _GEN_1938 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h3B;
  wire          compressDataVec_hitReq_24_59;
  assign compressDataVec_hitReq_24_59 = _GEN_1938;
  wire          compressDataVec_hitReq_24_187;
  assign compressDataVec_hitReq_24_187 = _GEN_1938;
  wire          _GEN_1939 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h3B;
  wire          compressDataVec_hitReq_25_59;
  assign compressDataVec_hitReq_25_59 = _GEN_1939;
  wire          compressDataVec_hitReq_25_187;
  assign compressDataVec_hitReq_25_187 = _GEN_1939;
  wire          _GEN_1940 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h3B;
  wire          compressDataVec_hitReq_26_59;
  assign compressDataVec_hitReq_26_59 = _GEN_1940;
  wire          compressDataVec_hitReq_26_187;
  assign compressDataVec_hitReq_26_187 = _GEN_1940;
  wire          _GEN_1941 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h3B;
  wire          compressDataVec_hitReq_27_59;
  assign compressDataVec_hitReq_27_59 = _GEN_1941;
  wire          compressDataVec_hitReq_27_187;
  assign compressDataVec_hitReq_27_187 = _GEN_1941;
  wire          _GEN_1942 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h3B;
  wire          compressDataVec_hitReq_28_59;
  assign compressDataVec_hitReq_28_59 = _GEN_1942;
  wire          compressDataVec_hitReq_28_187;
  assign compressDataVec_hitReq_28_187 = _GEN_1942;
  wire          _GEN_1943 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h3B;
  wire          compressDataVec_hitReq_29_59;
  assign compressDataVec_hitReq_29_59 = _GEN_1943;
  wire          compressDataVec_hitReq_29_187;
  assign compressDataVec_hitReq_29_187 = _GEN_1943;
  wire          _GEN_1944 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h3B;
  wire          compressDataVec_hitReq_30_59;
  assign compressDataVec_hitReq_30_59 = _GEN_1944;
  wire          compressDataVec_hitReq_30_187;
  assign compressDataVec_hitReq_30_187 = _GEN_1944;
  wire          _GEN_1945 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h3B;
  wire          compressDataVec_hitReq_31_59;
  assign compressDataVec_hitReq_31_59 = _GEN_1945;
  wire          compressDataVec_hitReq_31_187;
  assign compressDataVec_hitReq_31_187 = _GEN_1945;
  wire          compressDataVec_hitReq_32_59 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h3B;
  wire          compressDataVec_hitReq_33_59 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h3B;
  wire          compressDataVec_hitReq_34_59 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h3B;
  wire          compressDataVec_hitReq_35_59 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h3B;
  wire          compressDataVec_hitReq_36_59 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h3B;
  wire          compressDataVec_hitReq_37_59 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h3B;
  wire          compressDataVec_hitReq_38_59 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h3B;
  wire          compressDataVec_hitReq_39_59 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h3B;
  wire          compressDataVec_hitReq_40_59 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h3B;
  wire          compressDataVec_hitReq_41_59 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h3B;
  wire          compressDataVec_hitReq_42_59 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h3B;
  wire          compressDataVec_hitReq_43_59 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h3B;
  wire          compressDataVec_hitReq_44_59 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h3B;
  wire          compressDataVec_hitReq_45_59 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h3B;
  wire          compressDataVec_hitReq_46_59 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h3B;
  wire          compressDataVec_hitReq_47_59 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h3B;
  wire          compressDataVec_hitReq_48_59 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h3B;
  wire          compressDataVec_hitReq_49_59 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h3B;
  wire          compressDataVec_hitReq_50_59 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h3B;
  wire          compressDataVec_hitReq_51_59 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h3B;
  wire          compressDataVec_hitReq_52_59 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h3B;
  wire          compressDataVec_hitReq_53_59 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h3B;
  wire          compressDataVec_hitReq_54_59 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h3B;
  wire          compressDataVec_hitReq_55_59 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h3B;
  wire          compressDataVec_hitReq_56_59 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h3B;
  wire          compressDataVec_hitReq_57_59 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h3B;
  wire          compressDataVec_hitReq_58_59 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h3B;
  wire          compressDataVec_hitReq_59_59 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h3B;
  wire          compressDataVec_hitReq_60_59 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h3B;
  wire          compressDataVec_hitReq_61_59 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h3B;
  wire          compressDataVec_hitReq_62_59 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h3B;
  wire          compressDataVec_hitReq_63_59 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h3B;
  wire [7:0]    compressDataVec_selectReqData_59 =
    (compressDataVec_hitReq_0_59 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_59 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_59 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_59 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_59 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_59 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_59 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_59 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_59 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_59 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_59 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_59 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_59 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_59 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_59 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_59 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_59 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_59 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_59 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_59 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_59 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_59 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_59 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_59 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_59 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_59 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_59 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_59 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_59 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_59 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_59 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_59 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_59 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_59 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_59 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_59 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_59 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_59 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_59 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_59 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_59 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_59 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_59 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_59 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_59 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_59 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_59 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_59 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_59 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_59 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_59 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_59 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_59 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_59 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_59 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_59 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_59 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_59 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_59 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_59 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_59 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_59 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_59 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_59 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_59 = tailCount > 6'h3B;
  wire          _GEN_1946 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h3C;
  wire          compressDataVec_hitReq_0_60;
  assign compressDataVec_hitReq_0_60 = _GEN_1946;
  wire          compressDataVec_hitReq_0_188;
  assign compressDataVec_hitReq_0_188 = _GEN_1946;
  wire          _GEN_1947 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h3C;
  wire          compressDataVec_hitReq_1_60;
  assign compressDataVec_hitReq_1_60 = _GEN_1947;
  wire          compressDataVec_hitReq_1_188;
  assign compressDataVec_hitReq_1_188 = _GEN_1947;
  wire          _GEN_1948 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h3C;
  wire          compressDataVec_hitReq_2_60;
  assign compressDataVec_hitReq_2_60 = _GEN_1948;
  wire          compressDataVec_hitReq_2_188;
  assign compressDataVec_hitReq_2_188 = _GEN_1948;
  wire          _GEN_1949 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h3C;
  wire          compressDataVec_hitReq_3_60;
  assign compressDataVec_hitReq_3_60 = _GEN_1949;
  wire          compressDataVec_hitReq_3_188;
  assign compressDataVec_hitReq_3_188 = _GEN_1949;
  wire          _GEN_1950 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h3C;
  wire          compressDataVec_hitReq_4_60;
  assign compressDataVec_hitReq_4_60 = _GEN_1950;
  wire          compressDataVec_hitReq_4_188;
  assign compressDataVec_hitReq_4_188 = _GEN_1950;
  wire          _GEN_1951 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h3C;
  wire          compressDataVec_hitReq_5_60;
  assign compressDataVec_hitReq_5_60 = _GEN_1951;
  wire          compressDataVec_hitReq_5_188;
  assign compressDataVec_hitReq_5_188 = _GEN_1951;
  wire          _GEN_1952 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h3C;
  wire          compressDataVec_hitReq_6_60;
  assign compressDataVec_hitReq_6_60 = _GEN_1952;
  wire          compressDataVec_hitReq_6_188;
  assign compressDataVec_hitReq_6_188 = _GEN_1952;
  wire          _GEN_1953 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h3C;
  wire          compressDataVec_hitReq_7_60;
  assign compressDataVec_hitReq_7_60 = _GEN_1953;
  wire          compressDataVec_hitReq_7_188;
  assign compressDataVec_hitReq_7_188 = _GEN_1953;
  wire          _GEN_1954 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h3C;
  wire          compressDataVec_hitReq_8_60;
  assign compressDataVec_hitReq_8_60 = _GEN_1954;
  wire          compressDataVec_hitReq_8_188;
  assign compressDataVec_hitReq_8_188 = _GEN_1954;
  wire          _GEN_1955 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h3C;
  wire          compressDataVec_hitReq_9_60;
  assign compressDataVec_hitReq_9_60 = _GEN_1955;
  wire          compressDataVec_hitReq_9_188;
  assign compressDataVec_hitReq_9_188 = _GEN_1955;
  wire          _GEN_1956 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h3C;
  wire          compressDataVec_hitReq_10_60;
  assign compressDataVec_hitReq_10_60 = _GEN_1956;
  wire          compressDataVec_hitReq_10_188;
  assign compressDataVec_hitReq_10_188 = _GEN_1956;
  wire          _GEN_1957 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h3C;
  wire          compressDataVec_hitReq_11_60;
  assign compressDataVec_hitReq_11_60 = _GEN_1957;
  wire          compressDataVec_hitReq_11_188;
  assign compressDataVec_hitReq_11_188 = _GEN_1957;
  wire          _GEN_1958 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h3C;
  wire          compressDataVec_hitReq_12_60;
  assign compressDataVec_hitReq_12_60 = _GEN_1958;
  wire          compressDataVec_hitReq_12_188;
  assign compressDataVec_hitReq_12_188 = _GEN_1958;
  wire          _GEN_1959 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h3C;
  wire          compressDataVec_hitReq_13_60;
  assign compressDataVec_hitReq_13_60 = _GEN_1959;
  wire          compressDataVec_hitReq_13_188;
  assign compressDataVec_hitReq_13_188 = _GEN_1959;
  wire          _GEN_1960 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h3C;
  wire          compressDataVec_hitReq_14_60;
  assign compressDataVec_hitReq_14_60 = _GEN_1960;
  wire          compressDataVec_hitReq_14_188;
  assign compressDataVec_hitReq_14_188 = _GEN_1960;
  wire          _GEN_1961 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h3C;
  wire          compressDataVec_hitReq_15_60;
  assign compressDataVec_hitReq_15_60 = _GEN_1961;
  wire          compressDataVec_hitReq_15_188;
  assign compressDataVec_hitReq_15_188 = _GEN_1961;
  wire          _GEN_1962 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h3C;
  wire          compressDataVec_hitReq_16_60;
  assign compressDataVec_hitReq_16_60 = _GEN_1962;
  wire          compressDataVec_hitReq_16_188;
  assign compressDataVec_hitReq_16_188 = _GEN_1962;
  wire          _GEN_1963 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h3C;
  wire          compressDataVec_hitReq_17_60;
  assign compressDataVec_hitReq_17_60 = _GEN_1963;
  wire          compressDataVec_hitReq_17_188;
  assign compressDataVec_hitReq_17_188 = _GEN_1963;
  wire          _GEN_1964 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h3C;
  wire          compressDataVec_hitReq_18_60;
  assign compressDataVec_hitReq_18_60 = _GEN_1964;
  wire          compressDataVec_hitReq_18_188;
  assign compressDataVec_hitReq_18_188 = _GEN_1964;
  wire          _GEN_1965 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h3C;
  wire          compressDataVec_hitReq_19_60;
  assign compressDataVec_hitReq_19_60 = _GEN_1965;
  wire          compressDataVec_hitReq_19_188;
  assign compressDataVec_hitReq_19_188 = _GEN_1965;
  wire          _GEN_1966 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h3C;
  wire          compressDataVec_hitReq_20_60;
  assign compressDataVec_hitReq_20_60 = _GEN_1966;
  wire          compressDataVec_hitReq_20_188;
  assign compressDataVec_hitReq_20_188 = _GEN_1966;
  wire          _GEN_1967 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h3C;
  wire          compressDataVec_hitReq_21_60;
  assign compressDataVec_hitReq_21_60 = _GEN_1967;
  wire          compressDataVec_hitReq_21_188;
  assign compressDataVec_hitReq_21_188 = _GEN_1967;
  wire          _GEN_1968 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h3C;
  wire          compressDataVec_hitReq_22_60;
  assign compressDataVec_hitReq_22_60 = _GEN_1968;
  wire          compressDataVec_hitReq_22_188;
  assign compressDataVec_hitReq_22_188 = _GEN_1968;
  wire          _GEN_1969 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h3C;
  wire          compressDataVec_hitReq_23_60;
  assign compressDataVec_hitReq_23_60 = _GEN_1969;
  wire          compressDataVec_hitReq_23_188;
  assign compressDataVec_hitReq_23_188 = _GEN_1969;
  wire          _GEN_1970 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h3C;
  wire          compressDataVec_hitReq_24_60;
  assign compressDataVec_hitReq_24_60 = _GEN_1970;
  wire          compressDataVec_hitReq_24_188;
  assign compressDataVec_hitReq_24_188 = _GEN_1970;
  wire          _GEN_1971 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h3C;
  wire          compressDataVec_hitReq_25_60;
  assign compressDataVec_hitReq_25_60 = _GEN_1971;
  wire          compressDataVec_hitReq_25_188;
  assign compressDataVec_hitReq_25_188 = _GEN_1971;
  wire          _GEN_1972 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h3C;
  wire          compressDataVec_hitReq_26_60;
  assign compressDataVec_hitReq_26_60 = _GEN_1972;
  wire          compressDataVec_hitReq_26_188;
  assign compressDataVec_hitReq_26_188 = _GEN_1972;
  wire          _GEN_1973 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h3C;
  wire          compressDataVec_hitReq_27_60;
  assign compressDataVec_hitReq_27_60 = _GEN_1973;
  wire          compressDataVec_hitReq_27_188;
  assign compressDataVec_hitReq_27_188 = _GEN_1973;
  wire          _GEN_1974 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h3C;
  wire          compressDataVec_hitReq_28_60;
  assign compressDataVec_hitReq_28_60 = _GEN_1974;
  wire          compressDataVec_hitReq_28_188;
  assign compressDataVec_hitReq_28_188 = _GEN_1974;
  wire          _GEN_1975 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h3C;
  wire          compressDataVec_hitReq_29_60;
  assign compressDataVec_hitReq_29_60 = _GEN_1975;
  wire          compressDataVec_hitReq_29_188;
  assign compressDataVec_hitReq_29_188 = _GEN_1975;
  wire          _GEN_1976 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h3C;
  wire          compressDataVec_hitReq_30_60;
  assign compressDataVec_hitReq_30_60 = _GEN_1976;
  wire          compressDataVec_hitReq_30_188;
  assign compressDataVec_hitReq_30_188 = _GEN_1976;
  wire          _GEN_1977 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h3C;
  wire          compressDataVec_hitReq_31_60;
  assign compressDataVec_hitReq_31_60 = _GEN_1977;
  wire          compressDataVec_hitReq_31_188;
  assign compressDataVec_hitReq_31_188 = _GEN_1977;
  wire          compressDataVec_hitReq_32_60 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h3C;
  wire          compressDataVec_hitReq_33_60 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h3C;
  wire          compressDataVec_hitReq_34_60 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h3C;
  wire          compressDataVec_hitReq_35_60 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h3C;
  wire          compressDataVec_hitReq_36_60 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h3C;
  wire          compressDataVec_hitReq_37_60 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h3C;
  wire          compressDataVec_hitReq_38_60 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h3C;
  wire          compressDataVec_hitReq_39_60 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h3C;
  wire          compressDataVec_hitReq_40_60 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h3C;
  wire          compressDataVec_hitReq_41_60 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h3C;
  wire          compressDataVec_hitReq_42_60 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h3C;
  wire          compressDataVec_hitReq_43_60 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h3C;
  wire          compressDataVec_hitReq_44_60 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h3C;
  wire          compressDataVec_hitReq_45_60 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h3C;
  wire          compressDataVec_hitReq_46_60 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h3C;
  wire          compressDataVec_hitReq_47_60 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h3C;
  wire          compressDataVec_hitReq_48_60 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h3C;
  wire          compressDataVec_hitReq_49_60 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h3C;
  wire          compressDataVec_hitReq_50_60 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h3C;
  wire          compressDataVec_hitReq_51_60 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h3C;
  wire          compressDataVec_hitReq_52_60 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h3C;
  wire          compressDataVec_hitReq_53_60 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h3C;
  wire          compressDataVec_hitReq_54_60 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h3C;
  wire          compressDataVec_hitReq_55_60 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h3C;
  wire          compressDataVec_hitReq_56_60 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h3C;
  wire          compressDataVec_hitReq_57_60 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h3C;
  wire          compressDataVec_hitReq_58_60 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h3C;
  wire          compressDataVec_hitReq_59_60 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h3C;
  wire          compressDataVec_hitReq_60_60 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h3C;
  wire          compressDataVec_hitReq_61_60 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h3C;
  wire          compressDataVec_hitReq_62_60 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h3C;
  wire          compressDataVec_hitReq_63_60 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h3C;
  wire [7:0]    compressDataVec_selectReqData_60 =
    (compressDataVec_hitReq_0_60 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_60 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_60 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_60 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_60 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_60 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_60 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_60 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_60 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_60 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_60 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_60 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_60 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_60 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_60 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_60 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_60 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_60 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_60 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_60 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_60 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_60 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_60 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_60 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_60 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_60 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_60 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_60 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_60 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_60 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_60 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_60 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_60 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_60 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_60 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_60 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_60 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_60 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_60 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_60 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_60 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_60 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_60 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_60 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_60 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_60 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_60 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_60 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_60 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_60 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_60 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_60 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_60 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_60 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_60 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_60 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_60 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_60 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_60 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_60 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_60 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_60 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_60 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_60 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_60 = tailCount > 6'h3C;
  wire          _GEN_1978 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h3D;
  wire          compressDataVec_hitReq_0_61;
  assign compressDataVec_hitReq_0_61 = _GEN_1978;
  wire          compressDataVec_hitReq_0_189;
  assign compressDataVec_hitReq_0_189 = _GEN_1978;
  wire          _GEN_1979 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h3D;
  wire          compressDataVec_hitReq_1_61;
  assign compressDataVec_hitReq_1_61 = _GEN_1979;
  wire          compressDataVec_hitReq_1_189;
  assign compressDataVec_hitReq_1_189 = _GEN_1979;
  wire          _GEN_1980 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h3D;
  wire          compressDataVec_hitReq_2_61;
  assign compressDataVec_hitReq_2_61 = _GEN_1980;
  wire          compressDataVec_hitReq_2_189;
  assign compressDataVec_hitReq_2_189 = _GEN_1980;
  wire          _GEN_1981 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h3D;
  wire          compressDataVec_hitReq_3_61;
  assign compressDataVec_hitReq_3_61 = _GEN_1981;
  wire          compressDataVec_hitReq_3_189;
  assign compressDataVec_hitReq_3_189 = _GEN_1981;
  wire          _GEN_1982 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h3D;
  wire          compressDataVec_hitReq_4_61;
  assign compressDataVec_hitReq_4_61 = _GEN_1982;
  wire          compressDataVec_hitReq_4_189;
  assign compressDataVec_hitReq_4_189 = _GEN_1982;
  wire          _GEN_1983 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h3D;
  wire          compressDataVec_hitReq_5_61;
  assign compressDataVec_hitReq_5_61 = _GEN_1983;
  wire          compressDataVec_hitReq_5_189;
  assign compressDataVec_hitReq_5_189 = _GEN_1983;
  wire          _GEN_1984 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h3D;
  wire          compressDataVec_hitReq_6_61;
  assign compressDataVec_hitReq_6_61 = _GEN_1984;
  wire          compressDataVec_hitReq_6_189;
  assign compressDataVec_hitReq_6_189 = _GEN_1984;
  wire          _GEN_1985 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h3D;
  wire          compressDataVec_hitReq_7_61;
  assign compressDataVec_hitReq_7_61 = _GEN_1985;
  wire          compressDataVec_hitReq_7_189;
  assign compressDataVec_hitReq_7_189 = _GEN_1985;
  wire          _GEN_1986 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h3D;
  wire          compressDataVec_hitReq_8_61;
  assign compressDataVec_hitReq_8_61 = _GEN_1986;
  wire          compressDataVec_hitReq_8_189;
  assign compressDataVec_hitReq_8_189 = _GEN_1986;
  wire          _GEN_1987 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h3D;
  wire          compressDataVec_hitReq_9_61;
  assign compressDataVec_hitReq_9_61 = _GEN_1987;
  wire          compressDataVec_hitReq_9_189;
  assign compressDataVec_hitReq_9_189 = _GEN_1987;
  wire          _GEN_1988 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h3D;
  wire          compressDataVec_hitReq_10_61;
  assign compressDataVec_hitReq_10_61 = _GEN_1988;
  wire          compressDataVec_hitReq_10_189;
  assign compressDataVec_hitReq_10_189 = _GEN_1988;
  wire          _GEN_1989 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h3D;
  wire          compressDataVec_hitReq_11_61;
  assign compressDataVec_hitReq_11_61 = _GEN_1989;
  wire          compressDataVec_hitReq_11_189;
  assign compressDataVec_hitReq_11_189 = _GEN_1989;
  wire          _GEN_1990 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h3D;
  wire          compressDataVec_hitReq_12_61;
  assign compressDataVec_hitReq_12_61 = _GEN_1990;
  wire          compressDataVec_hitReq_12_189;
  assign compressDataVec_hitReq_12_189 = _GEN_1990;
  wire          _GEN_1991 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h3D;
  wire          compressDataVec_hitReq_13_61;
  assign compressDataVec_hitReq_13_61 = _GEN_1991;
  wire          compressDataVec_hitReq_13_189;
  assign compressDataVec_hitReq_13_189 = _GEN_1991;
  wire          _GEN_1992 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h3D;
  wire          compressDataVec_hitReq_14_61;
  assign compressDataVec_hitReq_14_61 = _GEN_1992;
  wire          compressDataVec_hitReq_14_189;
  assign compressDataVec_hitReq_14_189 = _GEN_1992;
  wire          _GEN_1993 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h3D;
  wire          compressDataVec_hitReq_15_61;
  assign compressDataVec_hitReq_15_61 = _GEN_1993;
  wire          compressDataVec_hitReq_15_189;
  assign compressDataVec_hitReq_15_189 = _GEN_1993;
  wire          _GEN_1994 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h3D;
  wire          compressDataVec_hitReq_16_61;
  assign compressDataVec_hitReq_16_61 = _GEN_1994;
  wire          compressDataVec_hitReq_16_189;
  assign compressDataVec_hitReq_16_189 = _GEN_1994;
  wire          _GEN_1995 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h3D;
  wire          compressDataVec_hitReq_17_61;
  assign compressDataVec_hitReq_17_61 = _GEN_1995;
  wire          compressDataVec_hitReq_17_189;
  assign compressDataVec_hitReq_17_189 = _GEN_1995;
  wire          _GEN_1996 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h3D;
  wire          compressDataVec_hitReq_18_61;
  assign compressDataVec_hitReq_18_61 = _GEN_1996;
  wire          compressDataVec_hitReq_18_189;
  assign compressDataVec_hitReq_18_189 = _GEN_1996;
  wire          _GEN_1997 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h3D;
  wire          compressDataVec_hitReq_19_61;
  assign compressDataVec_hitReq_19_61 = _GEN_1997;
  wire          compressDataVec_hitReq_19_189;
  assign compressDataVec_hitReq_19_189 = _GEN_1997;
  wire          _GEN_1998 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h3D;
  wire          compressDataVec_hitReq_20_61;
  assign compressDataVec_hitReq_20_61 = _GEN_1998;
  wire          compressDataVec_hitReq_20_189;
  assign compressDataVec_hitReq_20_189 = _GEN_1998;
  wire          _GEN_1999 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h3D;
  wire          compressDataVec_hitReq_21_61;
  assign compressDataVec_hitReq_21_61 = _GEN_1999;
  wire          compressDataVec_hitReq_21_189;
  assign compressDataVec_hitReq_21_189 = _GEN_1999;
  wire          _GEN_2000 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h3D;
  wire          compressDataVec_hitReq_22_61;
  assign compressDataVec_hitReq_22_61 = _GEN_2000;
  wire          compressDataVec_hitReq_22_189;
  assign compressDataVec_hitReq_22_189 = _GEN_2000;
  wire          _GEN_2001 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h3D;
  wire          compressDataVec_hitReq_23_61;
  assign compressDataVec_hitReq_23_61 = _GEN_2001;
  wire          compressDataVec_hitReq_23_189;
  assign compressDataVec_hitReq_23_189 = _GEN_2001;
  wire          _GEN_2002 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h3D;
  wire          compressDataVec_hitReq_24_61;
  assign compressDataVec_hitReq_24_61 = _GEN_2002;
  wire          compressDataVec_hitReq_24_189;
  assign compressDataVec_hitReq_24_189 = _GEN_2002;
  wire          _GEN_2003 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h3D;
  wire          compressDataVec_hitReq_25_61;
  assign compressDataVec_hitReq_25_61 = _GEN_2003;
  wire          compressDataVec_hitReq_25_189;
  assign compressDataVec_hitReq_25_189 = _GEN_2003;
  wire          _GEN_2004 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h3D;
  wire          compressDataVec_hitReq_26_61;
  assign compressDataVec_hitReq_26_61 = _GEN_2004;
  wire          compressDataVec_hitReq_26_189;
  assign compressDataVec_hitReq_26_189 = _GEN_2004;
  wire          _GEN_2005 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h3D;
  wire          compressDataVec_hitReq_27_61;
  assign compressDataVec_hitReq_27_61 = _GEN_2005;
  wire          compressDataVec_hitReq_27_189;
  assign compressDataVec_hitReq_27_189 = _GEN_2005;
  wire          _GEN_2006 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h3D;
  wire          compressDataVec_hitReq_28_61;
  assign compressDataVec_hitReq_28_61 = _GEN_2006;
  wire          compressDataVec_hitReq_28_189;
  assign compressDataVec_hitReq_28_189 = _GEN_2006;
  wire          _GEN_2007 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h3D;
  wire          compressDataVec_hitReq_29_61;
  assign compressDataVec_hitReq_29_61 = _GEN_2007;
  wire          compressDataVec_hitReq_29_189;
  assign compressDataVec_hitReq_29_189 = _GEN_2007;
  wire          _GEN_2008 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h3D;
  wire          compressDataVec_hitReq_30_61;
  assign compressDataVec_hitReq_30_61 = _GEN_2008;
  wire          compressDataVec_hitReq_30_189;
  assign compressDataVec_hitReq_30_189 = _GEN_2008;
  wire          _GEN_2009 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h3D;
  wire          compressDataVec_hitReq_31_61;
  assign compressDataVec_hitReq_31_61 = _GEN_2009;
  wire          compressDataVec_hitReq_31_189;
  assign compressDataVec_hitReq_31_189 = _GEN_2009;
  wire          compressDataVec_hitReq_32_61 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h3D;
  wire          compressDataVec_hitReq_33_61 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h3D;
  wire          compressDataVec_hitReq_34_61 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h3D;
  wire          compressDataVec_hitReq_35_61 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h3D;
  wire          compressDataVec_hitReq_36_61 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h3D;
  wire          compressDataVec_hitReq_37_61 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h3D;
  wire          compressDataVec_hitReq_38_61 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h3D;
  wire          compressDataVec_hitReq_39_61 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h3D;
  wire          compressDataVec_hitReq_40_61 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h3D;
  wire          compressDataVec_hitReq_41_61 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h3D;
  wire          compressDataVec_hitReq_42_61 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h3D;
  wire          compressDataVec_hitReq_43_61 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h3D;
  wire          compressDataVec_hitReq_44_61 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h3D;
  wire          compressDataVec_hitReq_45_61 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h3D;
  wire          compressDataVec_hitReq_46_61 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h3D;
  wire          compressDataVec_hitReq_47_61 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h3D;
  wire          compressDataVec_hitReq_48_61 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h3D;
  wire          compressDataVec_hitReq_49_61 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h3D;
  wire          compressDataVec_hitReq_50_61 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h3D;
  wire          compressDataVec_hitReq_51_61 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h3D;
  wire          compressDataVec_hitReq_52_61 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h3D;
  wire          compressDataVec_hitReq_53_61 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h3D;
  wire          compressDataVec_hitReq_54_61 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h3D;
  wire          compressDataVec_hitReq_55_61 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h3D;
  wire          compressDataVec_hitReq_56_61 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h3D;
  wire          compressDataVec_hitReq_57_61 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h3D;
  wire          compressDataVec_hitReq_58_61 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h3D;
  wire          compressDataVec_hitReq_59_61 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h3D;
  wire          compressDataVec_hitReq_60_61 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h3D;
  wire          compressDataVec_hitReq_61_61 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h3D;
  wire          compressDataVec_hitReq_62_61 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h3D;
  wire          compressDataVec_hitReq_63_61 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h3D;
  wire [7:0]    compressDataVec_selectReqData_61 =
    (compressDataVec_hitReq_0_61 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_61 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_61 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_61 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_61 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_61 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_61 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_61 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_61 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_61 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_61 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_61 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_61 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_61 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_61 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_61 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_61 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_61 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_61 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_61 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_61 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_61 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_61 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_61 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_61 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_61 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_61 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_61 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_61 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_61 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_61 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_61 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_61 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_61 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_61 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_61 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_61 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_61 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_61 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_61 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_61 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_61 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_61 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_61 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_61 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_61 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_61 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_61 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_61 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_61 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_61 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_61 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_61 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_61 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_61 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_61 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_61 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_61 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_61 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_61 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_61 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_61 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_61 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_61 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_61 = tailCount > 6'h3D;
  wire          _GEN_2010 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h3E;
  wire          compressDataVec_hitReq_0_62;
  assign compressDataVec_hitReq_0_62 = _GEN_2010;
  wire          compressDataVec_hitReq_0_190;
  assign compressDataVec_hitReq_0_190 = _GEN_2010;
  wire          _GEN_2011 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h3E;
  wire          compressDataVec_hitReq_1_62;
  assign compressDataVec_hitReq_1_62 = _GEN_2011;
  wire          compressDataVec_hitReq_1_190;
  assign compressDataVec_hitReq_1_190 = _GEN_2011;
  wire          _GEN_2012 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h3E;
  wire          compressDataVec_hitReq_2_62;
  assign compressDataVec_hitReq_2_62 = _GEN_2012;
  wire          compressDataVec_hitReq_2_190;
  assign compressDataVec_hitReq_2_190 = _GEN_2012;
  wire          _GEN_2013 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h3E;
  wire          compressDataVec_hitReq_3_62;
  assign compressDataVec_hitReq_3_62 = _GEN_2013;
  wire          compressDataVec_hitReq_3_190;
  assign compressDataVec_hitReq_3_190 = _GEN_2013;
  wire          _GEN_2014 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h3E;
  wire          compressDataVec_hitReq_4_62;
  assign compressDataVec_hitReq_4_62 = _GEN_2014;
  wire          compressDataVec_hitReq_4_190;
  assign compressDataVec_hitReq_4_190 = _GEN_2014;
  wire          _GEN_2015 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h3E;
  wire          compressDataVec_hitReq_5_62;
  assign compressDataVec_hitReq_5_62 = _GEN_2015;
  wire          compressDataVec_hitReq_5_190;
  assign compressDataVec_hitReq_5_190 = _GEN_2015;
  wire          _GEN_2016 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h3E;
  wire          compressDataVec_hitReq_6_62;
  assign compressDataVec_hitReq_6_62 = _GEN_2016;
  wire          compressDataVec_hitReq_6_190;
  assign compressDataVec_hitReq_6_190 = _GEN_2016;
  wire          _GEN_2017 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h3E;
  wire          compressDataVec_hitReq_7_62;
  assign compressDataVec_hitReq_7_62 = _GEN_2017;
  wire          compressDataVec_hitReq_7_190;
  assign compressDataVec_hitReq_7_190 = _GEN_2017;
  wire          _GEN_2018 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h3E;
  wire          compressDataVec_hitReq_8_62;
  assign compressDataVec_hitReq_8_62 = _GEN_2018;
  wire          compressDataVec_hitReq_8_190;
  assign compressDataVec_hitReq_8_190 = _GEN_2018;
  wire          _GEN_2019 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h3E;
  wire          compressDataVec_hitReq_9_62;
  assign compressDataVec_hitReq_9_62 = _GEN_2019;
  wire          compressDataVec_hitReq_9_190;
  assign compressDataVec_hitReq_9_190 = _GEN_2019;
  wire          _GEN_2020 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h3E;
  wire          compressDataVec_hitReq_10_62;
  assign compressDataVec_hitReq_10_62 = _GEN_2020;
  wire          compressDataVec_hitReq_10_190;
  assign compressDataVec_hitReq_10_190 = _GEN_2020;
  wire          _GEN_2021 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h3E;
  wire          compressDataVec_hitReq_11_62;
  assign compressDataVec_hitReq_11_62 = _GEN_2021;
  wire          compressDataVec_hitReq_11_190;
  assign compressDataVec_hitReq_11_190 = _GEN_2021;
  wire          _GEN_2022 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h3E;
  wire          compressDataVec_hitReq_12_62;
  assign compressDataVec_hitReq_12_62 = _GEN_2022;
  wire          compressDataVec_hitReq_12_190;
  assign compressDataVec_hitReq_12_190 = _GEN_2022;
  wire          _GEN_2023 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h3E;
  wire          compressDataVec_hitReq_13_62;
  assign compressDataVec_hitReq_13_62 = _GEN_2023;
  wire          compressDataVec_hitReq_13_190;
  assign compressDataVec_hitReq_13_190 = _GEN_2023;
  wire          _GEN_2024 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h3E;
  wire          compressDataVec_hitReq_14_62;
  assign compressDataVec_hitReq_14_62 = _GEN_2024;
  wire          compressDataVec_hitReq_14_190;
  assign compressDataVec_hitReq_14_190 = _GEN_2024;
  wire          _GEN_2025 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h3E;
  wire          compressDataVec_hitReq_15_62;
  assign compressDataVec_hitReq_15_62 = _GEN_2025;
  wire          compressDataVec_hitReq_15_190;
  assign compressDataVec_hitReq_15_190 = _GEN_2025;
  wire          _GEN_2026 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h3E;
  wire          compressDataVec_hitReq_16_62;
  assign compressDataVec_hitReq_16_62 = _GEN_2026;
  wire          compressDataVec_hitReq_16_190;
  assign compressDataVec_hitReq_16_190 = _GEN_2026;
  wire          _GEN_2027 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h3E;
  wire          compressDataVec_hitReq_17_62;
  assign compressDataVec_hitReq_17_62 = _GEN_2027;
  wire          compressDataVec_hitReq_17_190;
  assign compressDataVec_hitReq_17_190 = _GEN_2027;
  wire          _GEN_2028 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h3E;
  wire          compressDataVec_hitReq_18_62;
  assign compressDataVec_hitReq_18_62 = _GEN_2028;
  wire          compressDataVec_hitReq_18_190;
  assign compressDataVec_hitReq_18_190 = _GEN_2028;
  wire          _GEN_2029 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h3E;
  wire          compressDataVec_hitReq_19_62;
  assign compressDataVec_hitReq_19_62 = _GEN_2029;
  wire          compressDataVec_hitReq_19_190;
  assign compressDataVec_hitReq_19_190 = _GEN_2029;
  wire          _GEN_2030 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h3E;
  wire          compressDataVec_hitReq_20_62;
  assign compressDataVec_hitReq_20_62 = _GEN_2030;
  wire          compressDataVec_hitReq_20_190;
  assign compressDataVec_hitReq_20_190 = _GEN_2030;
  wire          _GEN_2031 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h3E;
  wire          compressDataVec_hitReq_21_62;
  assign compressDataVec_hitReq_21_62 = _GEN_2031;
  wire          compressDataVec_hitReq_21_190;
  assign compressDataVec_hitReq_21_190 = _GEN_2031;
  wire          _GEN_2032 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h3E;
  wire          compressDataVec_hitReq_22_62;
  assign compressDataVec_hitReq_22_62 = _GEN_2032;
  wire          compressDataVec_hitReq_22_190;
  assign compressDataVec_hitReq_22_190 = _GEN_2032;
  wire          _GEN_2033 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h3E;
  wire          compressDataVec_hitReq_23_62;
  assign compressDataVec_hitReq_23_62 = _GEN_2033;
  wire          compressDataVec_hitReq_23_190;
  assign compressDataVec_hitReq_23_190 = _GEN_2033;
  wire          _GEN_2034 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h3E;
  wire          compressDataVec_hitReq_24_62;
  assign compressDataVec_hitReq_24_62 = _GEN_2034;
  wire          compressDataVec_hitReq_24_190;
  assign compressDataVec_hitReq_24_190 = _GEN_2034;
  wire          _GEN_2035 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h3E;
  wire          compressDataVec_hitReq_25_62;
  assign compressDataVec_hitReq_25_62 = _GEN_2035;
  wire          compressDataVec_hitReq_25_190;
  assign compressDataVec_hitReq_25_190 = _GEN_2035;
  wire          _GEN_2036 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h3E;
  wire          compressDataVec_hitReq_26_62;
  assign compressDataVec_hitReq_26_62 = _GEN_2036;
  wire          compressDataVec_hitReq_26_190;
  assign compressDataVec_hitReq_26_190 = _GEN_2036;
  wire          _GEN_2037 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h3E;
  wire          compressDataVec_hitReq_27_62;
  assign compressDataVec_hitReq_27_62 = _GEN_2037;
  wire          compressDataVec_hitReq_27_190;
  assign compressDataVec_hitReq_27_190 = _GEN_2037;
  wire          _GEN_2038 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h3E;
  wire          compressDataVec_hitReq_28_62;
  assign compressDataVec_hitReq_28_62 = _GEN_2038;
  wire          compressDataVec_hitReq_28_190;
  assign compressDataVec_hitReq_28_190 = _GEN_2038;
  wire          _GEN_2039 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h3E;
  wire          compressDataVec_hitReq_29_62;
  assign compressDataVec_hitReq_29_62 = _GEN_2039;
  wire          compressDataVec_hitReq_29_190;
  assign compressDataVec_hitReq_29_190 = _GEN_2039;
  wire          _GEN_2040 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h3E;
  wire          compressDataVec_hitReq_30_62;
  assign compressDataVec_hitReq_30_62 = _GEN_2040;
  wire          compressDataVec_hitReq_30_190;
  assign compressDataVec_hitReq_30_190 = _GEN_2040;
  wire          _GEN_2041 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h3E;
  wire          compressDataVec_hitReq_31_62;
  assign compressDataVec_hitReq_31_62 = _GEN_2041;
  wire          compressDataVec_hitReq_31_190;
  assign compressDataVec_hitReq_31_190 = _GEN_2041;
  wire          compressDataVec_hitReq_32_62 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h3E;
  wire          compressDataVec_hitReq_33_62 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h3E;
  wire          compressDataVec_hitReq_34_62 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h3E;
  wire          compressDataVec_hitReq_35_62 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h3E;
  wire          compressDataVec_hitReq_36_62 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h3E;
  wire          compressDataVec_hitReq_37_62 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h3E;
  wire          compressDataVec_hitReq_38_62 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h3E;
  wire          compressDataVec_hitReq_39_62 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h3E;
  wire          compressDataVec_hitReq_40_62 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h3E;
  wire          compressDataVec_hitReq_41_62 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h3E;
  wire          compressDataVec_hitReq_42_62 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h3E;
  wire          compressDataVec_hitReq_43_62 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h3E;
  wire          compressDataVec_hitReq_44_62 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h3E;
  wire          compressDataVec_hitReq_45_62 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h3E;
  wire          compressDataVec_hitReq_46_62 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h3E;
  wire          compressDataVec_hitReq_47_62 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h3E;
  wire          compressDataVec_hitReq_48_62 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h3E;
  wire          compressDataVec_hitReq_49_62 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h3E;
  wire          compressDataVec_hitReq_50_62 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h3E;
  wire          compressDataVec_hitReq_51_62 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h3E;
  wire          compressDataVec_hitReq_52_62 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h3E;
  wire          compressDataVec_hitReq_53_62 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h3E;
  wire          compressDataVec_hitReq_54_62 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h3E;
  wire          compressDataVec_hitReq_55_62 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h3E;
  wire          compressDataVec_hitReq_56_62 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h3E;
  wire          compressDataVec_hitReq_57_62 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h3E;
  wire          compressDataVec_hitReq_58_62 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h3E;
  wire          compressDataVec_hitReq_59_62 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h3E;
  wire          compressDataVec_hitReq_60_62 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h3E;
  wire          compressDataVec_hitReq_61_62 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h3E;
  wire          compressDataVec_hitReq_62_62 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h3E;
  wire          compressDataVec_hitReq_63_62 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h3E;
  wire [7:0]    compressDataVec_selectReqData_62 =
    (compressDataVec_hitReq_0_62 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_62 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_62 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_62 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_62 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_62 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_62 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_62 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_62 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_62 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_62 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_62 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_62 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_62 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_62 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_62 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_62 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_62 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_62 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_62 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_62 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_62 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_62 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_62 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_62 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_62 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_62 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_62 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_62 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_62 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_62 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_62 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_62 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_62 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_62 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_62 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_62 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_62 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_62 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_62 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_62 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_62 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_62 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_62 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_62 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_62 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_62 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_62 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_62 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_62 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_62 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_62 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_62 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_62 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_62 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_62 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_62 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_62 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_62 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_62 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_62 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_62 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_62 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_62 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_useTail_62 = &tailCount;
  wire          _GEN_2042 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h3F;
  wire          compressDataVec_hitReq_0_63;
  assign compressDataVec_hitReq_0_63 = _GEN_2042;
  wire          compressDataVec_hitReq_0_191;
  assign compressDataVec_hitReq_0_191 = _GEN_2042;
  wire          _GEN_2043 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h3F;
  wire          compressDataVec_hitReq_1_63;
  assign compressDataVec_hitReq_1_63 = _GEN_2043;
  wire          compressDataVec_hitReq_1_191;
  assign compressDataVec_hitReq_1_191 = _GEN_2043;
  wire          _GEN_2044 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h3F;
  wire          compressDataVec_hitReq_2_63;
  assign compressDataVec_hitReq_2_63 = _GEN_2044;
  wire          compressDataVec_hitReq_2_191;
  assign compressDataVec_hitReq_2_191 = _GEN_2044;
  wire          _GEN_2045 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h3F;
  wire          compressDataVec_hitReq_3_63;
  assign compressDataVec_hitReq_3_63 = _GEN_2045;
  wire          compressDataVec_hitReq_3_191;
  assign compressDataVec_hitReq_3_191 = _GEN_2045;
  wire          _GEN_2046 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h3F;
  wire          compressDataVec_hitReq_4_63;
  assign compressDataVec_hitReq_4_63 = _GEN_2046;
  wire          compressDataVec_hitReq_4_191;
  assign compressDataVec_hitReq_4_191 = _GEN_2046;
  wire          _GEN_2047 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h3F;
  wire          compressDataVec_hitReq_5_63;
  assign compressDataVec_hitReq_5_63 = _GEN_2047;
  wire          compressDataVec_hitReq_5_191;
  assign compressDataVec_hitReq_5_191 = _GEN_2047;
  wire          _GEN_2048 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h3F;
  wire          compressDataVec_hitReq_6_63;
  assign compressDataVec_hitReq_6_63 = _GEN_2048;
  wire          compressDataVec_hitReq_6_191;
  assign compressDataVec_hitReq_6_191 = _GEN_2048;
  wire          _GEN_2049 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h3F;
  wire          compressDataVec_hitReq_7_63;
  assign compressDataVec_hitReq_7_63 = _GEN_2049;
  wire          compressDataVec_hitReq_7_191;
  assign compressDataVec_hitReq_7_191 = _GEN_2049;
  wire          _GEN_2050 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h3F;
  wire          compressDataVec_hitReq_8_63;
  assign compressDataVec_hitReq_8_63 = _GEN_2050;
  wire          compressDataVec_hitReq_8_191;
  assign compressDataVec_hitReq_8_191 = _GEN_2050;
  wire          _GEN_2051 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h3F;
  wire          compressDataVec_hitReq_9_63;
  assign compressDataVec_hitReq_9_63 = _GEN_2051;
  wire          compressDataVec_hitReq_9_191;
  assign compressDataVec_hitReq_9_191 = _GEN_2051;
  wire          _GEN_2052 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h3F;
  wire          compressDataVec_hitReq_10_63;
  assign compressDataVec_hitReq_10_63 = _GEN_2052;
  wire          compressDataVec_hitReq_10_191;
  assign compressDataVec_hitReq_10_191 = _GEN_2052;
  wire          _GEN_2053 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h3F;
  wire          compressDataVec_hitReq_11_63;
  assign compressDataVec_hitReq_11_63 = _GEN_2053;
  wire          compressDataVec_hitReq_11_191;
  assign compressDataVec_hitReq_11_191 = _GEN_2053;
  wire          _GEN_2054 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h3F;
  wire          compressDataVec_hitReq_12_63;
  assign compressDataVec_hitReq_12_63 = _GEN_2054;
  wire          compressDataVec_hitReq_12_191;
  assign compressDataVec_hitReq_12_191 = _GEN_2054;
  wire          _GEN_2055 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h3F;
  wire          compressDataVec_hitReq_13_63;
  assign compressDataVec_hitReq_13_63 = _GEN_2055;
  wire          compressDataVec_hitReq_13_191;
  assign compressDataVec_hitReq_13_191 = _GEN_2055;
  wire          _GEN_2056 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h3F;
  wire          compressDataVec_hitReq_14_63;
  assign compressDataVec_hitReq_14_63 = _GEN_2056;
  wire          compressDataVec_hitReq_14_191;
  assign compressDataVec_hitReq_14_191 = _GEN_2056;
  wire          _GEN_2057 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h3F;
  wire          compressDataVec_hitReq_15_63;
  assign compressDataVec_hitReq_15_63 = _GEN_2057;
  wire          compressDataVec_hitReq_15_191;
  assign compressDataVec_hitReq_15_191 = _GEN_2057;
  wire          _GEN_2058 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h3F;
  wire          compressDataVec_hitReq_16_63;
  assign compressDataVec_hitReq_16_63 = _GEN_2058;
  wire          compressDataVec_hitReq_16_191;
  assign compressDataVec_hitReq_16_191 = _GEN_2058;
  wire          _GEN_2059 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h3F;
  wire          compressDataVec_hitReq_17_63;
  assign compressDataVec_hitReq_17_63 = _GEN_2059;
  wire          compressDataVec_hitReq_17_191;
  assign compressDataVec_hitReq_17_191 = _GEN_2059;
  wire          _GEN_2060 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h3F;
  wire          compressDataVec_hitReq_18_63;
  assign compressDataVec_hitReq_18_63 = _GEN_2060;
  wire          compressDataVec_hitReq_18_191;
  assign compressDataVec_hitReq_18_191 = _GEN_2060;
  wire          _GEN_2061 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h3F;
  wire          compressDataVec_hitReq_19_63;
  assign compressDataVec_hitReq_19_63 = _GEN_2061;
  wire          compressDataVec_hitReq_19_191;
  assign compressDataVec_hitReq_19_191 = _GEN_2061;
  wire          _GEN_2062 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h3F;
  wire          compressDataVec_hitReq_20_63;
  assign compressDataVec_hitReq_20_63 = _GEN_2062;
  wire          compressDataVec_hitReq_20_191;
  assign compressDataVec_hitReq_20_191 = _GEN_2062;
  wire          _GEN_2063 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h3F;
  wire          compressDataVec_hitReq_21_63;
  assign compressDataVec_hitReq_21_63 = _GEN_2063;
  wire          compressDataVec_hitReq_21_191;
  assign compressDataVec_hitReq_21_191 = _GEN_2063;
  wire          _GEN_2064 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h3F;
  wire          compressDataVec_hitReq_22_63;
  assign compressDataVec_hitReq_22_63 = _GEN_2064;
  wire          compressDataVec_hitReq_22_191;
  assign compressDataVec_hitReq_22_191 = _GEN_2064;
  wire          _GEN_2065 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h3F;
  wire          compressDataVec_hitReq_23_63;
  assign compressDataVec_hitReq_23_63 = _GEN_2065;
  wire          compressDataVec_hitReq_23_191;
  assign compressDataVec_hitReq_23_191 = _GEN_2065;
  wire          _GEN_2066 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h3F;
  wire          compressDataVec_hitReq_24_63;
  assign compressDataVec_hitReq_24_63 = _GEN_2066;
  wire          compressDataVec_hitReq_24_191;
  assign compressDataVec_hitReq_24_191 = _GEN_2066;
  wire          _GEN_2067 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h3F;
  wire          compressDataVec_hitReq_25_63;
  assign compressDataVec_hitReq_25_63 = _GEN_2067;
  wire          compressDataVec_hitReq_25_191;
  assign compressDataVec_hitReq_25_191 = _GEN_2067;
  wire          _GEN_2068 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h3F;
  wire          compressDataVec_hitReq_26_63;
  assign compressDataVec_hitReq_26_63 = _GEN_2068;
  wire          compressDataVec_hitReq_26_191;
  assign compressDataVec_hitReq_26_191 = _GEN_2068;
  wire          _GEN_2069 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h3F;
  wire          compressDataVec_hitReq_27_63;
  assign compressDataVec_hitReq_27_63 = _GEN_2069;
  wire          compressDataVec_hitReq_27_191;
  assign compressDataVec_hitReq_27_191 = _GEN_2069;
  wire          _GEN_2070 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h3F;
  wire          compressDataVec_hitReq_28_63;
  assign compressDataVec_hitReq_28_63 = _GEN_2070;
  wire          compressDataVec_hitReq_28_191;
  assign compressDataVec_hitReq_28_191 = _GEN_2070;
  wire          _GEN_2071 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h3F;
  wire          compressDataVec_hitReq_29_63;
  assign compressDataVec_hitReq_29_63 = _GEN_2071;
  wire          compressDataVec_hitReq_29_191;
  assign compressDataVec_hitReq_29_191 = _GEN_2071;
  wire          _GEN_2072 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h3F;
  wire          compressDataVec_hitReq_30_63;
  assign compressDataVec_hitReq_30_63 = _GEN_2072;
  wire          compressDataVec_hitReq_30_191;
  assign compressDataVec_hitReq_30_191 = _GEN_2072;
  wire          _GEN_2073 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h3F;
  wire          compressDataVec_hitReq_31_63;
  assign compressDataVec_hitReq_31_63 = _GEN_2073;
  wire          compressDataVec_hitReq_31_191;
  assign compressDataVec_hitReq_31_191 = _GEN_2073;
  wire          compressDataVec_hitReq_32_63 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h3F;
  wire          compressDataVec_hitReq_33_63 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h3F;
  wire          compressDataVec_hitReq_34_63 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h3F;
  wire          compressDataVec_hitReq_35_63 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h3F;
  wire          compressDataVec_hitReq_36_63 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h3F;
  wire          compressDataVec_hitReq_37_63 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h3F;
  wire          compressDataVec_hitReq_38_63 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h3F;
  wire          compressDataVec_hitReq_39_63 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h3F;
  wire          compressDataVec_hitReq_40_63 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h3F;
  wire          compressDataVec_hitReq_41_63 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h3F;
  wire          compressDataVec_hitReq_42_63 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h3F;
  wire          compressDataVec_hitReq_43_63 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h3F;
  wire          compressDataVec_hitReq_44_63 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h3F;
  wire          compressDataVec_hitReq_45_63 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h3F;
  wire          compressDataVec_hitReq_46_63 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h3F;
  wire          compressDataVec_hitReq_47_63 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h3F;
  wire          compressDataVec_hitReq_48_63 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h3F;
  wire          compressDataVec_hitReq_49_63 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h3F;
  wire          compressDataVec_hitReq_50_63 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h3F;
  wire          compressDataVec_hitReq_51_63 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h3F;
  wire          compressDataVec_hitReq_52_63 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h3F;
  wire          compressDataVec_hitReq_53_63 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h3F;
  wire          compressDataVec_hitReq_54_63 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h3F;
  wire          compressDataVec_hitReq_55_63 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h3F;
  wire          compressDataVec_hitReq_56_63 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h3F;
  wire          compressDataVec_hitReq_57_63 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h3F;
  wire          compressDataVec_hitReq_58_63 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h3F;
  wire          compressDataVec_hitReq_59_63 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h3F;
  wire          compressDataVec_hitReq_60_63 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h3F;
  wire          compressDataVec_hitReq_61_63 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h3F;
  wire          compressDataVec_hitReq_62_63 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h3F;
  wire          compressDataVec_hitReq_63_63 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h3F;
  wire [7:0]    compressDataVec_selectReqData_63 =
    (compressDataVec_hitReq_0_63 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_63 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_63 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_63 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_63 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_63 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_63 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_63 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_63 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_63 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_63 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_63 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_63 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_63 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_63 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_63 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_63 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_63 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_63 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_63 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_63 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_63 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_63 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_63 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_63 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_63 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_63 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_63 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_63 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_63 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_63 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_63 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_63 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_63 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_63 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_63 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_63 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_63 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_63 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_63 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_63 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_63 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_63 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_63 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_63 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_63 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_63 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_63 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_63 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_63 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_63 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_63 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_63 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_63 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_63 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_63 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_63 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_63 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_63 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_63 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_63 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_63 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_63 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_63 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_64 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h40;
  wire          compressDataVec_hitReq_1_64 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h40;
  wire          compressDataVec_hitReq_2_64 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h40;
  wire          compressDataVec_hitReq_3_64 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h40;
  wire          compressDataVec_hitReq_4_64 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h40;
  wire          compressDataVec_hitReq_5_64 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h40;
  wire          compressDataVec_hitReq_6_64 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h40;
  wire          compressDataVec_hitReq_7_64 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h40;
  wire          compressDataVec_hitReq_8_64 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h40;
  wire          compressDataVec_hitReq_9_64 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h40;
  wire          compressDataVec_hitReq_10_64 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h40;
  wire          compressDataVec_hitReq_11_64 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h40;
  wire          compressDataVec_hitReq_12_64 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h40;
  wire          compressDataVec_hitReq_13_64 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h40;
  wire          compressDataVec_hitReq_14_64 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h40;
  wire          compressDataVec_hitReq_15_64 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h40;
  wire          compressDataVec_hitReq_16_64 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h40;
  wire          compressDataVec_hitReq_17_64 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h40;
  wire          compressDataVec_hitReq_18_64 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h40;
  wire          compressDataVec_hitReq_19_64 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h40;
  wire          compressDataVec_hitReq_20_64 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h40;
  wire          compressDataVec_hitReq_21_64 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h40;
  wire          compressDataVec_hitReq_22_64 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h40;
  wire          compressDataVec_hitReq_23_64 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h40;
  wire          compressDataVec_hitReq_24_64 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h40;
  wire          compressDataVec_hitReq_25_64 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h40;
  wire          compressDataVec_hitReq_26_64 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h40;
  wire          compressDataVec_hitReq_27_64 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h40;
  wire          compressDataVec_hitReq_28_64 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h40;
  wire          compressDataVec_hitReq_29_64 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h40;
  wire          compressDataVec_hitReq_30_64 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h40;
  wire          compressDataVec_hitReq_31_64 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h40;
  wire          compressDataVec_hitReq_32_64 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h40;
  wire          compressDataVec_hitReq_33_64 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h40;
  wire          compressDataVec_hitReq_34_64 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h40;
  wire          compressDataVec_hitReq_35_64 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h40;
  wire          compressDataVec_hitReq_36_64 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h40;
  wire          compressDataVec_hitReq_37_64 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h40;
  wire          compressDataVec_hitReq_38_64 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h40;
  wire          compressDataVec_hitReq_39_64 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h40;
  wire          compressDataVec_hitReq_40_64 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h40;
  wire          compressDataVec_hitReq_41_64 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h40;
  wire          compressDataVec_hitReq_42_64 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h40;
  wire          compressDataVec_hitReq_43_64 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h40;
  wire          compressDataVec_hitReq_44_64 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h40;
  wire          compressDataVec_hitReq_45_64 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h40;
  wire          compressDataVec_hitReq_46_64 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h40;
  wire          compressDataVec_hitReq_47_64 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h40;
  wire          compressDataVec_hitReq_48_64 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h40;
  wire          compressDataVec_hitReq_49_64 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h40;
  wire          compressDataVec_hitReq_50_64 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h40;
  wire          compressDataVec_hitReq_51_64 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h40;
  wire          compressDataVec_hitReq_52_64 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h40;
  wire          compressDataVec_hitReq_53_64 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h40;
  wire          compressDataVec_hitReq_54_64 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h40;
  wire          compressDataVec_hitReq_55_64 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h40;
  wire          compressDataVec_hitReq_56_64 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h40;
  wire          compressDataVec_hitReq_57_64 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h40;
  wire          compressDataVec_hitReq_58_64 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h40;
  wire          compressDataVec_hitReq_59_64 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h40;
  wire          compressDataVec_hitReq_60_64 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h40;
  wire          compressDataVec_hitReq_61_64 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h40;
  wire          compressDataVec_hitReq_62_64 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h40;
  wire          compressDataVec_hitReq_63_64 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h40;
  wire [7:0]    compressDataVec_selectReqData_64 =
    (compressDataVec_hitReq_0_64 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_64 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_64 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_64 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_64 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_64 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_64 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_64 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_64 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_64 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_64 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_64 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_64 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_64 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_64 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_64 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_64 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_64 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_64 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_64 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_64 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_64 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_64 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_64 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_64 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_64 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_64 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_64 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_64 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_64 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_64 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_64 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_64 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_64 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_64 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_64 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_64 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_64 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_64 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_64 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_64 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_64 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_64 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_64 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_64 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_64 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_64 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_64 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_64 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_64 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_64 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_64 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_64 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_64 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_64 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_64 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_64 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_64 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_64 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_64 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_64 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_64 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_64 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_64 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_65 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h41;
  wire          compressDataVec_hitReq_1_65 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h41;
  wire          compressDataVec_hitReq_2_65 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h41;
  wire          compressDataVec_hitReq_3_65 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h41;
  wire          compressDataVec_hitReq_4_65 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h41;
  wire          compressDataVec_hitReq_5_65 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h41;
  wire          compressDataVec_hitReq_6_65 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h41;
  wire          compressDataVec_hitReq_7_65 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h41;
  wire          compressDataVec_hitReq_8_65 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h41;
  wire          compressDataVec_hitReq_9_65 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h41;
  wire          compressDataVec_hitReq_10_65 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h41;
  wire          compressDataVec_hitReq_11_65 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h41;
  wire          compressDataVec_hitReq_12_65 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h41;
  wire          compressDataVec_hitReq_13_65 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h41;
  wire          compressDataVec_hitReq_14_65 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h41;
  wire          compressDataVec_hitReq_15_65 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h41;
  wire          compressDataVec_hitReq_16_65 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h41;
  wire          compressDataVec_hitReq_17_65 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h41;
  wire          compressDataVec_hitReq_18_65 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h41;
  wire          compressDataVec_hitReq_19_65 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h41;
  wire          compressDataVec_hitReq_20_65 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h41;
  wire          compressDataVec_hitReq_21_65 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h41;
  wire          compressDataVec_hitReq_22_65 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h41;
  wire          compressDataVec_hitReq_23_65 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h41;
  wire          compressDataVec_hitReq_24_65 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h41;
  wire          compressDataVec_hitReq_25_65 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h41;
  wire          compressDataVec_hitReq_26_65 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h41;
  wire          compressDataVec_hitReq_27_65 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h41;
  wire          compressDataVec_hitReq_28_65 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h41;
  wire          compressDataVec_hitReq_29_65 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h41;
  wire          compressDataVec_hitReq_30_65 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h41;
  wire          compressDataVec_hitReq_31_65 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h41;
  wire          compressDataVec_hitReq_32_65 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h41;
  wire          compressDataVec_hitReq_33_65 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h41;
  wire          compressDataVec_hitReq_34_65 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h41;
  wire          compressDataVec_hitReq_35_65 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h41;
  wire          compressDataVec_hitReq_36_65 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h41;
  wire          compressDataVec_hitReq_37_65 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h41;
  wire          compressDataVec_hitReq_38_65 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h41;
  wire          compressDataVec_hitReq_39_65 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h41;
  wire          compressDataVec_hitReq_40_65 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h41;
  wire          compressDataVec_hitReq_41_65 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h41;
  wire          compressDataVec_hitReq_42_65 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h41;
  wire          compressDataVec_hitReq_43_65 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h41;
  wire          compressDataVec_hitReq_44_65 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h41;
  wire          compressDataVec_hitReq_45_65 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h41;
  wire          compressDataVec_hitReq_46_65 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h41;
  wire          compressDataVec_hitReq_47_65 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h41;
  wire          compressDataVec_hitReq_48_65 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h41;
  wire          compressDataVec_hitReq_49_65 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h41;
  wire          compressDataVec_hitReq_50_65 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h41;
  wire          compressDataVec_hitReq_51_65 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h41;
  wire          compressDataVec_hitReq_52_65 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h41;
  wire          compressDataVec_hitReq_53_65 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h41;
  wire          compressDataVec_hitReq_54_65 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h41;
  wire          compressDataVec_hitReq_55_65 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h41;
  wire          compressDataVec_hitReq_56_65 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h41;
  wire          compressDataVec_hitReq_57_65 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h41;
  wire          compressDataVec_hitReq_58_65 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h41;
  wire          compressDataVec_hitReq_59_65 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h41;
  wire          compressDataVec_hitReq_60_65 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h41;
  wire          compressDataVec_hitReq_61_65 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h41;
  wire          compressDataVec_hitReq_62_65 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h41;
  wire          compressDataVec_hitReq_63_65 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h41;
  wire [7:0]    compressDataVec_selectReqData_65 =
    (compressDataVec_hitReq_0_65 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_65 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_65 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_65 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_65 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_65 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_65 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_65 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_65 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_65 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_65 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_65 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_65 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_65 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_65 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_65 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_65 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_65 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_65 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_65 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_65 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_65 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_65 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_65 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_65 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_65 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_65 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_65 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_65 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_65 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_65 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_65 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_65 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_65 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_65 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_65 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_65 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_65 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_65 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_65 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_65 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_65 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_65 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_65 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_65 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_65 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_65 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_65 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_65 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_65 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_65 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_65 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_65 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_65 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_65 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_65 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_65 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_65 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_65 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_65 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_65 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_65 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_65 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_65 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_66 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h42;
  wire          compressDataVec_hitReq_1_66 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h42;
  wire          compressDataVec_hitReq_2_66 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h42;
  wire          compressDataVec_hitReq_3_66 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h42;
  wire          compressDataVec_hitReq_4_66 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h42;
  wire          compressDataVec_hitReq_5_66 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h42;
  wire          compressDataVec_hitReq_6_66 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h42;
  wire          compressDataVec_hitReq_7_66 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h42;
  wire          compressDataVec_hitReq_8_66 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h42;
  wire          compressDataVec_hitReq_9_66 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h42;
  wire          compressDataVec_hitReq_10_66 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h42;
  wire          compressDataVec_hitReq_11_66 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h42;
  wire          compressDataVec_hitReq_12_66 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h42;
  wire          compressDataVec_hitReq_13_66 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h42;
  wire          compressDataVec_hitReq_14_66 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h42;
  wire          compressDataVec_hitReq_15_66 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h42;
  wire          compressDataVec_hitReq_16_66 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h42;
  wire          compressDataVec_hitReq_17_66 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h42;
  wire          compressDataVec_hitReq_18_66 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h42;
  wire          compressDataVec_hitReq_19_66 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h42;
  wire          compressDataVec_hitReq_20_66 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h42;
  wire          compressDataVec_hitReq_21_66 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h42;
  wire          compressDataVec_hitReq_22_66 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h42;
  wire          compressDataVec_hitReq_23_66 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h42;
  wire          compressDataVec_hitReq_24_66 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h42;
  wire          compressDataVec_hitReq_25_66 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h42;
  wire          compressDataVec_hitReq_26_66 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h42;
  wire          compressDataVec_hitReq_27_66 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h42;
  wire          compressDataVec_hitReq_28_66 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h42;
  wire          compressDataVec_hitReq_29_66 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h42;
  wire          compressDataVec_hitReq_30_66 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h42;
  wire          compressDataVec_hitReq_31_66 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h42;
  wire          compressDataVec_hitReq_32_66 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h42;
  wire          compressDataVec_hitReq_33_66 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h42;
  wire          compressDataVec_hitReq_34_66 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h42;
  wire          compressDataVec_hitReq_35_66 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h42;
  wire          compressDataVec_hitReq_36_66 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h42;
  wire          compressDataVec_hitReq_37_66 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h42;
  wire          compressDataVec_hitReq_38_66 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h42;
  wire          compressDataVec_hitReq_39_66 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h42;
  wire          compressDataVec_hitReq_40_66 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h42;
  wire          compressDataVec_hitReq_41_66 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h42;
  wire          compressDataVec_hitReq_42_66 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h42;
  wire          compressDataVec_hitReq_43_66 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h42;
  wire          compressDataVec_hitReq_44_66 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h42;
  wire          compressDataVec_hitReq_45_66 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h42;
  wire          compressDataVec_hitReq_46_66 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h42;
  wire          compressDataVec_hitReq_47_66 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h42;
  wire          compressDataVec_hitReq_48_66 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h42;
  wire          compressDataVec_hitReq_49_66 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h42;
  wire          compressDataVec_hitReq_50_66 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h42;
  wire          compressDataVec_hitReq_51_66 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h42;
  wire          compressDataVec_hitReq_52_66 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h42;
  wire          compressDataVec_hitReq_53_66 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h42;
  wire          compressDataVec_hitReq_54_66 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h42;
  wire          compressDataVec_hitReq_55_66 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h42;
  wire          compressDataVec_hitReq_56_66 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h42;
  wire          compressDataVec_hitReq_57_66 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h42;
  wire          compressDataVec_hitReq_58_66 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h42;
  wire          compressDataVec_hitReq_59_66 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h42;
  wire          compressDataVec_hitReq_60_66 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h42;
  wire          compressDataVec_hitReq_61_66 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h42;
  wire          compressDataVec_hitReq_62_66 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h42;
  wire          compressDataVec_hitReq_63_66 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h42;
  wire [7:0]    compressDataVec_selectReqData_66 =
    (compressDataVec_hitReq_0_66 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_66 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_66 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_66 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_66 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_66 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_66 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_66 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_66 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_66 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_66 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_66 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_66 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_66 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_66 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_66 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_66 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_66 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_66 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_66 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_66 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_66 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_66 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_66 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_66 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_66 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_66 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_66 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_66 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_66 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_66 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_66 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_66 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_66 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_66 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_66 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_66 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_66 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_66 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_66 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_66 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_66 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_66 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_66 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_66 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_66 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_66 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_66 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_66 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_66 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_66 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_66 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_66 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_66 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_66 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_66 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_66 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_66 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_66 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_66 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_66 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_66 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_66 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_66 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_67 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h43;
  wire          compressDataVec_hitReq_1_67 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h43;
  wire          compressDataVec_hitReq_2_67 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h43;
  wire          compressDataVec_hitReq_3_67 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h43;
  wire          compressDataVec_hitReq_4_67 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h43;
  wire          compressDataVec_hitReq_5_67 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h43;
  wire          compressDataVec_hitReq_6_67 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h43;
  wire          compressDataVec_hitReq_7_67 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h43;
  wire          compressDataVec_hitReq_8_67 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h43;
  wire          compressDataVec_hitReq_9_67 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h43;
  wire          compressDataVec_hitReq_10_67 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h43;
  wire          compressDataVec_hitReq_11_67 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h43;
  wire          compressDataVec_hitReq_12_67 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h43;
  wire          compressDataVec_hitReq_13_67 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h43;
  wire          compressDataVec_hitReq_14_67 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h43;
  wire          compressDataVec_hitReq_15_67 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h43;
  wire          compressDataVec_hitReq_16_67 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h43;
  wire          compressDataVec_hitReq_17_67 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h43;
  wire          compressDataVec_hitReq_18_67 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h43;
  wire          compressDataVec_hitReq_19_67 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h43;
  wire          compressDataVec_hitReq_20_67 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h43;
  wire          compressDataVec_hitReq_21_67 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h43;
  wire          compressDataVec_hitReq_22_67 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h43;
  wire          compressDataVec_hitReq_23_67 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h43;
  wire          compressDataVec_hitReq_24_67 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h43;
  wire          compressDataVec_hitReq_25_67 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h43;
  wire          compressDataVec_hitReq_26_67 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h43;
  wire          compressDataVec_hitReq_27_67 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h43;
  wire          compressDataVec_hitReq_28_67 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h43;
  wire          compressDataVec_hitReq_29_67 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h43;
  wire          compressDataVec_hitReq_30_67 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h43;
  wire          compressDataVec_hitReq_31_67 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h43;
  wire          compressDataVec_hitReq_32_67 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h43;
  wire          compressDataVec_hitReq_33_67 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h43;
  wire          compressDataVec_hitReq_34_67 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h43;
  wire          compressDataVec_hitReq_35_67 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h43;
  wire          compressDataVec_hitReq_36_67 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h43;
  wire          compressDataVec_hitReq_37_67 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h43;
  wire          compressDataVec_hitReq_38_67 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h43;
  wire          compressDataVec_hitReq_39_67 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h43;
  wire          compressDataVec_hitReq_40_67 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h43;
  wire          compressDataVec_hitReq_41_67 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h43;
  wire          compressDataVec_hitReq_42_67 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h43;
  wire          compressDataVec_hitReq_43_67 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h43;
  wire          compressDataVec_hitReq_44_67 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h43;
  wire          compressDataVec_hitReq_45_67 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h43;
  wire          compressDataVec_hitReq_46_67 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h43;
  wire          compressDataVec_hitReq_47_67 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h43;
  wire          compressDataVec_hitReq_48_67 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h43;
  wire          compressDataVec_hitReq_49_67 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h43;
  wire          compressDataVec_hitReq_50_67 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h43;
  wire          compressDataVec_hitReq_51_67 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h43;
  wire          compressDataVec_hitReq_52_67 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h43;
  wire          compressDataVec_hitReq_53_67 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h43;
  wire          compressDataVec_hitReq_54_67 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h43;
  wire          compressDataVec_hitReq_55_67 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h43;
  wire          compressDataVec_hitReq_56_67 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h43;
  wire          compressDataVec_hitReq_57_67 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h43;
  wire          compressDataVec_hitReq_58_67 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h43;
  wire          compressDataVec_hitReq_59_67 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h43;
  wire          compressDataVec_hitReq_60_67 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h43;
  wire          compressDataVec_hitReq_61_67 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h43;
  wire          compressDataVec_hitReq_62_67 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h43;
  wire          compressDataVec_hitReq_63_67 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h43;
  wire [7:0]    compressDataVec_selectReqData_67 =
    (compressDataVec_hitReq_0_67 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_67 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_67 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_67 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_67 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_67 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_67 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_67 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_67 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_67 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_67 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_67 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_67 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_67 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_67 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_67 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_67 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_67 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_67 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_67 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_67 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_67 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_67 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_67 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_67 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_67 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_67 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_67 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_67 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_67 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_67 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_67 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_67 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_67 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_67 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_67 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_67 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_67 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_67 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_67 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_67 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_67 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_67 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_67 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_67 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_67 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_67 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_67 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_67 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_67 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_67 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_67 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_67 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_67 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_67 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_67 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_67 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_67 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_67 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_67 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_67 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_67 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_67 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_67 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_68 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h44;
  wire          compressDataVec_hitReq_1_68 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h44;
  wire          compressDataVec_hitReq_2_68 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h44;
  wire          compressDataVec_hitReq_3_68 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h44;
  wire          compressDataVec_hitReq_4_68 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h44;
  wire          compressDataVec_hitReq_5_68 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h44;
  wire          compressDataVec_hitReq_6_68 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h44;
  wire          compressDataVec_hitReq_7_68 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h44;
  wire          compressDataVec_hitReq_8_68 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h44;
  wire          compressDataVec_hitReq_9_68 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h44;
  wire          compressDataVec_hitReq_10_68 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h44;
  wire          compressDataVec_hitReq_11_68 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h44;
  wire          compressDataVec_hitReq_12_68 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h44;
  wire          compressDataVec_hitReq_13_68 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h44;
  wire          compressDataVec_hitReq_14_68 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h44;
  wire          compressDataVec_hitReq_15_68 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h44;
  wire          compressDataVec_hitReq_16_68 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h44;
  wire          compressDataVec_hitReq_17_68 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h44;
  wire          compressDataVec_hitReq_18_68 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h44;
  wire          compressDataVec_hitReq_19_68 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h44;
  wire          compressDataVec_hitReq_20_68 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h44;
  wire          compressDataVec_hitReq_21_68 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h44;
  wire          compressDataVec_hitReq_22_68 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h44;
  wire          compressDataVec_hitReq_23_68 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h44;
  wire          compressDataVec_hitReq_24_68 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h44;
  wire          compressDataVec_hitReq_25_68 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h44;
  wire          compressDataVec_hitReq_26_68 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h44;
  wire          compressDataVec_hitReq_27_68 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h44;
  wire          compressDataVec_hitReq_28_68 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h44;
  wire          compressDataVec_hitReq_29_68 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h44;
  wire          compressDataVec_hitReq_30_68 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h44;
  wire          compressDataVec_hitReq_31_68 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h44;
  wire          compressDataVec_hitReq_32_68 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h44;
  wire          compressDataVec_hitReq_33_68 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h44;
  wire          compressDataVec_hitReq_34_68 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h44;
  wire          compressDataVec_hitReq_35_68 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h44;
  wire          compressDataVec_hitReq_36_68 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h44;
  wire          compressDataVec_hitReq_37_68 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h44;
  wire          compressDataVec_hitReq_38_68 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h44;
  wire          compressDataVec_hitReq_39_68 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h44;
  wire          compressDataVec_hitReq_40_68 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h44;
  wire          compressDataVec_hitReq_41_68 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h44;
  wire          compressDataVec_hitReq_42_68 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h44;
  wire          compressDataVec_hitReq_43_68 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h44;
  wire          compressDataVec_hitReq_44_68 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h44;
  wire          compressDataVec_hitReq_45_68 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h44;
  wire          compressDataVec_hitReq_46_68 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h44;
  wire          compressDataVec_hitReq_47_68 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h44;
  wire          compressDataVec_hitReq_48_68 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h44;
  wire          compressDataVec_hitReq_49_68 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h44;
  wire          compressDataVec_hitReq_50_68 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h44;
  wire          compressDataVec_hitReq_51_68 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h44;
  wire          compressDataVec_hitReq_52_68 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h44;
  wire          compressDataVec_hitReq_53_68 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h44;
  wire          compressDataVec_hitReq_54_68 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h44;
  wire          compressDataVec_hitReq_55_68 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h44;
  wire          compressDataVec_hitReq_56_68 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h44;
  wire          compressDataVec_hitReq_57_68 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h44;
  wire          compressDataVec_hitReq_58_68 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h44;
  wire          compressDataVec_hitReq_59_68 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h44;
  wire          compressDataVec_hitReq_60_68 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h44;
  wire          compressDataVec_hitReq_61_68 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h44;
  wire          compressDataVec_hitReq_62_68 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h44;
  wire          compressDataVec_hitReq_63_68 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h44;
  wire [7:0]    compressDataVec_selectReqData_68 =
    (compressDataVec_hitReq_0_68 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_68 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_68 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_68 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_68 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_68 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_68 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_68 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_68 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_68 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_68 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_68 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_68 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_68 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_68 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_68 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_68 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_68 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_68 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_68 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_68 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_68 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_68 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_68 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_68 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_68 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_68 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_68 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_68 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_68 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_68 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_68 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_68 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_68 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_68 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_68 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_68 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_68 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_68 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_68 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_68 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_68 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_68 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_68 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_68 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_68 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_68 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_68 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_68 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_68 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_68 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_68 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_68 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_68 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_68 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_68 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_68 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_68 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_68 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_68 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_68 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_68 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_68 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_68 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_69 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h45;
  wire          compressDataVec_hitReq_1_69 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h45;
  wire          compressDataVec_hitReq_2_69 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h45;
  wire          compressDataVec_hitReq_3_69 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h45;
  wire          compressDataVec_hitReq_4_69 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h45;
  wire          compressDataVec_hitReq_5_69 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h45;
  wire          compressDataVec_hitReq_6_69 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h45;
  wire          compressDataVec_hitReq_7_69 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h45;
  wire          compressDataVec_hitReq_8_69 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h45;
  wire          compressDataVec_hitReq_9_69 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h45;
  wire          compressDataVec_hitReq_10_69 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h45;
  wire          compressDataVec_hitReq_11_69 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h45;
  wire          compressDataVec_hitReq_12_69 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h45;
  wire          compressDataVec_hitReq_13_69 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h45;
  wire          compressDataVec_hitReq_14_69 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h45;
  wire          compressDataVec_hitReq_15_69 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h45;
  wire          compressDataVec_hitReq_16_69 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h45;
  wire          compressDataVec_hitReq_17_69 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h45;
  wire          compressDataVec_hitReq_18_69 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h45;
  wire          compressDataVec_hitReq_19_69 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h45;
  wire          compressDataVec_hitReq_20_69 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h45;
  wire          compressDataVec_hitReq_21_69 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h45;
  wire          compressDataVec_hitReq_22_69 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h45;
  wire          compressDataVec_hitReq_23_69 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h45;
  wire          compressDataVec_hitReq_24_69 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h45;
  wire          compressDataVec_hitReq_25_69 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h45;
  wire          compressDataVec_hitReq_26_69 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h45;
  wire          compressDataVec_hitReq_27_69 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h45;
  wire          compressDataVec_hitReq_28_69 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h45;
  wire          compressDataVec_hitReq_29_69 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h45;
  wire          compressDataVec_hitReq_30_69 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h45;
  wire          compressDataVec_hitReq_31_69 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h45;
  wire          compressDataVec_hitReq_32_69 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h45;
  wire          compressDataVec_hitReq_33_69 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h45;
  wire          compressDataVec_hitReq_34_69 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h45;
  wire          compressDataVec_hitReq_35_69 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h45;
  wire          compressDataVec_hitReq_36_69 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h45;
  wire          compressDataVec_hitReq_37_69 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h45;
  wire          compressDataVec_hitReq_38_69 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h45;
  wire          compressDataVec_hitReq_39_69 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h45;
  wire          compressDataVec_hitReq_40_69 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h45;
  wire          compressDataVec_hitReq_41_69 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h45;
  wire          compressDataVec_hitReq_42_69 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h45;
  wire          compressDataVec_hitReq_43_69 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h45;
  wire          compressDataVec_hitReq_44_69 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h45;
  wire          compressDataVec_hitReq_45_69 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h45;
  wire          compressDataVec_hitReq_46_69 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h45;
  wire          compressDataVec_hitReq_47_69 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h45;
  wire          compressDataVec_hitReq_48_69 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h45;
  wire          compressDataVec_hitReq_49_69 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h45;
  wire          compressDataVec_hitReq_50_69 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h45;
  wire          compressDataVec_hitReq_51_69 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h45;
  wire          compressDataVec_hitReq_52_69 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h45;
  wire          compressDataVec_hitReq_53_69 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h45;
  wire          compressDataVec_hitReq_54_69 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h45;
  wire          compressDataVec_hitReq_55_69 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h45;
  wire          compressDataVec_hitReq_56_69 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h45;
  wire          compressDataVec_hitReq_57_69 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h45;
  wire          compressDataVec_hitReq_58_69 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h45;
  wire          compressDataVec_hitReq_59_69 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h45;
  wire          compressDataVec_hitReq_60_69 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h45;
  wire          compressDataVec_hitReq_61_69 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h45;
  wire          compressDataVec_hitReq_62_69 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h45;
  wire          compressDataVec_hitReq_63_69 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h45;
  wire [7:0]    compressDataVec_selectReqData_69 =
    (compressDataVec_hitReq_0_69 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_69 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_69 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_69 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_69 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_69 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_69 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_69 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_69 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_69 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_69 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_69 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_69 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_69 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_69 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_69 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_69 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_69 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_69 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_69 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_69 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_69 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_69 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_69 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_69 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_69 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_69 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_69 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_69 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_69 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_69 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_69 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_69 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_69 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_69 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_69 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_69 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_69 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_69 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_69 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_69 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_69 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_69 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_69 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_69 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_69 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_69 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_69 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_69 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_69 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_69 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_69 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_69 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_69 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_69 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_69 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_69 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_69 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_69 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_69 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_69 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_69 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_69 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_69 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_70 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h46;
  wire          compressDataVec_hitReq_1_70 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h46;
  wire          compressDataVec_hitReq_2_70 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h46;
  wire          compressDataVec_hitReq_3_70 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h46;
  wire          compressDataVec_hitReq_4_70 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h46;
  wire          compressDataVec_hitReq_5_70 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h46;
  wire          compressDataVec_hitReq_6_70 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h46;
  wire          compressDataVec_hitReq_7_70 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h46;
  wire          compressDataVec_hitReq_8_70 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h46;
  wire          compressDataVec_hitReq_9_70 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h46;
  wire          compressDataVec_hitReq_10_70 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h46;
  wire          compressDataVec_hitReq_11_70 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h46;
  wire          compressDataVec_hitReq_12_70 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h46;
  wire          compressDataVec_hitReq_13_70 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h46;
  wire          compressDataVec_hitReq_14_70 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h46;
  wire          compressDataVec_hitReq_15_70 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h46;
  wire          compressDataVec_hitReq_16_70 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h46;
  wire          compressDataVec_hitReq_17_70 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h46;
  wire          compressDataVec_hitReq_18_70 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h46;
  wire          compressDataVec_hitReq_19_70 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h46;
  wire          compressDataVec_hitReq_20_70 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h46;
  wire          compressDataVec_hitReq_21_70 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h46;
  wire          compressDataVec_hitReq_22_70 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h46;
  wire          compressDataVec_hitReq_23_70 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h46;
  wire          compressDataVec_hitReq_24_70 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h46;
  wire          compressDataVec_hitReq_25_70 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h46;
  wire          compressDataVec_hitReq_26_70 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h46;
  wire          compressDataVec_hitReq_27_70 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h46;
  wire          compressDataVec_hitReq_28_70 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h46;
  wire          compressDataVec_hitReq_29_70 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h46;
  wire          compressDataVec_hitReq_30_70 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h46;
  wire          compressDataVec_hitReq_31_70 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h46;
  wire          compressDataVec_hitReq_32_70 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h46;
  wire          compressDataVec_hitReq_33_70 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h46;
  wire          compressDataVec_hitReq_34_70 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h46;
  wire          compressDataVec_hitReq_35_70 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h46;
  wire          compressDataVec_hitReq_36_70 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h46;
  wire          compressDataVec_hitReq_37_70 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h46;
  wire          compressDataVec_hitReq_38_70 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h46;
  wire          compressDataVec_hitReq_39_70 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h46;
  wire          compressDataVec_hitReq_40_70 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h46;
  wire          compressDataVec_hitReq_41_70 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h46;
  wire          compressDataVec_hitReq_42_70 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h46;
  wire          compressDataVec_hitReq_43_70 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h46;
  wire          compressDataVec_hitReq_44_70 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h46;
  wire          compressDataVec_hitReq_45_70 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h46;
  wire          compressDataVec_hitReq_46_70 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h46;
  wire          compressDataVec_hitReq_47_70 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h46;
  wire          compressDataVec_hitReq_48_70 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h46;
  wire          compressDataVec_hitReq_49_70 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h46;
  wire          compressDataVec_hitReq_50_70 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h46;
  wire          compressDataVec_hitReq_51_70 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h46;
  wire          compressDataVec_hitReq_52_70 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h46;
  wire          compressDataVec_hitReq_53_70 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h46;
  wire          compressDataVec_hitReq_54_70 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h46;
  wire          compressDataVec_hitReq_55_70 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h46;
  wire          compressDataVec_hitReq_56_70 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h46;
  wire          compressDataVec_hitReq_57_70 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h46;
  wire          compressDataVec_hitReq_58_70 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h46;
  wire          compressDataVec_hitReq_59_70 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h46;
  wire          compressDataVec_hitReq_60_70 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h46;
  wire          compressDataVec_hitReq_61_70 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h46;
  wire          compressDataVec_hitReq_62_70 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h46;
  wire          compressDataVec_hitReq_63_70 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h46;
  wire [7:0]    compressDataVec_selectReqData_70 =
    (compressDataVec_hitReq_0_70 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_70 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_70 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_70 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_70 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_70 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_70 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_70 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_70 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_70 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_70 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_70 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_70 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_70 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_70 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_70 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_70 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_70 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_70 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_70 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_70 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_70 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_70 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_70 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_70 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_70 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_70 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_70 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_70 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_70 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_70 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_70 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_70 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_70 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_70 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_70 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_70 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_70 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_70 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_70 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_70 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_70 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_70 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_70 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_70 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_70 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_70 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_70 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_70 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_70 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_70 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_70 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_70 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_70 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_70 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_70 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_70 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_70 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_70 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_70 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_70 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_70 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_70 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_70 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_71 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h47;
  wire          compressDataVec_hitReq_1_71 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h47;
  wire          compressDataVec_hitReq_2_71 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h47;
  wire          compressDataVec_hitReq_3_71 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h47;
  wire          compressDataVec_hitReq_4_71 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h47;
  wire          compressDataVec_hitReq_5_71 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h47;
  wire          compressDataVec_hitReq_6_71 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h47;
  wire          compressDataVec_hitReq_7_71 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h47;
  wire          compressDataVec_hitReq_8_71 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h47;
  wire          compressDataVec_hitReq_9_71 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h47;
  wire          compressDataVec_hitReq_10_71 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h47;
  wire          compressDataVec_hitReq_11_71 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h47;
  wire          compressDataVec_hitReq_12_71 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h47;
  wire          compressDataVec_hitReq_13_71 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h47;
  wire          compressDataVec_hitReq_14_71 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h47;
  wire          compressDataVec_hitReq_15_71 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h47;
  wire          compressDataVec_hitReq_16_71 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h47;
  wire          compressDataVec_hitReq_17_71 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h47;
  wire          compressDataVec_hitReq_18_71 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h47;
  wire          compressDataVec_hitReq_19_71 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h47;
  wire          compressDataVec_hitReq_20_71 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h47;
  wire          compressDataVec_hitReq_21_71 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h47;
  wire          compressDataVec_hitReq_22_71 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h47;
  wire          compressDataVec_hitReq_23_71 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h47;
  wire          compressDataVec_hitReq_24_71 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h47;
  wire          compressDataVec_hitReq_25_71 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h47;
  wire          compressDataVec_hitReq_26_71 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h47;
  wire          compressDataVec_hitReq_27_71 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h47;
  wire          compressDataVec_hitReq_28_71 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h47;
  wire          compressDataVec_hitReq_29_71 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h47;
  wire          compressDataVec_hitReq_30_71 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h47;
  wire          compressDataVec_hitReq_31_71 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h47;
  wire          compressDataVec_hitReq_32_71 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h47;
  wire          compressDataVec_hitReq_33_71 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h47;
  wire          compressDataVec_hitReq_34_71 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h47;
  wire          compressDataVec_hitReq_35_71 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h47;
  wire          compressDataVec_hitReq_36_71 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h47;
  wire          compressDataVec_hitReq_37_71 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h47;
  wire          compressDataVec_hitReq_38_71 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h47;
  wire          compressDataVec_hitReq_39_71 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h47;
  wire          compressDataVec_hitReq_40_71 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h47;
  wire          compressDataVec_hitReq_41_71 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h47;
  wire          compressDataVec_hitReq_42_71 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h47;
  wire          compressDataVec_hitReq_43_71 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h47;
  wire          compressDataVec_hitReq_44_71 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h47;
  wire          compressDataVec_hitReq_45_71 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h47;
  wire          compressDataVec_hitReq_46_71 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h47;
  wire          compressDataVec_hitReq_47_71 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h47;
  wire          compressDataVec_hitReq_48_71 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h47;
  wire          compressDataVec_hitReq_49_71 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h47;
  wire          compressDataVec_hitReq_50_71 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h47;
  wire          compressDataVec_hitReq_51_71 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h47;
  wire          compressDataVec_hitReq_52_71 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h47;
  wire          compressDataVec_hitReq_53_71 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h47;
  wire          compressDataVec_hitReq_54_71 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h47;
  wire          compressDataVec_hitReq_55_71 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h47;
  wire          compressDataVec_hitReq_56_71 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h47;
  wire          compressDataVec_hitReq_57_71 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h47;
  wire          compressDataVec_hitReq_58_71 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h47;
  wire          compressDataVec_hitReq_59_71 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h47;
  wire          compressDataVec_hitReq_60_71 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h47;
  wire          compressDataVec_hitReq_61_71 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h47;
  wire          compressDataVec_hitReq_62_71 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h47;
  wire          compressDataVec_hitReq_63_71 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h47;
  wire [7:0]    compressDataVec_selectReqData_71 =
    (compressDataVec_hitReq_0_71 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_71 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_71 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_71 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_71 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_71 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_71 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_71 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_71 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_71 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_71 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_71 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_71 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_71 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_71 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_71 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_71 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_71 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_71 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_71 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_71 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_71 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_71 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_71 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_71 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_71 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_71 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_71 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_71 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_71 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_71 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_71 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_71 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_71 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_71 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_71 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_71 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_71 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_71 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_71 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_71 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_71 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_71 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_71 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_71 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_71 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_71 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_71 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_71 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_71 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_71 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_71 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_71 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_71 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_71 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_71 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_71 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_71 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_71 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_71 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_71 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_71 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_71 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_71 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_72 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h48;
  wire          compressDataVec_hitReq_1_72 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h48;
  wire          compressDataVec_hitReq_2_72 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h48;
  wire          compressDataVec_hitReq_3_72 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h48;
  wire          compressDataVec_hitReq_4_72 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h48;
  wire          compressDataVec_hitReq_5_72 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h48;
  wire          compressDataVec_hitReq_6_72 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h48;
  wire          compressDataVec_hitReq_7_72 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h48;
  wire          compressDataVec_hitReq_8_72 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h48;
  wire          compressDataVec_hitReq_9_72 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h48;
  wire          compressDataVec_hitReq_10_72 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h48;
  wire          compressDataVec_hitReq_11_72 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h48;
  wire          compressDataVec_hitReq_12_72 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h48;
  wire          compressDataVec_hitReq_13_72 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h48;
  wire          compressDataVec_hitReq_14_72 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h48;
  wire          compressDataVec_hitReq_15_72 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h48;
  wire          compressDataVec_hitReq_16_72 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h48;
  wire          compressDataVec_hitReq_17_72 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h48;
  wire          compressDataVec_hitReq_18_72 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h48;
  wire          compressDataVec_hitReq_19_72 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h48;
  wire          compressDataVec_hitReq_20_72 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h48;
  wire          compressDataVec_hitReq_21_72 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h48;
  wire          compressDataVec_hitReq_22_72 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h48;
  wire          compressDataVec_hitReq_23_72 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h48;
  wire          compressDataVec_hitReq_24_72 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h48;
  wire          compressDataVec_hitReq_25_72 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h48;
  wire          compressDataVec_hitReq_26_72 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h48;
  wire          compressDataVec_hitReq_27_72 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h48;
  wire          compressDataVec_hitReq_28_72 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h48;
  wire          compressDataVec_hitReq_29_72 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h48;
  wire          compressDataVec_hitReq_30_72 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h48;
  wire          compressDataVec_hitReq_31_72 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h48;
  wire          compressDataVec_hitReq_32_72 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h48;
  wire          compressDataVec_hitReq_33_72 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h48;
  wire          compressDataVec_hitReq_34_72 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h48;
  wire          compressDataVec_hitReq_35_72 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h48;
  wire          compressDataVec_hitReq_36_72 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h48;
  wire          compressDataVec_hitReq_37_72 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h48;
  wire          compressDataVec_hitReq_38_72 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h48;
  wire          compressDataVec_hitReq_39_72 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h48;
  wire          compressDataVec_hitReq_40_72 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h48;
  wire          compressDataVec_hitReq_41_72 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h48;
  wire          compressDataVec_hitReq_42_72 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h48;
  wire          compressDataVec_hitReq_43_72 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h48;
  wire          compressDataVec_hitReq_44_72 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h48;
  wire          compressDataVec_hitReq_45_72 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h48;
  wire          compressDataVec_hitReq_46_72 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h48;
  wire          compressDataVec_hitReq_47_72 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h48;
  wire          compressDataVec_hitReq_48_72 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h48;
  wire          compressDataVec_hitReq_49_72 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h48;
  wire          compressDataVec_hitReq_50_72 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h48;
  wire          compressDataVec_hitReq_51_72 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h48;
  wire          compressDataVec_hitReq_52_72 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h48;
  wire          compressDataVec_hitReq_53_72 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h48;
  wire          compressDataVec_hitReq_54_72 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h48;
  wire          compressDataVec_hitReq_55_72 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h48;
  wire          compressDataVec_hitReq_56_72 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h48;
  wire          compressDataVec_hitReq_57_72 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h48;
  wire          compressDataVec_hitReq_58_72 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h48;
  wire          compressDataVec_hitReq_59_72 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h48;
  wire          compressDataVec_hitReq_60_72 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h48;
  wire          compressDataVec_hitReq_61_72 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h48;
  wire          compressDataVec_hitReq_62_72 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h48;
  wire          compressDataVec_hitReq_63_72 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h48;
  wire [7:0]    compressDataVec_selectReqData_72 =
    (compressDataVec_hitReq_0_72 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_72 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_72 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_72 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_72 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_72 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_72 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_72 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_72 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_72 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_72 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_72 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_72 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_72 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_72 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_72 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_72 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_72 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_72 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_72 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_72 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_72 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_72 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_72 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_72 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_72 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_72 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_72 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_72 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_72 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_72 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_72 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_72 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_72 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_72 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_72 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_72 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_72 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_72 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_72 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_72 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_72 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_72 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_72 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_72 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_72 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_72 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_72 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_72 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_72 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_72 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_72 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_72 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_72 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_72 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_72 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_72 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_72 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_72 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_72 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_72 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_72 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_72 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_72 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_73 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h49;
  wire          compressDataVec_hitReq_1_73 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h49;
  wire          compressDataVec_hitReq_2_73 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h49;
  wire          compressDataVec_hitReq_3_73 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h49;
  wire          compressDataVec_hitReq_4_73 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h49;
  wire          compressDataVec_hitReq_5_73 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h49;
  wire          compressDataVec_hitReq_6_73 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h49;
  wire          compressDataVec_hitReq_7_73 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h49;
  wire          compressDataVec_hitReq_8_73 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h49;
  wire          compressDataVec_hitReq_9_73 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h49;
  wire          compressDataVec_hitReq_10_73 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h49;
  wire          compressDataVec_hitReq_11_73 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h49;
  wire          compressDataVec_hitReq_12_73 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h49;
  wire          compressDataVec_hitReq_13_73 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h49;
  wire          compressDataVec_hitReq_14_73 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h49;
  wire          compressDataVec_hitReq_15_73 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h49;
  wire          compressDataVec_hitReq_16_73 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h49;
  wire          compressDataVec_hitReq_17_73 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h49;
  wire          compressDataVec_hitReq_18_73 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h49;
  wire          compressDataVec_hitReq_19_73 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h49;
  wire          compressDataVec_hitReq_20_73 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h49;
  wire          compressDataVec_hitReq_21_73 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h49;
  wire          compressDataVec_hitReq_22_73 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h49;
  wire          compressDataVec_hitReq_23_73 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h49;
  wire          compressDataVec_hitReq_24_73 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h49;
  wire          compressDataVec_hitReq_25_73 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h49;
  wire          compressDataVec_hitReq_26_73 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h49;
  wire          compressDataVec_hitReq_27_73 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h49;
  wire          compressDataVec_hitReq_28_73 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h49;
  wire          compressDataVec_hitReq_29_73 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h49;
  wire          compressDataVec_hitReq_30_73 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h49;
  wire          compressDataVec_hitReq_31_73 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h49;
  wire          compressDataVec_hitReq_32_73 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h49;
  wire          compressDataVec_hitReq_33_73 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h49;
  wire          compressDataVec_hitReq_34_73 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h49;
  wire          compressDataVec_hitReq_35_73 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h49;
  wire          compressDataVec_hitReq_36_73 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h49;
  wire          compressDataVec_hitReq_37_73 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h49;
  wire          compressDataVec_hitReq_38_73 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h49;
  wire          compressDataVec_hitReq_39_73 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h49;
  wire          compressDataVec_hitReq_40_73 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h49;
  wire          compressDataVec_hitReq_41_73 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h49;
  wire          compressDataVec_hitReq_42_73 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h49;
  wire          compressDataVec_hitReq_43_73 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h49;
  wire          compressDataVec_hitReq_44_73 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h49;
  wire          compressDataVec_hitReq_45_73 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h49;
  wire          compressDataVec_hitReq_46_73 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h49;
  wire          compressDataVec_hitReq_47_73 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h49;
  wire          compressDataVec_hitReq_48_73 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h49;
  wire          compressDataVec_hitReq_49_73 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h49;
  wire          compressDataVec_hitReq_50_73 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h49;
  wire          compressDataVec_hitReq_51_73 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h49;
  wire          compressDataVec_hitReq_52_73 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h49;
  wire          compressDataVec_hitReq_53_73 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h49;
  wire          compressDataVec_hitReq_54_73 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h49;
  wire          compressDataVec_hitReq_55_73 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h49;
  wire          compressDataVec_hitReq_56_73 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h49;
  wire          compressDataVec_hitReq_57_73 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h49;
  wire          compressDataVec_hitReq_58_73 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h49;
  wire          compressDataVec_hitReq_59_73 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h49;
  wire          compressDataVec_hitReq_60_73 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h49;
  wire          compressDataVec_hitReq_61_73 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h49;
  wire          compressDataVec_hitReq_62_73 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h49;
  wire          compressDataVec_hitReq_63_73 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h49;
  wire [7:0]    compressDataVec_selectReqData_73 =
    (compressDataVec_hitReq_0_73 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_73 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_73 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_73 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_73 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_73 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_73 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_73 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_73 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_73 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_73 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_73 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_73 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_73 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_73 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_73 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_73 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_73 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_73 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_73 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_73 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_73 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_73 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_73 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_73 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_73 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_73 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_73 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_73 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_73 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_73 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_73 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_73 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_73 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_73 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_73 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_73 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_73 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_73 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_73 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_73 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_73 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_73 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_73 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_73 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_73 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_73 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_73 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_73 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_73 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_73 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_73 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_73 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_73 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_73 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_73 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_73 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_73 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_73 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_73 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_73 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_73 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_73 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_73 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_74 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h4A;
  wire          compressDataVec_hitReq_1_74 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h4A;
  wire          compressDataVec_hitReq_2_74 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h4A;
  wire          compressDataVec_hitReq_3_74 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h4A;
  wire          compressDataVec_hitReq_4_74 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h4A;
  wire          compressDataVec_hitReq_5_74 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h4A;
  wire          compressDataVec_hitReq_6_74 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h4A;
  wire          compressDataVec_hitReq_7_74 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h4A;
  wire          compressDataVec_hitReq_8_74 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h4A;
  wire          compressDataVec_hitReq_9_74 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h4A;
  wire          compressDataVec_hitReq_10_74 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h4A;
  wire          compressDataVec_hitReq_11_74 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h4A;
  wire          compressDataVec_hitReq_12_74 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h4A;
  wire          compressDataVec_hitReq_13_74 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h4A;
  wire          compressDataVec_hitReq_14_74 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h4A;
  wire          compressDataVec_hitReq_15_74 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h4A;
  wire          compressDataVec_hitReq_16_74 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h4A;
  wire          compressDataVec_hitReq_17_74 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h4A;
  wire          compressDataVec_hitReq_18_74 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h4A;
  wire          compressDataVec_hitReq_19_74 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h4A;
  wire          compressDataVec_hitReq_20_74 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h4A;
  wire          compressDataVec_hitReq_21_74 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h4A;
  wire          compressDataVec_hitReq_22_74 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h4A;
  wire          compressDataVec_hitReq_23_74 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h4A;
  wire          compressDataVec_hitReq_24_74 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h4A;
  wire          compressDataVec_hitReq_25_74 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h4A;
  wire          compressDataVec_hitReq_26_74 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h4A;
  wire          compressDataVec_hitReq_27_74 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h4A;
  wire          compressDataVec_hitReq_28_74 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h4A;
  wire          compressDataVec_hitReq_29_74 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h4A;
  wire          compressDataVec_hitReq_30_74 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h4A;
  wire          compressDataVec_hitReq_31_74 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h4A;
  wire          compressDataVec_hitReq_32_74 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h4A;
  wire          compressDataVec_hitReq_33_74 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h4A;
  wire          compressDataVec_hitReq_34_74 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h4A;
  wire          compressDataVec_hitReq_35_74 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h4A;
  wire          compressDataVec_hitReq_36_74 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h4A;
  wire          compressDataVec_hitReq_37_74 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h4A;
  wire          compressDataVec_hitReq_38_74 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h4A;
  wire          compressDataVec_hitReq_39_74 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h4A;
  wire          compressDataVec_hitReq_40_74 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h4A;
  wire          compressDataVec_hitReq_41_74 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h4A;
  wire          compressDataVec_hitReq_42_74 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h4A;
  wire          compressDataVec_hitReq_43_74 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h4A;
  wire          compressDataVec_hitReq_44_74 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h4A;
  wire          compressDataVec_hitReq_45_74 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h4A;
  wire          compressDataVec_hitReq_46_74 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h4A;
  wire          compressDataVec_hitReq_47_74 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h4A;
  wire          compressDataVec_hitReq_48_74 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h4A;
  wire          compressDataVec_hitReq_49_74 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h4A;
  wire          compressDataVec_hitReq_50_74 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h4A;
  wire          compressDataVec_hitReq_51_74 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h4A;
  wire          compressDataVec_hitReq_52_74 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h4A;
  wire          compressDataVec_hitReq_53_74 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h4A;
  wire          compressDataVec_hitReq_54_74 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h4A;
  wire          compressDataVec_hitReq_55_74 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h4A;
  wire          compressDataVec_hitReq_56_74 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h4A;
  wire          compressDataVec_hitReq_57_74 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h4A;
  wire          compressDataVec_hitReq_58_74 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h4A;
  wire          compressDataVec_hitReq_59_74 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h4A;
  wire          compressDataVec_hitReq_60_74 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h4A;
  wire          compressDataVec_hitReq_61_74 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h4A;
  wire          compressDataVec_hitReq_62_74 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h4A;
  wire          compressDataVec_hitReq_63_74 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h4A;
  wire [7:0]    compressDataVec_selectReqData_74 =
    (compressDataVec_hitReq_0_74 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_74 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_74 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_74 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_74 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_74 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_74 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_74 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_74 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_74 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_74 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_74 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_74 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_74 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_74 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_74 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_74 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_74 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_74 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_74 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_74 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_74 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_74 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_74 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_74 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_74 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_74 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_74 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_74 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_74 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_74 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_74 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_74 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_74 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_74 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_74 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_74 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_74 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_74 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_74 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_74 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_74 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_74 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_74 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_74 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_74 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_74 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_74 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_74 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_74 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_74 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_74 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_74 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_74 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_74 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_74 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_74 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_74 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_74 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_74 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_74 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_74 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_74 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_74 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_75 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h4B;
  wire          compressDataVec_hitReq_1_75 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h4B;
  wire          compressDataVec_hitReq_2_75 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h4B;
  wire          compressDataVec_hitReq_3_75 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h4B;
  wire          compressDataVec_hitReq_4_75 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h4B;
  wire          compressDataVec_hitReq_5_75 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h4B;
  wire          compressDataVec_hitReq_6_75 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h4B;
  wire          compressDataVec_hitReq_7_75 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h4B;
  wire          compressDataVec_hitReq_8_75 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h4B;
  wire          compressDataVec_hitReq_9_75 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h4B;
  wire          compressDataVec_hitReq_10_75 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h4B;
  wire          compressDataVec_hitReq_11_75 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h4B;
  wire          compressDataVec_hitReq_12_75 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h4B;
  wire          compressDataVec_hitReq_13_75 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h4B;
  wire          compressDataVec_hitReq_14_75 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h4B;
  wire          compressDataVec_hitReq_15_75 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h4B;
  wire          compressDataVec_hitReq_16_75 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h4B;
  wire          compressDataVec_hitReq_17_75 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h4B;
  wire          compressDataVec_hitReq_18_75 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h4B;
  wire          compressDataVec_hitReq_19_75 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h4B;
  wire          compressDataVec_hitReq_20_75 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h4B;
  wire          compressDataVec_hitReq_21_75 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h4B;
  wire          compressDataVec_hitReq_22_75 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h4B;
  wire          compressDataVec_hitReq_23_75 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h4B;
  wire          compressDataVec_hitReq_24_75 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h4B;
  wire          compressDataVec_hitReq_25_75 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h4B;
  wire          compressDataVec_hitReq_26_75 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h4B;
  wire          compressDataVec_hitReq_27_75 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h4B;
  wire          compressDataVec_hitReq_28_75 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h4B;
  wire          compressDataVec_hitReq_29_75 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h4B;
  wire          compressDataVec_hitReq_30_75 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h4B;
  wire          compressDataVec_hitReq_31_75 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h4B;
  wire          compressDataVec_hitReq_32_75 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h4B;
  wire          compressDataVec_hitReq_33_75 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h4B;
  wire          compressDataVec_hitReq_34_75 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h4B;
  wire          compressDataVec_hitReq_35_75 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h4B;
  wire          compressDataVec_hitReq_36_75 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h4B;
  wire          compressDataVec_hitReq_37_75 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h4B;
  wire          compressDataVec_hitReq_38_75 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h4B;
  wire          compressDataVec_hitReq_39_75 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h4B;
  wire          compressDataVec_hitReq_40_75 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h4B;
  wire          compressDataVec_hitReq_41_75 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h4B;
  wire          compressDataVec_hitReq_42_75 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h4B;
  wire          compressDataVec_hitReq_43_75 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h4B;
  wire          compressDataVec_hitReq_44_75 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h4B;
  wire          compressDataVec_hitReq_45_75 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h4B;
  wire          compressDataVec_hitReq_46_75 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h4B;
  wire          compressDataVec_hitReq_47_75 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h4B;
  wire          compressDataVec_hitReq_48_75 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h4B;
  wire          compressDataVec_hitReq_49_75 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h4B;
  wire          compressDataVec_hitReq_50_75 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h4B;
  wire          compressDataVec_hitReq_51_75 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h4B;
  wire          compressDataVec_hitReq_52_75 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h4B;
  wire          compressDataVec_hitReq_53_75 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h4B;
  wire          compressDataVec_hitReq_54_75 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h4B;
  wire          compressDataVec_hitReq_55_75 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h4B;
  wire          compressDataVec_hitReq_56_75 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h4B;
  wire          compressDataVec_hitReq_57_75 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h4B;
  wire          compressDataVec_hitReq_58_75 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h4B;
  wire          compressDataVec_hitReq_59_75 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h4B;
  wire          compressDataVec_hitReq_60_75 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h4B;
  wire          compressDataVec_hitReq_61_75 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h4B;
  wire          compressDataVec_hitReq_62_75 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h4B;
  wire          compressDataVec_hitReq_63_75 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h4B;
  wire [7:0]    compressDataVec_selectReqData_75 =
    (compressDataVec_hitReq_0_75 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_75 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_75 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_75 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_75 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_75 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_75 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_75 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_75 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_75 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_75 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_75 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_75 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_75 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_75 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_75 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_75 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_75 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_75 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_75 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_75 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_75 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_75 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_75 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_75 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_75 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_75 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_75 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_75 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_75 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_75 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_75 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_75 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_75 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_75 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_75 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_75 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_75 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_75 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_75 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_75 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_75 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_75 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_75 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_75 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_75 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_75 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_75 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_75 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_75 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_75 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_75 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_75 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_75 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_75 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_75 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_75 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_75 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_75 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_75 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_75 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_75 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_75 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_75 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_76 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h4C;
  wire          compressDataVec_hitReq_1_76 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h4C;
  wire          compressDataVec_hitReq_2_76 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h4C;
  wire          compressDataVec_hitReq_3_76 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h4C;
  wire          compressDataVec_hitReq_4_76 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h4C;
  wire          compressDataVec_hitReq_5_76 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h4C;
  wire          compressDataVec_hitReq_6_76 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h4C;
  wire          compressDataVec_hitReq_7_76 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h4C;
  wire          compressDataVec_hitReq_8_76 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h4C;
  wire          compressDataVec_hitReq_9_76 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h4C;
  wire          compressDataVec_hitReq_10_76 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h4C;
  wire          compressDataVec_hitReq_11_76 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h4C;
  wire          compressDataVec_hitReq_12_76 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h4C;
  wire          compressDataVec_hitReq_13_76 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h4C;
  wire          compressDataVec_hitReq_14_76 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h4C;
  wire          compressDataVec_hitReq_15_76 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h4C;
  wire          compressDataVec_hitReq_16_76 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h4C;
  wire          compressDataVec_hitReq_17_76 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h4C;
  wire          compressDataVec_hitReq_18_76 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h4C;
  wire          compressDataVec_hitReq_19_76 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h4C;
  wire          compressDataVec_hitReq_20_76 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h4C;
  wire          compressDataVec_hitReq_21_76 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h4C;
  wire          compressDataVec_hitReq_22_76 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h4C;
  wire          compressDataVec_hitReq_23_76 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h4C;
  wire          compressDataVec_hitReq_24_76 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h4C;
  wire          compressDataVec_hitReq_25_76 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h4C;
  wire          compressDataVec_hitReq_26_76 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h4C;
  wire          compressDataVec_hitReq_27_76 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h4C;
  wire          compressDataVec_hitReq_28_76 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h4C;
  wire          compressDataVec_hitReq_29_76 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h4C;
  wire          compressDataVec_hitReq_30_76 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h4C;
  wire          compressDataVec_hitReq_31_76 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h4C;
  wire          compressDataVec_hitReq_32_76 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h4C;
  wire          compressDataVec_hitReq_33_76 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h4C;
  wire          compressDataVec_hitReq_34_76 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h4C;
  wire          compressDataVec_hitReq_35_76 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h4C;
  wire          compressDataVec_hitReq_36_76 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h4C;
  wire          compressDataVec_hitReq_37_76 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h4C;
  wire          compressDataVec_hitReq_38_76 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h4C;
  wire          compressDataVec_hitReq_39_76 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h4C;
  wire          compressDataVec_hitReq_40_76 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h4C;
  wire          compressDataVec_hitReq_41_76 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h4C;
  wire          compressDataVec_hitReq_42_76 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h4C;
  wire          compressDataVec_hitReq_43_76 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h4C;
  wire          compressDataVec_hitReq_44_76 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h4C;
  wire          compressDataVec_hitReq_45_76 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h4C;
  wire          compressDataVec_hitReq_46_76 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h4C;
  wire          compressDataVec_hitReq_47_76 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h4C;
  wire          compressDataVec_hitReq_48_76 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h4C;
  wire          compressDataVec_hitReq_49_76 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h4C;
  wire          compressDataVec_hitReq_50_76 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h4C;
  wire          compressDataVec_hitReq_51_76 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h4C;
  wire          compressDataVec_hitReq_52_76 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h4C;
  wire          compressDataVec_hitReq_53_76 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h4C;
  wire          compressDataVec_hitReq_54_76 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h4C;
  wire          compressDataVec_hitReq_55_76 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h4C;
  wire          compressDataVec_hitReq_56_76 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h4C;
  wire          compressDataVec_hitReq_57_76 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h4C;
  wire          compressDataVec_hitReq_58_76 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h4C;
  wire          compressDataVec_hitReq_59_76 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h4C;
  wire          compressDataVec_hitReq_60_76 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h4C;
  wire          compressDataVec_hitReq_61_76 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h4C;
  wire          compressDataVec_hitReq_62_76 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h4C;
  wire          compressDataVec_hitReq_63_76 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h4C;
  wire [7:0]    compressDataVec_selectReqData_76 =
    (compressDataVec_hitReq_0_76 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_76 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_76 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_76 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_76 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_76 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_76 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_76 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_76 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_76 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_76 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_76 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_76 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_76 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_76 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_76 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_76 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_76 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_76 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_76 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_76 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_76 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_76 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_76 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_76 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_76 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_76 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_76 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_76 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_76 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_76 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_76 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_76 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_76 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_76 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_76 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_76 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_76 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_76 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_76 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_76 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_76 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_76 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_76 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_76 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_76 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_76 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_76 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_76 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_76 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_76 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_76 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_76 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_76 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_76 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_76 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_76 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_76 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_76 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_76 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_76 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_76 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_76 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_76 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_77 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h4D;
  wire          compressDataVec_hitReq_1_77 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h4D;
  wire          compressDataVec_hitReq_2_77 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h4D;
  wire          compressDataVec_hitReq_3_77 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h4D;
  wire          compressDataVec_hitReq_4_77 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h4D;
  wire          compressDataVec_hitReq_5_77 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h4D;
  wire          compressDataVec_hitReq_6_77 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h4D;
  wire          compressDataVec_hitReq_7_77 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h4D;
  wire          compressDataVec_hitReq_8_77 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h4D;
  wire          compressDataVec_hitReq_9_77 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h4D;
  wire          compressDataVec_hitReq_10_77 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h4D;
  wire          compressDataVec_hitReq_11_77 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h4D;
  wire          compressDataVec_hitReq_12_77 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h4D;
  wire          compressDataVec_hitReq_13_77 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h4D;
  wire          compressDataVec_hitReq_14_77 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h4D;
  wire          compressDataVec_hitReq_15_77 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h4D;
  wire          compressDataVec_hitReq_16_77 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h4D;
  wire          compressDataVec_hitReq_17_77 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h4D;
  wire          compressDataVec_hitReq_18_77 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h4D;
  wire          compressDataVec_hitReq_19_77 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h4D;
  wire          compressDataVec_hitReq_20_77 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h4D;
  wire          compressDataVec_hitReq_21_77 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h4D;
  wire          compressDataVec_hitReq_22_77 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h4D;
  wire          compressDataVec_hitReq_23_77 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h4D;
  wire          compressDataVec_hitReq_24_77 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h4D;
  wire          compressDataVec_hitReq_25_77 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h4D;
  wire          compressDataVec_hitReq_26_77 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h4D;
  wire          compressDataVec_hitReq_27_77 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h4D;
  wire          compressDataVec_hitReq_28_77 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h4D;
  wire          compressDataVec_hitReq_29_77 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h4D;
  wire          compressDataVec_hitReq_30_77 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h4D;
  wire          compressDataVec_hitReq_31_77 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h4D;
  wire          compressDataVec_hitReq_32_77 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h4D;
  wire          compressDataVec_hitReq_33_77 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h4D;
  wire          compressDataVec_hitReq_34_77 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h4D;
  wire          compressDataVec_hitReq_35_77 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h4D;
  wire          compressDataVec_hitReq_36_77 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h4D;
  wire          compressDataVec_hitReq_37_77 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h4D;
  wire          compressDataVec_hitReq_38_77 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h4D;
  wire          compressDataVec_hitReq_39_77 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h4D;
  wire          compressDataVec_hitReq_40_77 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h4D;
  wire          compressDataVec_hitReq_41_77 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h4D;
  wire          compressDataVec_hitReq_42_77 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h4D;
  wire          compressDataVec_hitReq_43_77 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h4D;
  wire          compressDataVec_hitReq_44_77 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h4D;
  wire          compressDataVec_hitReq_45_77 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h4D;
  wire          compressDataVec_hitReq_46_77 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h4D;
  wire          compressDataVec_hitReq_47_77 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h4D;
  wire          compressDataVec_hitReq_48_77 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h4D;
  wire          compressDataVec_hitReq_49_77 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h4D;
  wire          compressDataVec_hitReq_50_77 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h4D;
  wire          compressDataVec_hitReq_51_77 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h4D;
  wire          compressDataVec_hitReq_52_77 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h4D;
  wire          compressDataVec_hitReq_53_77 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h4D;
  wire          compressDataVec_hitReq_54_77 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h4D;
  wire          compressDataVec_hitReq_55_77 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h4D;
  wire          compressDataVec_hitReq_56_77 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h4D;
  wire          compressDataVec_hitReq_57_77 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h4D;
  wire          compressDataVec_hitReq_58_77 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h4D;
  wire          compressDataVec_hitReq_59_77 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h4D;
  wire          compressDataVec_hitReq_60_77 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h4D;
  wire          compressDataVec_hitReq_61_77 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h4D;
  wire          compressDataVec_hitReq_62_77 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h4D;
  wire          compressDataVec_hitReq_63_77 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h4D;
  wire [7:0]    compressDataVec_selectReqData_77 =
    (compressDataVec_hitReq_0_77 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_77 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_77 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_77 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_77 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_77 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_77 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_77 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_77 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_77 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_77 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_77 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_77 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_77 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_77 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_77 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_77 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_77 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_77 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_77 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_77 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_77 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_77 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_77 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_77 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_77 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_77 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_77 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_77 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_77 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_77 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_77 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_77 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_77 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_77 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_77 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_77 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_77 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_77 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_77 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_77 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_77 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_77 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_77 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_77 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_77 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_77 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_77 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_77 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_77 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_77 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_77 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_77 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_77 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_77 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_77 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_77 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_77 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_77 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_77 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_77 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_77 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_77 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_77 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_78 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h4E;
  wire          compressDataVec_hitReq_1_78 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h4E;
  wire          compressDataVec_hitReq_2_78 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h4E;
  wire          compressDataVec_hitReq_3_78 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h4E;
  wire          compressDataVec_hitReq_4_78 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h4E;
  wire          compressDataVec_hitReq_5_78 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h4E;
  wire          compressDataVec_hitReq_6_78 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h4E;
  wire          compressDataVec_hitReq_7_78 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h4E;
  wire          compressDataVec_hitReq_8_78 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h4E;
  wire          compressDataVec_hitReq_9_78 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h4E;
  wire          compressDataVec_hitReq_10_78 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h4E;
  wire          compressDataVec_hitReq_11_78 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h4E;
  wire          compressDataVec_hitReq_12_78 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h4E;
  wire          compressDataVec_hitReq_13_78 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h4E;
  wire          compressDataVec_hitReq_14_78 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h4E;
  wire          compressDataVec_hitReq_15_78 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h4E;
  wire          compressDataVec_hitReq_16_78 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h4E;
  wire          compressDataVec_hitReq_17_78 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h4E;
  wire          compressDataVec_hitReq_18_78 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h4E;
  wire          compressDataVec_hitReq_19_78 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h4E;
  wire          compressDataVec_hitReq_20_78 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h4E;
  wire          compressDataVec_hitReq_21_78 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h4E;
  wire          compressDataVec_hitReq_22_78 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h4E;
  wire          compressDataVec_hitReq_23_78 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h4E;
  wire          compressDataVec_hitReq_24_78 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h4E;
  wire          compressDataVec_hitReq_25_78 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h4E;
  wire          compressDataVec_hitReq_26_78 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h4E;
  wire          compressDataVec_hitReq_27_78 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h4E;
  wire          compressDataVec_hitReq_28_78 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h4E;
  wire          compressDataVec_hitReq_29_78 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h4E;
  wire          compressDataVec_hitReq_30_78 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h4E;
  wire          compressDataVec_hitReq_31_78 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h4E;
  wire          compressDataVec_hitReq_32_78 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h4E;
  wire          compressDataVec_hitReq_33_78 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h4E;
  wire          compressDataVec_hitReq_34_78 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h4E;
  wire          compressDataVec_hitReq_35_78 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h4E;
  wire          compressDataVec_hitReq_36_78 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h4E;
  wire          compressDataVec_hitReq_37_78 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h4E;
  wire          compressDataVec_hitReq_38_78 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h4E;
  wire          compressDataVec_hitReq_39_78 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h4E;
  wire          compressDataVec_hitReq_40_78 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h4E;
  wire          compressDataVec_hitReq_41_78 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h4E;
  wire          compressDataVec_hitReq_42_78 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h4E;
  wire          compressDataVec_hitReq_43_78 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h4E;
  wire          compressDataVec_hitReq_44_78 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h4E;
  wire          compressDataVec_hitReq_45_78 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h4E;
  wire          compressDataVec_hitReq_46_78 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h4E;
  wire          compressDataVec_hitReq_47_78 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h4E;
  wire          compressDataVec_hitReq_48_78 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h4E;
  wire          compressDataVec_hitReq_49_78 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h4E;
  wire          compressDataVec_hitReq_50_78 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h4E;
  wire          compressDataVec_hitReq_51_78 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h4E;
  wire          compressDataVec_hitReq_52_78 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h4E;
  wire          compressDataVec_hitReq_53_78 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h4E;
  wire          compressDataVec_hitReq_54_78 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h4E;
  wire          compressDataVec_hitReq_55_78 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h4E;
  wire          compressDataVec_hitReq_56_78 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h4E;
  wire          compressDataVec_hitReq_57_78 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h4E;
  wire          compressDataVec_hitReq_58_78 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h4E;
  wire          compressDataVec_hitReq_59_78 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h4E;
  wire          compressDataVec_hitReq_60_78 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h4E;
  wire          compressDataVec_hitReq_61_78 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h4E;
  wire          compressDataVec_hitReq_62_78 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h4E;
  wire          compressDataVec_hitReq_63_78 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h4E;
  wire [7:0]    compressDataVec_selectReqData_78 =
    (compressDataVec_hitReq_0_78 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_78 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_78 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_78 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_78 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_78 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_78 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_78 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_78 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_78 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_78 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_78 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_78 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_78 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_78 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_78 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_78 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_78 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_78 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_78 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_78 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_78 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_78 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_78 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_78 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_78 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_78 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_78 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_78 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_78 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_78 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_78 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_78 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_78 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_78 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_78 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_78 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_78 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_78 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_78 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_78 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_78 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_78 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_78 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_78 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_78 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_78 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_78 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_78 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_78 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_78 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_78 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_78 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_78 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_78 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_78 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_78 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_78 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_78 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_78 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_78 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_78 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_78 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_78 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_79 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h4F;
  wire          compressDataVec_hitReq_1_79 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h4F;
  wire          compressDataVec_hitReq_2_79 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h4F;
  wire          compressDataVec_hitReq_3_79 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h4F;
  wire          compressDataVec_hitReq_4_79 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h4F;
  wire          compressDataVec_hitReq_5_79 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h4F;
  wire          compressDataVec_hitReq_6_79 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h4F;
  wire          compressDataVec_hitReq_7_79 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h4F;
  wire          compressDataVec_hitReq_8_79 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h4F;
  wire          compressDataVec_hitReq_9_79 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h4F;
  wire          compressDataVec_hitReq_10_79 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h4F;
  wire          compressDataVec_hitReq_11_79 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h4F;
  wire          compressDataVec_hitReq_12_79 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h4F;
  wire          compressDataVec_hitReq_13_79 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h4F;
  wire          compressDataVec_hitReq_14_79 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h4F;
  wire          compressDataVec_hitReq_15_79 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h4F;
  wire          compressDataVec_hitReq_16_79 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h4F;
  wire          compressDataVec_hitReq_17_79 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h4F;
  wire          compressDataVec_hitReq_18_79 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h4F;
  wire          compressDataVec_hitReq_19_79 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h4F;
  wire          compressDataVec_hitReq_20_79 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h4F;
  wire          compressDataVec_hitReq_21_79 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h4F;
  wire          compressDataVec_hitReq_22_79 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h4F;
  wire          compressDataVec_hitReq_23_79 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h4F;
  wire          compressDataVec_hitReq_24_79 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h4F;
  wire          compressDataVec_hitReq_25_79 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h4F;
  wire          compressDataVec_hitReq_26_79 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h4F;
  wire          compressDataVec_hitReq_27_79 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h4F;
  wire          compressDataVec_hitReq_28_79 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h4F;
  wire          compressDataVec_hitReq_29_79 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h4F;
  wire          compressDataVec_hitReq_30_79 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h4F;
  wire          compressDataVec_hitReq_31_79 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h4F;
  wire          compressDataVec_hitReq_32_79 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h4F;
  wire          compressDataVec_hitReq_33_79 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h4F;
  wire          compressDataVec_hitReq_34_79 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h4F;
  wire          compressDataVec_hitReq_35_79 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h4F;
  wire          compressDataVec_hitReq_36_79 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h4F;
  wire          compressDataVec_hitReq_37_79 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h4F;
  wire          compressDataVec_hitReq_38_79 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h4F;
  wire          compressDataVec_hitReq_39_79 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h4F;
  wire          compressDataVec_hitReq_40_79 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h4F;
  wire          compressDataVec_hitReq_41_79 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h4F;
  wire          compressDataVec_hitReq_42_79 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h4F;
  wire          compressDataVec_hitReq_43_79 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h4F;
  wire          compressDataVec_hitReq_44_79 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h4F;
  wire          compressDataVec_hitReq_45_79 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h4F;
  wire          compressDataVec_hitReq_46_79 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h4F;
  wire          compressDataVec_hitReq_47_79 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h4F;
  wire          compressDataVec_hitReq_48_79 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h4F;
  wire          compressDataVec_hitReq_49_79 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h4F;
  wire          compressDataVec_hitReq_50_79 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h4F;
  wire          compressDataVec_hitReq_51_79 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h4F;
  wire          compressDataVec_hitReq_52_79 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h4F;
  wire          compressDataVec_hitReq_53_79 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h4F;
  wire          compressDataVec_hitReq_54_79 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h4F;
  wire          compressDataVec_hitReq_55_79 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h4F;
  wire          compressDataVec_hitReq_56_79 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h4F;
  wire          compressDataVec_hitReq_57_79 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h4F;
  wire          compressDataVec_hitReq_58_79 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h4F;
  wire          compressDataVec_hitReq_59_79 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h4F;
  wire          compressDataVec_hitReq_60_79 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h4F;
  wire          compressDataVec_hitReq_61_79 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h4F;
  wire          compressDataVec_hitReq_62_79 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h4F;
  wire          compressDataVec_hitReq_63_79 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h4F;
  wire [7:0]    compressDataVec_selectReqData_79 =
    (compressDataVec_hitReq_0_79 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_79 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_79 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_79 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_79 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_79 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_79 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_79 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_79 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_79 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_79 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_79 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_79 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_79 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_79 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_79 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_79 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_79 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_79 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_79 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_79 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_79 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_79 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_79 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_79 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_79 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_79 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_79 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_79 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_79 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_79 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_79 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_79 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_79 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_79 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_79 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_79 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_79 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_79 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_79 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_79 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_79 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_79 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_79 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_79 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_79 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_79 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_79 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_79 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_79 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_79 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_79 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_79 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_79 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_79 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_79 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_79 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_79 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_79 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_79 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_79 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_79 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_79 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_79 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_80 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h50;
  wire          compressDataVec_hitReq_1_80 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h50;
  wire          compressDataVec_hitReq_2_80 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h50;
  wire          compressDataVec_hitReq_3_80 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h50;
  wire          compressDataVec_hitReq_4_80 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h50;
  wire          compressDataVec_hitReq_5_80 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h50;
  wire          compressDataVec_hitReq_6_80 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h50;
  wire          compressDataVec_hitReq_7_80 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h50;
  wire          compressDataVec_hitReq_8_80 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h50;
  wire          compressDataVec_hitReq_9_80 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h50;
  wire          compressDataVec_hitReq_10_80 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h50;
  wire          compressDataVec_hitReq_11_80 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h50;
  wire          compressDataVec_hitReq_12_80 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h50;
  wire          compressDataVec_hitReq_13_80 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h50;
  wire          compressDataVec_hitReq_14_80 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h50;
  wire          compressDataVec_hitReq_15_80 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h50;
  wire          compressDataVec_hitReq_16_80 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h50;
  wire          compressDataVec_hitReq_17_80 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h50;
  wire          compressDataVec_hitReq_18_80 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h50;
  wire          compressDataVec_hitReq_19_80 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h50;
  wire          compressDataVec_hitReq_20_80 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h50;
  wire          compressDataVec_hitReq_21_80 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h50;
  wire          compressDataVec_hitReq_22_80 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h50;
  wire          compressDataVec_hitReq_23_80 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h50;
  wire          compressDataVec_hitReq_24_80 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h50;
  wire          compressDataVec_hitReq_25_80 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h50;
  wire          compressDataVec_hitReq_26_80 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h50;
  wire          compressDataVec_hitReq_27_80 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h50;
  wire          compressDataVec_hitReq_28_80 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h50;
  wire          compressDataVec_hitReq_29_80 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h50;
  wire          compressDataVec_hitReq_30_80 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h50;
  wire          compressDataVec_hitReq_31_80 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h50;
  wire          compressDataVec_hitReq_32_80 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h50;
  wire          compressDataVec_hitReq_33_80 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h50;
  wire          compressDataVec_hitReq_34_80 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h50;
  wire          compressDataVec_hitReq_35_80 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h50;
  wire          compressDataVec_hitReq_36_80 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h50;
  wire          compressDataVec_hitReq_37_80 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h50;
  wire          compressDataVec_hitReq_38_80 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h50;
  wire          compressDataVec_hitReq_39_80 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h50;
  wire          compressDataVec_hitReq_40_80 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h50;
  wire          compressDataVec_hitReq_41_80 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h50;
  wire          compressDataVec_hitReq_42_80 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h50;
  wire          compressDataVec_hitReq_43_80 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h50;
  wire          compressDataVec_hitReq_44_80 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h50;
  wire          compressDataVec_hitReq_45_80 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h50;
  wire          compressDataVec_hitReq_46_80 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h50;
  wire          compressDataVec_hitReq_47_80 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h50;
  wire          compressDataVec_hitReq_48_80 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h50;
  wire          compressDataVec_hitReq_49_80 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h50;
  wire          compressDataVec_hitReq_50_80 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h50;
  wire          compressDataVec_hitReq_51_80 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h50;
  wire          compressDataVec_hitReq_52_80 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h50;
  wire          compressDataVec_hitReq_53_80 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h50;
  wire          compressDataVec_hitReq_54_80 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h50;
  wire          compressDataVec_hitReq_55_80 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h50;
  wire          compressDataVec_hitReq_56_80 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h50;
  wire          compressDataVec_hitReq_57_80 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h50;
  wire          compressDataVec_hitReq_58_80 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h50;
  wire          compressDataVec_hitReq_59_80 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h50;
  wire          compressDataVec_hitReq_60_80 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h50;
  wire          compressDataVec_hitReq_61_80 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h50;
  wire          compressDataVec_hitReq_62_80 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h50;
  wire          compressDataVec_hitReq_63_80 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h50;
  wire [7:0]    compressDataVec_selectReqData_80 =
    (compressDataVec_hitReq_0_80 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_80 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_80 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_80 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_80 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_80 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_80 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_80 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_80 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_80 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_80 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_80 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_80 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_80 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_80 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_80 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_80 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_80 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_80 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_80 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_80 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_80 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_80 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_80 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_80 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_80 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_80 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_80 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_80 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_80 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_80 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_80 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_80 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_80 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_80 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_80 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_80 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_80 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_80 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_80 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_80 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_80 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_80 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_80 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_80 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_80 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_80 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_80 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_80 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_80 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_80 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_80 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_80 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_80 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_80 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_80 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_80 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_80 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_80 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_80 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_80 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_80 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_80 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_80 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_81 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h51;
  wire          compressDataVec_hitReq_1_81 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h51;
  wire          compressDataVec_hitReq_2_81 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h51;
  wire          compressDataVec_hitReq_3_81 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h51;
  wire          compressDataVec_hitReq_4_81 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h51;
  wire          compressDataVec_hitReq_5_81 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h51;
  wire          compressDataVec_hitReq_6_81 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h51;
  wire          compressDataVec_hitReq_7_81 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h51;
  wire          compressDataVec_hitReq_8_81 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h51;
  wire          compressDataVec_hitReq_9_81 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h51;
  wire          compressDataVec_hitReq_10_81 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h51;
  wire          compressDataVec_hitReq_11_81 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h51;
  wire          compressDataVec_hitReq_12_81 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h51;
  wire          compressDataVec_hitReq_13_81 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h51;
  wire          compressDataVec_hitReq_14_81 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h51;
  wire          compressDataVec_hitReq_15_81 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h51;
  wire          compressDataVec_hitReq_16_81 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h51;
  wire          compressDataVec_hitReq_17_81 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h51;
  wire          compressDataVec_hitReq_18_81 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h51;
  wire          compressDataVec_hitReq_19_81 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h51;
  wire          compressDataVec_hitReq_20_81 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h51;
  wire          compressDataVec_hitReq_21_81 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h51;
  wire          compressDataVec_hitReq_22_81 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h51;
  wire          compressDataVec_hitReq_23_81 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h51;
  wire          compressDataVec_hitReq_24_81 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h51;
  wire          compressDataVec_hitReq_25_81 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h51;
  wire          compressDataVec_hitReq_26_81 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h51;
  wire          compressDataVec_hitReq_27_81 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h51;
  wire          compressDataVec_hitReq_28_81 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h51;
  wire          compressDataVec_hitReq_29_81 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h51;
  wire          compressDataVec_hitReq_30_81 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h51;
  wire          compressDataVec_hitReq_31_81 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h51;
  wire          compressDataVec_hitReq_32_81 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h51;
  wire          compressDataVec_hitReq_33_81 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h51;
  wire          compressDataVec_hitReq_34_81 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h51;
  wire          compressDataVec_hitReq_35_81 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h51;
  wire          compressDataVec_hitReq_36_81 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h51;
  wire          compressDataVec_hitReq_37_81 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h51;
  wire          compressDataVec_hitReq_38_81 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h51;
  wire          compressDataVec_hitReq_39_81 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h51;
  wire          compressDataVec_hitReq_40_81 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h51;
  wire          compressDataVec_hitReq_41_81 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h51;
  wire          compressDataVec_hitReq_42_81 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h51;
  wire          compressDataVec_hitReq_43_81 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h51;
  wire          compressDataVec_hitReq_44_81 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h51;
  wire          compressDataVec_hitReq_45_81 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h51;
  wire          compressDataVec_hitReq_46_81 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h51;
  wire          compressDataVec_hitReq_47_81 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h51;
  wire          compressDataVec_hitReq_48_81 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h51;
  wire          compressDataVec_hitReq_49_81 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h51;
  wire          compressDataVec_hitReq_50_81 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h51;
  wire          compressDataVec_hitReq_51_81 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h51;
  wire          compressDataVec_hitReq_52_81 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h51;
  wire          compressDataVec_hitReq_53_81 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h51;
  wire          compressDataVec_hitReq_54_81 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h51;
  wire          compressDataVec_hitReq_55_81 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h51;
  wire          compressDataVec_hitReq_56_81 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h51;
  wire          compressDataVec_hitReq_57_81 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h51;
  wire          compressDataVec_hitReq_58_81 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h51;
  wire          compressDataVec_hitReq_59_81 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h51;
  wire          compressDataVec_hitReq_60_81 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h51;
  wire          compressDataVec_hitReq_61_81 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h51;
  wire          compressDataVec_hitReq_62_81 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h51;
  wire          compressDataVec_hitReq_63_81 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h51;
  wire [7:0]    compressDataVec_selectReqData_81 =
    (compressDataVec_hitReq_0_81 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_81 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_81 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_81 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_81 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_81 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_81 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_81 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_81 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_81 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_81 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_81 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_81 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_81 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_81 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_81 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_81 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_81 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_81 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_81 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_81 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_81 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_81 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_81 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_81 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_81 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_81 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_81 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_81 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_81 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_81 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_81 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_81 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_81 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_81 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_81 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_81 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_81 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_81 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_81 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_81 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_81 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_81 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_81 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_81 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_81 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_81 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_81 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_81 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_81 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_81 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_81 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_81 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_81 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_81 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_81 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_81 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_81 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_81 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_81 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_81 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_81 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_81 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_81 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_82 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h52;
  wire          compressDataVec_hitReq_1_82 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h52;
  wire          compressDataVec_hitReq_2_82 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h52;
  wire          compressDataVec_hitReq_3_82 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h52;
  wire          compressDataVec_hitReq_4_82 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h52;
  wire          compressDataVec_hitReq_5_82 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h52;
  wire          compressDataVec_hitReq_6_82 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h52;
  wire          compressDataVec_hitReq_7_82 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h52;
  wire          compressDataVec_hitReq_8_82 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h52;
  wire          compressDataVec_hitReq_9_82 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h52;
  wire          compressDataVec_hitReq_10_82 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h52;
  wire          compressDataVec_hitReq_11_82 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h52;
  wire          compressDataVec_hitReq_12_82 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h52;
  wire          compressDataVec_hitReq_13_82 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h52;
  wire          compressDataVec_hitReq_14_82 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h52;
  wire          compressDataVec_hitReq_15_82 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h52;
  wire          compressDataVec_hitReq_16_82 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h52;
  wire          compressDataVec_hitReq_17_82 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h52;
  wire          compressDataVec_hitReq_18_82 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h52;
  wire          compressDataVec_hitReq_19_82 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h52;
  wire          compressDataVec_hitReq_20_82 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h52;
  wire          compressDataVec_hitReq_21_82 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h52;
  wire          compressDataVec_hitReq_22_82 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h52;
  wire          compressDataVec_hitReq_23_82 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h52;
  wire          compressDataVec_hitReq_24_82 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h52;
  wire          compressDataVec_hitReq_25_82 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h52;
  wire          compressDataVec_hitReq_26_82 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h52;
  wire          compressDataVec_hitReq_27_82 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h52;
  wire          compressDataVec_hitReq_28_82 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h52;
  wire          compressDataVec_hitReq_29_82 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h52;
  wire          compressDataVec_hitReq_30_82 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h52;
  wire          compressDataVec_hitReq_31_82 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h52;
  wire          compressDataVec_hitReq_32_82 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h52;
  wire          compressDataVec_hitReq_33_82 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h52;
  wire          compressDataVec_hitReq_34_82 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h52;
  wire          compressDataVec_hitReq_35_82 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h52;
  wire          compressDataVec_hitReq_36_82 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h52;
  wire          compressDataVec_hitReq_37_82 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h52;
  wire          compressDataVec_hitReq_38_82 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h52;
  wire          compressDataVec_hitReq_39_82 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h52;
  wire          compressDataVec_hitReq_40_82 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h52;
  wire          compressDataVec_hitReq_41_82 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h52;
  wire          compressDataVec_hitReq_42_82 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h52;
  wire          compressDataVec_hitReq_43_82 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h52;
  wire          compressDataVec_hitReq_44_82 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h52;
  wire          compressDataVec_hitReq_45_82 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h52;
  wire          compressDataVec_hitReq_46_82 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h52;
  wire          compressDataVec_hitReq_47_82 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h52;
  wire          compressDataVec_hitReq_48_82 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h52;
  wire          compressDataVec_hitReq_49_82 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h52;
  wire          compressDataVec_hitReq_50_82 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h52;
  wire          compressDataVec_hitReq_51_82 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h52;
  wire          compressDataVec_hitReq_52_82 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h52;
  wire          compressDataVec_hitReq_53_82 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h52;
  wire          compressDataVec_hitReq_54_82 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h52;
  wire          compressDataVec_hitReq_55_82 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h52;
  wire          compressDataVec_hitReq_56_82 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h52;
  wire          compressDataVec_hitReq_57_82 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h52;
  wire          compressDataVec_hitReq_58_82 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h52;
  wire          compressDataVec_hitReq_59_82 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h52;
  wire          compressDataVec_hitReq_60_82 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h52;
  wire          compressDataVec_hitReq_61_82 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h52;
  wire          compressDataVec_hitReq_62_82 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h52;
  wire          compressDataVec_hitReq_63_82 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h52;
  wire [7:0]    compressDataVec_selectReqData_82 =
    (compressDataVec_hitReq_0_82 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_82 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_82 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_82 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_82 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_82 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_82 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_82 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_82 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_82 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_82 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_82 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_82 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_82 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_82 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_82 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_82 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_82 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_82 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_82 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_82 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_82 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_82 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_82 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_82 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_82 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_82 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_82 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_82 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_82 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_82 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_82 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_82 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_82 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_82 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_82 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_82 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_82 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_82 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_82 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_82 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_82 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_82 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_82 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_82 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_82 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_82 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_82 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_82 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_82 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_82 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_82 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_82 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_82 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_82 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_82 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_82 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_82 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_82 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_82 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_82 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_82 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_82 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_82 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_83 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h53;
  wire          compressDataVec_hitReq_1_83 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h53;
  wire          compressDataVec_hitReq_2_83 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h53;
  wire          compressDataVec_hitReq_3_83 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h53;
  wire          compressDataVec_hitReq_4_83 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h53;
  wire          compressDataVec_hitReq_5_83 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h53;
  wire          compressDataVec_hitReq_6_83 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h53;
  wire          compressDataVec_hitReq_7_83 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h53;
  wire          compressDataVec_hitReq_8_83 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h53;
  wire          compressDataVec_hitReq_9_83 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h53;
  wire          compressDataVec_hitReq_10_83 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h53;
  wire          compressDataVec_hitReq_11_83 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h53;
  wire          compressDataVec_hitReq_12_83 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h53;
  wire          compressDataVec_hitReq_13_83 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h53;
  wire          compressDataVec_hitReq_14_83 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h53;
  wire          compressDataVec_hitReq_15_83 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h53;
  wire          compressDataVec_hitReq_16_83 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h53;
  wire          compressDataVec_hitReq_17_83 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h53;
  wire          compressDataVec_hitReq_18_83 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h53;
  wire          compressDataVec_hitReq_19_83 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h53;
  wire          compressDataVec_hitReq_20_83 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h53;
  wire          compressDataVec_hitReq_21_83 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h53;
  wire          compressDataVec_hitReq_22_83 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h53;
  wire          compressDataVec_hitReq_23_83 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h53;
  wire          compressDataVec_hitReq_24_83 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h53;
  wire          compressDataVec_hitReq_25_83 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h53;
  wire          compressDataVec_hitReq_26_83 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h53;
  wire          compressDataVec_hitReq_27_83 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h53;
  wire          compressDataVec_hitReq_28_83 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h53;
  wire          compressDataVec_hitReq_29_83 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h53;
  wire          compressDataVec_hitReq_30_83 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h53;
  wire          compressDataVec_hitReq_31_83 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h53;
  wire          compressDataVec_hitReq_32_83 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h53;
  wire          compressDataVec_hitReq_33_83 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h53;
  wire          compressDataVec_hitReq_34_83 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h53;
  wire          compressDataVec_hitReq_35_83 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h53;
  wire          compressDataVec_hitReq_36_83 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h53;
  wire          compressDataVec_hitReq_37_83 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h53;
  wire          compressDataVec_hitReq_38_83 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h53;
  wire          compressDataVec_hitReq_39_83 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h53;
  wire          compressDataVec_hitReq_40_83 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h53;
  wire          compressDataVec_hitReq_41_83 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h53;
  wire          compressDataVec_hitReq_42_83 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h53;
  wire          compressDataVec_hitReq_43_83 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h53;
  wire          compressDataVec_hitReq_44_83 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h53;
  wire          compressDataVec_hitReq_45_83 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h53;
  wire          compressDataVec_hitReq_46_83 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h53;
  wire          compressDataVec_hitReq_47_83 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h53;
  wire          compressDataVec_hitReq_48_83 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h53;
  wire          compressDataVec_hitReq_49_83 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h53;
  wire          compressDataVec_hitReq_50_83 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h53;
  wire          compressDataVec_hitReq_51_83 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h53;
  wire          compressDataVec_hitReq_52_83 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h53;
  wire          compressDataVec_hitReq_53_83 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h53;
  wire          compressDataVec_hitReq_54_83 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h53;
  wire          compressDataVec_hitReq_55_83 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h53;
  wire          compressDataVec_hitReq_56_83 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h53;
  wire          compressDataVec_hitReq_57_83 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h53;
  wire          compressDataVec_hitReq_58_83 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h53;
  wire          compressDataVec_hitReq_59_83 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h53;
  wire          compressDataVec_hitReq_60_83 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h53;
  wire          compressDataVec_hitReq_61_83 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h53;
  wire          compressDataVec_hitReq_62_83 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h53;
  wire          compressDataVec_hitReq_63_83 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h53;
  wire [7:0]    compressDataVec_selectReqData_83 =
    (compressDataVec_hitReq_0_83 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_83 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_83 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_83 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_83 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_83 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_83 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_83 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_83 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_83 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_83 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_83 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_83 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_83 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_83 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_83 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_83 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_83 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_83 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_83 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_83 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_83 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_83 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_83 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_83 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_83 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_83 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_83 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_83 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_83 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_83 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_83 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_83 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_83 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_83 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_83 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_83 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_83 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_83 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_83 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_83 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_83 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_83 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_83 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_83 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_83 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_83 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_83 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_83 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_83 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_83 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_83 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_83 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_83 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_83 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_83 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_83 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_83 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_83 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_83 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_83 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_83 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_83 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_83 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_84 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h54;
  wire          compressDataVec_hitReq_1_84 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h54;
  wire          compressDataVec_hitReq_2_84 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h54;
  wire          compressDataVec_hitReq_3_84 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h54;
  wire          compressDataVec_hitReq_4_84 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h54;
  wire          compressDataVec_hitReq_5_84 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h54;
  wire          compressDataVec_hitReq_6_84 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h54;
  wire          compressDataVec_hitReq_7_84 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h54;
  wire          compressDataVec_hitReq_8_84 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h54;
  wire          compressDataVec_hitReq_9_84 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h54;
  wire          compressDataVec_hitReq_10_84 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h54;
  wire          compressDataVec_hitReq_11_84 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h54;
  wire          compressDataVec_hitReq_12_84 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h54;
  wire          compressDataVec_hitReq_13_84 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h54;
  wire          compressDataVec_hitReq_14_84 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h54;
  wire          compressDataVec_hitReq_15_84 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h54;
  wire          compressDataVec_hitReq_16_84 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h54;
  wire          compressDataVec_hitReq_17_84 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h54;
  wire          compressDataVec_hitReq_18_84 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h54;
  wire          compressDataVec_hitReq_19_84 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h54;
  wire          compressDataVec_hitReq_20_84 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h54;
  wire          compressDataVec_hitReq_21_84 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h54;
  wire          compressDataVec_hitReq_22_84 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h54;
  wire          compressDataVec_hitReq_23_84 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h54;
  wire          compressDataVec_hitReq_24_84 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h54;
  wire          compressDataVec_hitReq_25_84 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h54;
  wire          compressDataVec_hitReq_26_84 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h54;
  wire          compressDataVec_hitReq_27_84 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h54;
  wire          compressDataVec_hitReq_28_84 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h54;
  wire          compressDataVec_hitReq_29_84 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h54;
  wire          compressDataVec_hitReq_30_84 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h54;
  wire          compressDataVec_hitReq_31_84 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h54;
  wire          compressDataVec_hitReq_32_84 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h54;
  wire          compressDataVec_hitReq_33_84 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h54;
  wire          compressDataVec_hitReq_34_84 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h54;
  wire          compressDataVec_hitReq_35_84 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h54;
  wire          compressDataVec_hitReq_36_84 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h54;
  wire          compressDataVec_hitReq_37_84 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h54;
  wire          compressDataVec_hitReq_38_84 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h54;
  wire          compressDataVec_hitReq_39_84 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h54;
  wire          compressDataVec_hitReq_40_84 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h54;
  wire          compressDataVec_hitReq_41_84 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h54;
  wire          compressDataVec_hitReq_42_84 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h54;
  wire          compressDataVec_hitReq_43_84 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h54;
  wire          compressDataVec_hitReq_44_84 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h54;
  wire          compressDataVec_hitReq_45_84 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h54;
  wire          compressDataVec_hitReq_46_84 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h54;
  wire          compressDataVec_hitReq_47_84 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h54;
  wire          compressDataVec_hitReq_48_84 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h54;
  wire          compressDataVec_hitReq_49_84 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h54;
  wire          compressDataVec_hitReq_50_84 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h54;
  wire          compressDataVec_hitReq_51_84 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h54;
  wire          compressDataVec_hitReq_52_84 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h54;
  wire          compressDataVec_hitReq_53_84 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h54;
  wire          compressDataVec_hitReq_54_84 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h54;
  wire          compressDataVec_hitReq_55_84 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h54;
  wire          compressDataVec_hitReq_56_84 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h54;
  wire          compressDataVec_hitReq_57_84 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h54;
  wire          compressDataVec_hitReq_58_84 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h54;
  wire          compressDataVec_hitReq_59_84 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h54;
  wire          compressDataVec_hitReq_60_84 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h54;
  wire          compressDataVec_hitReq_61_84 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h54;
  wire          compressDataVec_hitReq_62_84 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h54;
  wire          compressDataVec_hitReq_63_84 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h54;
  wire [7:0]    compressDataVec_selectReqData_84 =
    (compressDataVec_hitReq_0_84 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_84 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_84 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_84 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_84 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_84 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_84 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_84 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_84 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_84 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_84 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_84 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_84 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_84 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_84 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_84 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_84 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_84 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_84 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_84 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_84 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_84 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_84 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_84 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_84 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_84 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_84 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_84 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_84 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_84 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_84 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_84 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_84 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_84 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_84 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_84 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_84 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_84 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_84 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_84 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_84 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_84 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_84 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_84 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_84 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_84 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_84 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_84 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_84 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_84 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_84 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_84 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_84 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_84 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_84 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_84 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_84 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_84 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_84 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_84 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_84 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_84 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_84 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_84 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_85 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h55;
  wire          compressDataVec_hitReq_1_85 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h55;
  wire          compressDataVec_hitReq_2_85 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h55;
  wire          compressDataVec_hitReq_3_85 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h55;
  wire          compressDataVec_hitReq_4_85 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h55;
  wire          compressDataVec_hitReq_5_85 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h55;
  wire          compressDataVec_hitReq_6_85 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h55;
  wire          compressDataVec_hitReq_7_85 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h55;
  wire          compressDataVec_hitReq_8_85 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h55;
  wire          compressDataVec_hitReq_9_85 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h55;
  wire          compressDataVec_hitReq_10_85 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h55;
  wire          compressDataVec_hitReq_11_85 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h55;
  wire          compressDataVec_hitReq_12_85 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h55;
  wire          compressDataVec_hitReq_13_85 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h55;
  wire          compressDataVec_hitReq_14_85 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h55;
  wire          compressDataVec_hitReq_15_85 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h55;
  wire          compressDataVec_hitReq_16_85 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h55;
  wire          compressDataVec_hitReq_17_85 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h55;
  wire          compressDataVec_hitReq_18_85 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h55;
  wire          compressDataVec_hitReq_19_85 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h55;
  wire          compressDataVec_hitReq_20_85 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h55;
  wire          compressDataVec_hitReq_21_85 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h55;
  wire          compressDataVec_hitReq_22_85 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h55;
  wire          compressDataVec_hitReq_23_85 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h55;
  wire          compressDataVec_hitReq_24_85 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h55;
  wire          compressDataVec_hitReq_25_85 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h55;
  wire          compressDataVec_hitReq_26_85 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h55;
  wire          compressDataVec_hitReq_27_85 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h55;
  wire          compressDataVec_hitReq_28_85 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h55;
  wire          compressDataVec_hitReq_29_85 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h55;
  wire          compressDataVec_hitReq_30_85 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h55;
  wire          compressDataVec_hitReq_31_85 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h55;
  wire          compressDataVec_hitReq_32_85 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h55;
  wire          compressDataVec_hitReq_33_85 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h55;
  wire          compressDataVec_hitReq_34_85 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h55;
  wire          compressDataVec_hitReq_35_85 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h55;
  wire          compressDataVec_hitReq_36_85 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h55;
  wire          compressDataVec_hitReq_37_85 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h55;
  wire          compressDataVec_hitReq_38_85 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h55;
  wire          compressDataVec_hitReq_39_85 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h55;
  wire          compressDataVec_hitReq_40_85 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h55;
  wire          compressDataVec_hitReq_41_85 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h55;
  wire          compressDataVec_hitReq_42_85 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h55;
  wire          compressDataVec_hitReq_43_85 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h55;
  wire          compressDataVec_hitReq_44_85 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h55;
  wire          compressDataVec_hitReq_45_85 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h55;
  wire          compressDataVec_hitReq_46_85 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h55;
  wire          compressDataVec_hitReq_47_85 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h55;
  wire          compressDataVec_hitReq_48_85 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h55;
  wire          compressDataVec_hitReq_49_85 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h55;
  wire          compressDataVec_hitReq_50_85 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h55;
  wire          compressDataVec_hitReq_51_85 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h55;
  wire          compressDataVec_hitReq_52_85 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h55;
  wire          compressDataVec_hitReq_53_85 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h55;
  wire          compressDataVec_hitReq_54_85 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h55;
  wire          compressDataVec_hitReq_55_85 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h55;
  wire          compressDataVec_hitReq_56_85 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h55;
  wire          compressDataVec_hitReq_57_85 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h55;
  wire          compressDataVec_hitReq_58_85 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h55;
  wire          compressDataVec_hitReq_59_85 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h55;
  wire          compressDataVec_hitReq_60_85 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h55;
  wire          compressDataVec_hitReq_61_85 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h55;
  wire          compressDataVec_hitReq_62_85 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h55;
  wire          compressDataVec_hitReq_63_85 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h55;
  wire [7:0]    compressDataVec_selectReqData_85 =
    (compressDataVec_hitReq_0_85 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_85 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_85 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_85 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_85 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_85 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_85 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_85 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_85 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_85 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_85 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_85 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_85 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_85 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_85 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_85 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_85 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_85 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_85 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_85 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_85 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_85 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_85 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_85 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_85 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_85 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_85 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_85 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_85 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_85 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_85 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_85 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_85 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_85 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_85 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_85 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_85 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_85 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_85 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_85 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_85 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_85 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_85 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_85 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_85 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_85 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_85 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_85 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_85 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_85 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_85 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_85 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_85 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_85 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_85 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_85 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_85 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_85 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_85 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_85 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_85 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_85 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_85 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_85 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_86 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h56;
  wire          compressDataVec_hitReq_1_86 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h56;
  wire          compressDataVec_hitReq_2_86 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h56;
  wire          compressDataVec_hitReq_3_86 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h56;
  wire          compressDataVec_hitReq_4_86 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h56;
  wire          compressDataVec_hitReq_5_86 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h56;
  wire          compressDataVec_hitReq_6_86 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h56;
  wire          compressDataVec_hitReq_7_86 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h56;
  wire          compressDataVec_hitReq_8_86 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h56;
  wire          compressDataVec_hitReq_9_86 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h56;
  wire          compressDataVec_hitReq_10_86 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h56;
  wire          compressDataVec_hitReq_11_86 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h56;
  wire          compressDataVec_hitReq_12_86 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h56;
  wire          compressDataVec_hitReq_13_86 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h56;
  wire          compressDataVec_hitReq_14_86 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h56;
  wire          compressDataVec_hitReq_15_86 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h56;
  wire          compressDataVec_hitReq_16_86 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h56;
  wire          compressDataVec_hitReq_17_86 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h56;
  wire          compressDataVec_hitReq_18_86 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h56;
  wire          compressDataVec_hitReq_19_86 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h56;
  wire          compressDataVec_hitReq_20_86 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h56;
  wire          compressDataVec_hitReq_21_86 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h56;
  wire          compressDataVec_hitReq_22_86 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h56;
  wire          compressDataVec_hitReq_23_86 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h56;
  wire          compressDataVec_hitReq_24_86 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h56;
  wire          compressDataVec_hitReq_25_86 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h56;
  wire          compressDataVec_hitReq_26_86 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h56;
  wire          compressDataVec_hitReq_27_86 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h56;
  wire          compressDataVec_hitReq_28_86 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h56;
  wire          compressDataVec_hitReq_29_86 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h56;
  wire          compressDataVec_hitReq_30_86 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h56;
  wire          compressDataVec_hitReq_31_86 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h56;
  wire          compressDataVec_hitReq_32_86 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h56;
  wire          compressDataVec_hitReq_33_86 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h56;
  wire          compressDataVec_hitReq_34_86 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h56;
  wire          compressDataVec_hitReq_35_86 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h56;
  wire          compressDataVec_hitReq_36_86 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h56;
  wire          compressDataVec_hitReq_37_86 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h56;
  wire          compressDataVec_hitReq_38_86 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h56;
  wire          compressDataVec_hitReq_39_86 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h56;
  wire          compressDataVec_hitReq_40_86 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h56;
  wire          compressDataVec_hitReq_41_86 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h56;
  wire          compressDataVec_hitReq_42_86 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h56;
  wire          compressDataVec_hitReq_43_86 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h56;
  wire          compressDataVec_hitReq_44_86 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h56;
  wire          compressDataVec_hitReq_45_86 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h56;
  wire          compressDataVec_hitReq_46_86 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h56;
  wire          compressDataVec_hitReq_47_86 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h56;
  wire          compressDataVec_hitReq_48_86 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h56;
  wire          compressDataVec_hitReq_49_86 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h56;
  wire          compressDataVec_hitReq_50_86 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h56;
  wire          compressDataVec_hitReq_51_86 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h56;
  wire          compressDataVec_hitReq_52_86 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h56;
  wire          compressDataVec_hitReq_53_86 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h56;
  wire          compressDataVec_hitReq_54_86 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h56;
  wire          compressDataVec_hitReq_55_86 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h56;
  wire          compressDataVec_hitReq_56_86 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h56;
  wire          compressDataVec_hitReq_57_86 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h56;
  wire          compressDataVec_hitReq_58_86 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h56;
  wire          compressDataVec_hitReq_59_86 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h56;
  wire          compressDataVec_hitReq_60_86 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h56;
  wire          compressDataVec_hitReq_61_86 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h56;
  wire          compressDataVec_hitReq_62_86 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h56;
  wire          compressDataVec_hitReq_63_86 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h56;
  wire [7:0]    compressDataVec_selectReqData_86 =
    (compressDataVec_hitReq_0_86 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_86 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_86 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_86 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_86 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_86 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_86 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_86 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_86 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_86 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_86 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_86 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_86 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_86 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_86 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_86 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_86 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_86 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_86 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_86 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_86 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_86 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_86 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_86 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_86 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_86 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_86 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_86 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_86 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_86 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_86 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_86 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_86 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_86 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_86 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_86 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_86 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_86 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_86 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_86 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_86 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_86 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_86 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_86 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_86 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_86 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_86 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_86 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_86 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_86 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_86 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_86 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_86 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_86 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_86 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_86 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_86 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_86 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_86 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_86 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_86 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_86 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_86 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_86 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_87 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h57;
  wire          compressDataVec_hitReq_1_87 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h57;
  wire          compressDataVec_hitReq_2_87 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h57;
  wire          compressDataVec_hitReq_3_87 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h57;
  wire          compressDataVec_hitReq_4_87 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h57;
  wire          compressDataVec_hitReq_5_87 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h57;
  wire          compressDataVec_hitReq_6_87 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h57;
  wire          compressDataVec_hitReq_7_87 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h57;
  wire          compressDataVec_hitReq_8_87 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h57;
  wire          compressDataVec_hitReq_9_87 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h57;
  wire          compressDataVec_hitReq_10_87 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h57;
  wire          compressDataVec_hitReq_11_87 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h57;
  wire          compressDataVec_hitReq_12_87 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h57;
  wire          compressDataVec_hitReq_13_87 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h57;
  wire          compressDataVec_hitReq_14_87 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h57;
  wire          compressDataVec_hitReq_15_87 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h57;
  wire          compressDataVec_hitReq_16_87 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h57;
  wire          compressDataVec_hitReq_17_87 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h57;
  wire          compressDataVec_hitReq_18_87 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h57;
  wire          compressDataVec_hitReq_19_87 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h57;
  wire          compressDataVec_hitReq_20_87 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h57;
  wire          compressDataVec_hitReq_21_87 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h57;
  wire          compressDataVec_hitReq_22_87 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h57;
  wire          compressDataVec_hitReq_23_87 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h57;
  wire          compressDataVec_hitReq_24_87 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h57;
  wire          compressDataVec_hitReq_25_87 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h57;
  wire          compressDataVec_hitReq_26_87 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h57;
  wire          compressDataVec_hitReq_27_87 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h57;
  wire          compressDataVec_hitReq_28_87 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h57;
  wire          compressDataVec_hitReq_29_87 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h57;
  wire          compressDataVec_hitReq_30_87 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h57;
  wire          compressDataVec_hitReq_31_87 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h57;
  wire          compressDataVec_hitReq_32_87 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h57;
  wire          compressDataVec_hitReq_33_87 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h57;
  wire          compressDataVec_hitReq_34_87 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h57;
  wire          compressDataVec_hitReq_35_87 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h57;
  wire          compressDataVec_hitReq_36_87 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h57;
  wire          compressDataVec_hitReq_37_87 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h57;
  wire          compressDataVec_hitReq_38_87 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h57;
  wire          compressDataVec_hitReq_39_87 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h57;
  wire          compressDataVec_hitReq_40_87 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h57;
  wire          compressDataVec_hitReq_41_87 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h57;
  wire          compressDataVec_hitReq_42_87 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h57;
  wire          compressDataVec_hitReq_43_87 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h57;
  wire          compressDataVec_hitReq_44_87 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h57;
  wire          compressDataVec_hitReq_45_87 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h57;
  wire          compressDataVec_hitReq_46_87 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h57;
  wire          compressDataVec_hitReq_47_87 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h57;
  wire          compressDataVec_hitReq_48_87 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h57;
  wire          compressDataVec_hitReq_49_87 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h57;
  wire          compressDataVec_hitReq_50_87 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h57;
  wire          compressDataVec_hitReq_51_87 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h57;
  wire          compressDataVec_hitReq_52_87 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h57;
  wire          compressDataVec_hitReq_53_87 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h57;
  wire          compressDataVec_hitReq_54_87 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h57;
  wire          compressDataVec_hitReq_55_87 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h57;
  wire          compressDataVec_hitReq_56_87 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h57;
  wire          compressDataVec_hitReq_57_87 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h57;
  wire          compressDataVec_hitReq_58_87 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h57;
  wire          compressDataVec_hitReq_59_87 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h57;
  wire          compressDataVec_hitReq_60_87 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h57;
  wire          compressDataVec_hitReq_61_87 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h57;
  wire          compressDataVec_hitReq_62_87 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h57;
  wire          compressDataVec_hitReq_63_87 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h57;
  wire [7:0]    compressDataVec_selectReqData_87 =
    (compressDataVec_hitReq_0_87 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_87 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_87 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_87 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_87 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_87 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_87 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_87 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_87 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_87 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_87 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_87 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_87 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_87 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_87 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_87 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_87 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_87 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_87 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_87 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_87 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_87 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_87 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_87 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_87 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_87 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_87 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_87 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_87 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_87 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_87 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_87 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_87 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_87 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_87 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_87 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_87 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_87 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_87 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_87 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_87 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_87 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_87 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_87 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_87 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_87 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_87 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_87 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_87 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_87 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_87 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_87 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_87 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_87 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_87 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_87 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_87 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_87 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_87 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_87 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_87 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_87 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_87 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_87 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_88 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h58;
  wire          compressDataVec_hitReq_1_88 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h58;
  wire          compressDataVec_hitReq_2_88 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h58;
  wire          compressDataVec_hitReq_3_88 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h58;
  wire          compressDataVec_hitReq_4_88 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h58;
  wire          compressDataVec_hitReq_5_88 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h58;
  wire          compressDataVec_hitReq_6_88 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h58;
  wire          compressDataVec_hitReq_7_88 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h58;
  wire          compressDataVec_hitReq_8_88 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h58;
  wire          compressDataVec_hitReq_9_88 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h58;
  wire          compressDataVec_hitReq_10_88 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h58;
  wire          compressDataVec_hitReq_11_88 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h58;
  wire          compressDataVec_hitReq_12_88 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h58;
  wire          compressDataVec_hitReq_13_88 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h58;
  wire          compressDataVec_hitReq_14_88 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h58;
  wire          compressDataVec_hitReq_15_88 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h58;
  wire          compressDataVec_hitReq_16_88 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h58;
  wire          compressDataVec_hitReq_17_88 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h58;
  wire          compressDataVec_hitReq_18_88 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h58;
  wire          compressDataVec_hitReq_19_88 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h58;
  wire          compressDataVec_hitReq_20_88 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h58;
  wire          compressDataVec_hitReq_21_88 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h58;
  wire          compressDataVec_hitReq_22_88 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h58;
  wire          compressDataVec_hitReq_23_88 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h58;
  wire          compressDataVec_hitReq_24_88 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h58;
  wire          compressDataVec_hitReq_25_88 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h58;
  wire          compressDataVec_hitReq_26_88 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h58;
  wire          compressDataVec_hitReq_27_88 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h58;
  wire          compressDataVec_hitReq_28_88 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h58;
  wire          compressDataVec_hitReq_29_88 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h58;
  wire          compressDataVec_hitReq_30_88 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h58;
  wire          compressDataVec_hitReq_31_88 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h58;
  wire          compressDataVec_hitReq_32_88 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h58;
  wire          compressDataVec_hitReq_33_88 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h58;
  wire          compressDataVec_hitReq_34_88 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h58;
  wire          compressDataVec_hitReq_35_88 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h58;
  wire          compressDataVec_hitReq_36_88 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h58;
  wire          compressDataVec_hitReq_37_88 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h58;
  wire          compressDataVec_hitReq_38_88 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h58;
  wire          compressDataVec_hitReq_39_88 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h58;
  wire          compressDataVec_hitReq_40_88 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h58;
  wire          compressDataVec_hitReq_41_88 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h58;
  wire          compressDataVec_hitReq_42_88 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h58;
  wire          compressDataVec_hitReq_43_88 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h58;
  wire          compressDataVec_hitReq_44_88 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h58;
  wire          compressDataVec_hitReq_45_88 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h58;
  wire          compressDataVec_hitReq_46_88 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h58;
  wire          compressDataVec_hitReq_47_88 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h58;
  wire          compressDataVec_hitReq_48_88 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h58;
  wire          compressDataVec_hitReq_49_88 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h58;
  wire          compressDataVec_hitReq_50_88 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h58;
  wire          compressDataVec_hitReq_51_88 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h58;
  wire          compressDataVec_hitReq_52_88 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h58;
  wire          compressDataVec_hitReq_53_88 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h58;
  wire          compressDataVec_hitReq_54_88 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h58;
  wire          compressDataVec_hitReq_55_88 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h58;
  wire          compressDataVec_hitReq_56_88 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h58;
  wire          compressDataVec_hitReq_57_88 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h58;
  wire          compressDataVec_hitReq_58_88 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h58;
  wire          compressDataVec_hitReq_59_88 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h58;
  wire          compressDataVec_hitReq_60_88 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h58;
  wire          compressDataVec_hitReq_61_88 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h58;
  wire          compressDataVec_hitReq_62_88 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h58;
  wire          compressDataVec_hitReq_63_88 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h58;
  wire [7:0]    compressDataVec_selectReqData_88 =
    (compressDataVec_hitReq_0_88 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_88 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_88 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_88 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_88 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_88 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_88 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_88 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_88 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_88 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_88 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_88 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_88 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_88 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_88 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_88 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_88 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_88 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_88 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_88 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_88 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_88 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_88 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_88 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_88 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_88 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_88 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_88 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_88 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_88 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_88 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_88 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_88 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_88 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_88 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_88 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_88 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_88 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_88 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_88 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_88 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_88 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_88 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_88 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_88 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_88 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_88 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_88 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_88 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_88 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_88 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_88 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_88 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_88 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_88 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_88 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_88 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_88 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_88 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_88 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_88 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_88 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_88 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_88 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_89 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h59;
  wire          compressDataVec_hitReq_1_89 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h59;
  wire          compressDataVec_hitReq_2_89 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h59;
  wire          compressDataVec_hitReq_3_89 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h59;
  wire          compressDataVec_hitReq_4_89 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h59;
  wire          compressDataVec_hitReq_5_89 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h59;
  wire          compressDataVec_hitReq_6_89 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h59;
  wire          compressDataVec_hitReq_7_89 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h59;
  wire          compressDataVec_hitReq_8_89 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h59;
  wire          compressDataVec_hitReq_9_89 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h59;
  wire          compressDataVec_hitReq_10_89 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h59;
  wire          compressDataVec_hitReq_11_89 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h59;
  wire          compressDataVec_hitReq_12_89 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h59;
  wire          compressDataVec_hitReq_13_89 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h59;
  wire          compressDataVec_hitReq_14_89 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h59;
  wire          compressDataVec_hitReq_15_89 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h59;
  wire          compressDataVec_hitReq_16_89 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h59;
  wire          compressDataVec_hitReq_17_89 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h59;
  wire          compressDataVec_hitReq_18_89 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h59;
  wire          compressDataVec_hitReq_19_89 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h59;
  wire          compressDataVec_hitReq_20_89 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h59;
  wire          compressDataVec_hitReq_21_89 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h59;
  wire          compressDataVec_hitReq_22_89 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h59;
  wire          compressDataVec_hitReq_23_89 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h59;
  wire          compressDataVec_hitReq_24_89 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h59;
  wire          compressDataVec_hitReq_25_89 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h59;
  wire          compressDataVec_hitReq_26_89 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h59;
  wire          compressDataVec_hitReq_27_89 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h59;
  wire          compressDataVec_hitReq_28_89 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h59;
  wire          compressDataVec_hitReq_29_89 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h59;
  wire          compressDataVec_hitReq_30_89 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h59;
  wire          compressDataVec_hitReq_31_89 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h59;
  wire          compressDataVec_hitReq_32_89 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h59;
  wire          compressDataVec_hitReq_33_89 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h59;
  wire          compressDataVec_hitReq_34_89 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h59;
  wire          compressDataVec_hitReq_35_89 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h59;
  wire          compressDataVec_hitReq_36_89 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h59;
  wire          compressDataVec_hitReq_37_89 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h59;
  wire          compressDataVec_hitReq_38_89 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h59;
  wire          compressDataVec_hitReq_39_89 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h59;
  wire          compressDataVec_hitReq_40_89 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h59;
  wire          compressDataVec_hitReq_41_89 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h59;
  wire          compressDataVec_hitReq_42_89 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h59;
  wire          compressDataVec_hitReq_43_89 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h59;
  wire          compressDataVec_hitReq_44_89 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h59;
  wire          compressDataVec_hitReq_45_89 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h59;
  wire          compressDataVec_hitReq_46_89 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h59;
  wire          compressDataVec_hitReq_47_89 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h59;
  wire          compressDataVec_hitReq_48_89 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h59;
  wire          compressDataVec_hitReq_49_89 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h59;
  wire          compressDataVec_hitReq_50_89 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h59;
  wire          compressDataVec_hitReq_51_89 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h59;
  wire          compressDataVec_hitReq_52_89 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h59;
  wire          compressDataVec_hitReq_53_89 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h59;
  wire          compressDataVec_hitReq_54_89 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h59;
  wire          compressDataVec_hitReq_55_89 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h59;
  wire          compressDataVec_hitReq_56_89 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h59;
  wire          compressDataVec_hitReq_57_89 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h59;
  wire          compressDataVec_hitReq_58_89 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h59;
  wire          compressDataVec_hitReq_59_89 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h59;
  wire          compressDataVec_hitReq_60_89 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h59;
  wire          compressDataVec_hitReq_61_89 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h59;
  wire          compressDataVec_hitReq_62_89 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h59;
  wire          compressDataVec_hitReq_63_89 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h59;
  wire [7:0]    compressDataVec_selectReqData_89 =
    (compressDataVec_hitReq_0_89 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_89 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_89 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_89 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_89 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_89 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_89 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_89 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_89 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_89 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_89 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_89 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_89 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_89 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_89 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_89 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_89 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_89 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_89 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_89 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_89 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_89 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_89 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_89 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_89 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_89 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_89 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_89 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_89 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_89 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_89 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_89 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_89 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_89 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_89 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_89 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_89 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_89 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_89 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_89 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_89 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_89 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_89 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_89 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_89 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_89 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_89 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_89 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_89 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_89 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_89 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_89 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_89 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_89 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_89 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_89 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_89 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_89 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_89 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_89 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_89 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_89 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_89 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_89 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_90 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h5A;
  wire          compressDataVec_hitReq_1_90 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h5A;
  wire          compressDataVec_hitReq_2_90 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h5A;
  wire          compressDataVec_hitReq_3_90 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h5A;
  wire          compressDataVec_hitReq_4_90 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h5A;
  wire          compressDataVec_hitReq_5_90 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h5A;
  wire          compressDataVec_hitReq_6_90 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h5A;
  wire          compressDataVec_hitReq_7_90 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h5A;
  wire          compressDataVec_hitReq_8_90 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h5A;
  wire          compressDataVec_hitReq_9_90 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h5A;
  wire          compressDataVec_hitReq_10_90 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h5A;
  wire          compressDataVec_hitReq_11_90 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h5A;
  wire          compressDataVec_hitReq_12_90 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h5A;
  wire          compressDataVec_hitReq_13_90 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h5A;
  wire          compressDataVec_hitReq_14_90 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h5A;
  wire          compressDataVec_hitReq_15_90 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h5A;
  wire          compressDataVec_hitReq_16_90 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h5A;
  wire          compressDataVec_hitReq_17_90 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h5A;
  wire          compressDataVec_hitReq_18_90 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h5A;
  wire          compressDataVec_hitReq_19_90 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h5A;
  wire          compressDataVec_hitReq_20_90 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h5A;
  wire          compressDataVec_hitReq_21_90 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h5A;
  wire          compressDataVec_hitReq_22_90 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h5A;
  wire          compressDataVec_hitReq_23_90 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h5A;
  wire          compressDataVec_hitReq_24_90 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h5A;
  wire          compressDataVec_hitReq_25_90 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h5A;
  wire          compressDataVec_hitReq_26_90 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h5A;
  wire          compressDataVec_hitReq_27_90 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h5A;
  wire          compressDataVec_hitReq_28_90 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h5A;
  wire          compressDataVec_hitReq_29_90 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h5A;
  wire          compressDataVec_hitReq_30_90 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h5A;
  wire          compressDataVec_hitReq_31_90 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h5A;
  wire          compressDataVec_hitReq_32_90 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h5A;
  wire          compressDataVec_hitReq_33_90 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h5A;
  wire          compressDataVec_hitReq_34_90 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h5A;
  wire          compressDataVec_hitReq_35_90 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h5A;
  wire          compressDataVec_hitReq_36_90 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h5A;
  wire          compressDataVec_hitReq_37_90 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h5A;
  wire          compressDataVec_hitReq_38_90 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h5A;
  wire          compressDataVec_hitReq_39_90 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h5A;
  wire          compressDataVec_hitReq_40_90 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h5A;
  wire          compressDataVec_hitReq_41_90 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h5A;
  wire          compressDataVec_hitReq_42_90 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h5A;
  wire          compressDataVec_hitReq_43_90 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h5A;
  wire          compressDataVec_hitReq_44_90 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h5A;
  wire          compressDataVec_hitReq_45_90 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h5A;
  wire          compressDataVec_hitReq_46_90 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h5A;
  wire          compressDataVec_hitReq_47_90 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h5A;
  wire          compressDataVec_hitReq_48_90 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h5A;
  wire          compressDataVec_hitReq_49_90 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h5A;
  wire          compressDataVec_hitReq_50_90 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h5A;
  wire          compressDataVec_hitReq_51_90 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h5A;
  wire          compressDataVec_hitReq_52_90 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h5A;
  wire          compressDataVec_hitReq_53_90 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h5A;
  wire          compressDataVec_hitReq_54_90 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h5A;
  wire          compressDataVec_hitReq_55_90 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h5A;
  wire          compressDataVec_hitReq_56_90 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h5A;
  wire          compressDataVec_hitReq_57_90 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h5A;
  wire          compressDataVec_hitReq_58_90 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h5A;
  wire          compressDataVec_hitReq_59_90 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h5A;
  wire          compressDataVec_hitReq_60_90 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h5A;
  wire          compressDataVec_hitReq_61_90 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h5A;
  wire          compressDataVec_hitReq_62_90 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h5A;
  wire          compressDataVec_hitReq_63_90 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h5A;
  wire [7:0]    compressDataVec_selectReqData_90 =
    (compressDataVec_hitReq_0_90 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_90 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_90 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_90 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_90 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_90 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_90 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_90 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_90 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_90 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_90 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_90 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_90 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_90 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_90 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_90 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_90 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_90 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_90 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_90 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_90 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_90 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_90 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_90 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_90 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_90 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_90 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_90 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_90 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_90 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_90 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_90 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_90 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_90 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_90 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_90 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_90 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_90 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_90 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_90 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_90 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_90 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_90 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_90 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_90 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_90 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_90 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_90 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_90 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_90 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_90 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_90 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_90 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_90 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_90 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_90 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_90 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_90 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_90 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_90 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_90 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_90 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_90 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_90 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_91 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h5B;
  wire          compressDataVec_hitReq_1_91 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h5B;
  wire          compressDataVec_hitReq_2_91 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h5B;
  wire          compressDataVec_hitReq_3_91 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h5B;
  wire          compressDataVec_hitReq_4_91 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h5B;
  wire          compressDataVec_hitReq_5_91 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h5B;
  wire          compressDataVec_hitReq_6_91 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h5B;
  wire          compressDataVec_hitReq_7_91 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h5B;
  wire          compressDataVec_hitReq_8_91 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h5B;
  wire          compressDataVec_hitReq_9_91 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h5B;
  wire          compressDataVec_hitReq_10_91 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h5B;
  wire          compressDataVec_hitReq_11_91 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h5B;
  wire          compressDataVec_hitReq_12_91 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h5B;
  wire          compressDataVec_hitReq_13_91 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h5B;
  wire          compressDataVec_hitReq_14_91 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h5B;
  wire          compressDataVec_hitReq_15_91 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h5B;
  wire          compressDataVec_hitReq_16_91 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h5B;
  wire          compressDataVec_hitReq_17_91 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h5B;
  wire          compressDataVec_hitReq_18_91 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h5B;
  wire          compressDataVec_hitReq_19_91 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h5B;
  wire          compressDataVec_hitReq_20_91 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h5B;
  wire          compressDataVec_hitReq_21_91 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h5B;
  wire          compressDataVec_hitReq_22_91 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h5B;
  wire          compressDataVec_hitReq_23_91 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h5B;
  wire          compressDataVec_hitReq_24_91 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h5B;
  wire          compressDataVec_hitReq_25_91 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h5B;
  wire          compressDataVec_hitReq_26_91 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h5B;
  wire          compressDataVec_hitReq_27_91 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h5B;
  wire          compressDataVec_hitReq_28_91 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h5B;
  wire          compressDataVec_hitReq_29_91 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h5B;
  wire          compressDataVec_hitReq_30_91 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h5B;
  wire          compressDataVec_hitReq_31_91 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h5B;
  wire          compressDataVec_hitReq_32_91 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h5B;
  wire          compressDataVec_hitReq_33_91 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h5B;
  wire          compressDataVec_hitReq_34_91 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h5B;
  wire          compressDataVec_hitReq_35_91 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h5B;
  wire          compressDataVec_hitReq_36_91 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h5B;
  wire          compressDataVec_hitReq_37_91 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h5B;
  wire          compressDataVec_hitReq_38_91 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h5B;
  wire          compressDataVec_hitReq_39_91 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h5B;
  wire          compressDataVec_hitReq_40_91 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h5B;
  wire          compressDataVec_hitReq_41_91 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h5B;
  wire          compressDataVec_hitReq_42_91 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h5B;
  wire          compressDataVec_hitReq_43_91 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h5B;
  wire          compressDataVec_hitReq_44_91 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h5B;
  wire          compressDataVec_hitReq_45_91 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h5B;
  wire          compressDataVec_hitReq_46_91 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h5B;
  wire          compressDataVec_hitReq_47_91 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h5B;
  wire          compressDataVec_hitReq_48_91 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h5B;
  wire          compressDataVec_hitReq_49_91 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h5B;
  wire          compressDataVec_hitReq_50_91 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h5B;
  wire          compressDataVec_hitReq_51_91 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h5B;
  wire          compressDataVec_hitReq_52_91 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h5B;
  wire          compressDataVec_hitReq_53_91 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h5B;
  wire          compressDataVec_hitReq_54_91 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h5B;
  wire          compressDataVec_hitReq_55_91 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h5B;
  wire          compressDataVec_hitReq_56_91 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h5B;
  wire          compressDataVec_hitReq_57_91 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h5B;
  wire          compressDataVec_hitReq_58_91 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h5B;
  wire          compressDataVec_hitReq_59_91 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h5B;
  wire          compressDataVec_hitReq_60_91 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h5B;
  wire          compressDataVec_hitReq_61_91 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h5B;
  wire          compressDataVec_hitReq_62_91 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h5B;
  wire          compressDataVec_hitReq_63_91 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h5B;
  wire [7:0]    compressDataVec_selectReqData_91 =
    (compressDataVec_hitReq_0_91 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_91 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_91 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_91 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_91 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_91 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_91 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_91 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_91 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_91 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_91 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_91 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_91 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_91 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_91 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_91 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_91 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_91 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_91 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_91 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_91 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_91 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_91 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_91 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_91 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_91 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_91 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_91 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_91 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_91 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_91 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_91 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_91 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_91 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_91 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_91 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_91 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_91 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_91 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_91 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_91 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_91 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_91 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_91 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_91 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_91 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_91 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_91 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_91 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_91 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_91 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_91 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_91 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_91 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_91 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_91 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_91 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_91 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_91 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_91 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_91 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_91 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_91 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_91 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_92 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h5C;
  wire          compressDataVec_hitReq_1_92 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h5C;
  wire          compressDataVec_hitReq_2_92 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h5C;
  wire          compressDataVec_hitReq_3_92 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h5C;
  wire          compressDataVec_hitReq_4_92 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h5C;
  wire          compressDataVec_hitReq_5_92 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h5C;
  wire          compressDataVec_hitReq_6_92 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h5C;
  wire          compressDataVec_hitReq_7_92 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h5C;
  wire          compressDataVec_hitReq_8_92 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h5C;
  wire          compressDataVec_hitReq_9_92 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h5C;
  wire          compressDataVec_hitReq_10_92 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h5C;
  wire          compressDataVec_hitReq_11_92 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h5C;
  wire          compressDataVec_hitReq_12_92 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h5C;
  wire          compressDataVec_hitReq_13_92 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h5C;
  wire          compressDataVec_hitReq_14_92 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h5C;
  wire          compressDataVec_hitReq_15_92 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h5C;
  wire          compressDataVec_hitReq_16_92 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h5C;
  wire          compressDataVec_hitReq_17_92 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h5C;
  wire          compressDataVec_hitReq_18_92 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h5C;
  wire          compressDataVec_hitReq_19_92 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h5C;
  wire          compressDataVec_hitReq_20_92 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h5C;
  wire          compressDataVec_hitReq_21_92 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h5C;
  wire          compressDataVec_hitReq_22_92 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h5C;
  wire          compressDataVec_hitReq_23_92 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h5C;
  wire          compressDataVec_hitReq_24_92 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h5C;
  wire          compressDataVec_hitReq_25_92 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h5C;
  wire          compressDataVec_hitReq_26_92 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h5C;
  wire          compressDataVec_hitReq_27_92 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h5C;
  wire          compressDataVec_hitReq_28_92 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h5C;
  wire          compressDataVec_hitReq_29_92 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h5C;
  wire          compressDataVec_hitReq_30_92 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h5C;
  wire          compressDataVec_hitReq_31_92 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h5C;
  wire          compressDataVec_hitReq_32_92 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h5C;
  wire          compressDataVec_hitReq_33_92 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h5C;
  wire          compressDataVec_hitReq_34_92 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h5C;
  wire          compressDataVec_hitReq_35_92 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h5C;
  wire          compressDataVec_hitReq_36_92 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h5C;
  wire          compressDataVec_hitReq_37_92 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h5C;
  wire          compressDataVec_hitReq_38_92 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h5C;
  wire          compressDataVec_hitReq_39_92 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h5C;
  wire          compressDataVec_hitReq_40_92 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h5C;
  wire          compressDataVec_hitReq_41_92 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h5C;
  wire          compressDataVec_hitReq_42_92 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h5C;
  wire          compressDataVec_hitReq_43_92 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h5C;
  wire          compressDataVec_hitReq_44_92 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h5C;
  wire          compressDataVec_hitReq_45_92 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h5C;
  wire          compressDataVec_hitReq_46_92 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h5C;
  wire          compressDataVec_hitReq_47_92 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h5C;
  wire          compressDataVec_hitReq_48_92 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h5C;
  wire          compressDataVec_hitReq_49_92 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h5C;
  wire          compressDataVec_hitReq_50_92 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h5C;
  wire          compressDataVec_hitReq_51_92 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h5C;
  wire          compressDataVec_hitReq_52_92 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h5C;
  wire          compressDataVec_hitReq_53_92 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h5C;
  wire          compressDataVec_hitReq_54_92 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h5C;
  wire          compressDataVec_hitReq_55_92 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h5C;
  wire          compressDataVec_hitReq_56_92 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h5C;
  wire          compressDataVec_hitReq_57_92 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h5C;
  wire          compressDataVec_hitReq_58_92 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h5C;
  wire          compressDataVec_hitReq_59_92 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h5C;
  wire          compressDataVec_hitReq_60_92 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h5C;
  wire          compressDataVec_hitReq_61_92 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h5C;
  wire          compressDataVec_hitReq_62_92 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h5C;
  wire          compressDataVec_hitReq_63_92 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h5C;
  wire [7:0]    compressDataVec_selectReqData_92 =
    (compressDataVec_hitReq_0_92 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_92 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_92 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_92 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_92 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_92 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_92 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_92 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_92 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_92 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_92 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_92 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_92 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_92 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_92 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_92 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_92 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_92 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_92 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_92 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_92 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_92 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_92 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_92 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_92 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_92 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_92 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_92 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_92 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_92 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_92 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_92 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_92 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_92 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_92 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_92 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_92 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_92 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_92 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_92 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_92 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_92 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_92 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_92 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_92 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_92 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_92 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_92 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_92 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_92 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_92 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_92 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_92 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_92 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_92 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_92 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_92 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_92 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_92 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_92 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_92 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_92 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_92 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_92 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_93 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h5D;
  wire          compressDataVec_hitReq_1_93 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h5D;
  wire          compressDataVec_hitReq_2_93 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h5D;
  wire          compressDataVec_hitReq_3_93 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h5D;
  wire          compressDataVec_hitReq_4_93 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h5D;
  wire          compressDataVec_hitReq_5_93 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h5D;
  wire          compressDataVec_hitReq_6_93 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h5D;
  wire          compressDataVec_hitReq_7_93 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h5D;
  wire          compressDataVec_hitReq_8_93 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h5D;
  wire          compressDataVec_hitReq_9_93 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h5D;
  wire          compressDataVec_hitReq_10_93 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h5D;
  wire          compressDataVec_hitReq_11_93 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h5D;
  wire          compressDataVec_hitReq_12_93 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h5D;
  wire          compressDataVec_hitReq_13_93 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h5D;
  wire          compressDataVec_hitReq_14_93 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h5D;
  wire          compressDataVec_hitReq_15_93 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h5D;
  wire          compressDataVec_hitReq_16_93 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h5D;
  wire          compressDataVec_hitReq_17_93 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h5D;
  wire          compressDataVec_hitReq_18_93 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h5D;
  wire          compressDataVec_hitReq_19_93 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h5D;
  wire          compressDataVec_hitReq_20_93 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h5D;
  wire          compressDataVec_hitReq_21_93 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h5D;
  wire          compressDataVec_hitReq_22_93 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h5D;
  wire          compressDataVec_hitReq_23_93 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h5D;
  wire          compressDataVec_hitReq_24_93 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h5D;
  wire          compressDataVec_hitReq_25_93 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h5D;
  wire          compressDataVec_hitReq_26_93 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h5D;
  wire          compressDataVec_hitReq_27_93 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h5D;
  wire          compressDataVec_hitReq_28_93 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h5D;
  wire          compressDataVec_hitReq_29_93 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h5D;
  wire          compressDataVec_hitReq_30_93 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h5D;
  wire          compressDataVec_hitReq_31_93 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h5D;
  wire          compressDataVec_hitReq_32_93 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h5D;
  wire          compressDataVec_hitReq_33_93 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h5D;
  wire          compressDataVec_hitReq_34_93 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h5D;
  wire          compressDataVec_hitReq_35_93 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h5D;
  wire          compressDataVec_hitReq_36_93 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h5D;
  wire          compressDataVec_hitReq_37_93 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h5D;
  wire          compressDataVec_hitReq_38_93 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h5D;
  wire          compressDataVec_hitReq_39_93 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h5D;
  wire          compressDataVec_hitReq_40_93 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h5D;
  wire          compressDataVec_hitReq_41_93 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h5D;
  wire          compressDataVec_hitReq_42_93 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h5D;
  wire          compressDataVec_hitReq_43_93 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h5D;
  wire          compressDataVec_hitReq_44_93 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h5D;
  wire          compressDataVec_hitReq_45_93 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h5D;
  wire          compressDataVec_hitReq_46_93 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h5D;
  wire          compressDataVec_hitReq_47_93 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h5D;
  wire          compressDataVec_hitReq_48_93 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h5D;
  wire          compressDataVec_hitReq_49_93 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h5D;
  wire          compressDataVec_hitReq_50_93 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h5D;
  wire          compressDataVec_hitReq_51_93 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h5D;
  wire          compressDataVec_hitReq_52_93 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h5D;
  wire          compressDataVec_hitReq_53_93 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h5D;
  wire          compressDataVec_hitReq_54_93 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h5D;
  wire          compressDataVec_hitReq_55_93 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h5D;
  wire          compressDataVec_hitReq_56_93 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h5D;
  wire          compressDataVec_hitReq_57_93 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h5D;
  wire          compressDataVec_hitReq_58_93 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h5D;
  wire          compressDataVec_hitReq_59_93 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h5D;
  wire          compressDataVec_hitReq_60_93 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h5D;
  wire          compressDataVec_hitReq_61_93 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h5D;
  wire          compressDataVec_hitReq_62_93 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h5D;
  wire          compressDataVec_hitReq_63_93 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h5D;
  wire [7:0]    compressDataVec_selectReqData_93 =
    (compressDataVec_hitReq_0_93 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_93 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_93 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_93 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_93 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_93 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_93 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_93 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_93 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_93 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_93 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_93 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_93 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_93 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_93 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_93 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_93 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_93 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_93 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_93 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_93 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_93 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_93 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_93 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_93 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_93 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_93 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_93 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_93 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_93 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_93 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_93 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_93 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_93 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_93 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_93 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_93 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_93 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_93 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_93 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_93 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_93 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_93 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_93 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_93 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_93 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_93 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_93 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_93 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_93 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_93 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_93 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_93 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_93 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_93 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_93 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_93 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_93 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_93 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_93 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_93 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_93 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_93 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_93 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_94 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h5E;
  wire          compressDataVec_hitReq_1_94 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h5E;
  wire          compressDataVec_hitReq_2_94 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h5E;
  wire          compressDataVec_hitReq_3_94 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h5E;
  wire          compressDataVec_hitReq_4_94 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h5E;
  wire          compressDataVec_hitReq_5_94 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h5E;
  wire          compressDataVec_hitReq_6_94 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h5E;
  wire          compressDataVec_hitReq_7_94 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h5E;
  wire          compressDataVec_hitReq_8_94 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h5E;
  wire          compressDataVec_hitReq_9_94 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h5E;
  wire          compressDataVec_hitReq_10_94 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h5E;
  wire          compressDataVec_hitReq_11_94 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h5E;
  wire          compressDataVec_hitReq_12_94 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h5E;
  wire          compressDataVec_hitReq_13_94 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h5E;
  wire          compressDataVec_hitReq_14_94 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h5E;
  wire          compressDataVec_hitReq_15_94 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h5E;
  wire          compressDataVec_hitReq_16_94 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h5E;
  wire          compressDataVec_hitReq_17_94 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h5E;
  wire          compressDataVec_hitReq_18_94 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h5E;
  wire          compressDataVec_hitReq_19_94 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h5E;
  wire          compressDataVec_hitReq_20_94 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h5E;
  wire          compressDataVec_hitReq_21_94 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h5E;
  wire          compressDataVec_hitReq_22_94 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h5E;
  wire          compressDataVec_hitReq_23_94 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h5E;
  wire          compressDataVec_hitReq_24_94 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h5E;
  wire          compressDataVec_hitReq_25_94 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h5E;
  wire          compressDataVec_hitReq_26_94 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h5E;
  wire          compressDataVec_hitReq_27_94 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h5E;
  wire          compressDataVec_hitReq_28_94 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h5E;
  wire          compressDataVec_hitReq_29_94 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h5E;
  wire          compressDataVec_hitReq_30_94 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h5E;
  wire          compressDataVec_hitReq_31_94 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h5E;
  wire          compressDataVec_hitReq_32_94 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h5E;
  wire          compressDataVec_hitReq_33_94 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h5E;
  wire          compressDataVec_hitReq_34_94 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h5E;
  wire          compressDataVec_hitReq_35_94 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h5E;
  wire          compressDataVec_hitReq_36_94 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h5E;
  wire          compressDataVec_hitReq_37_94 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h5E;
  wire          compressDataVec_hitReq_38_94 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h5E;
  wire          compressDataVec_hitReq_39_94 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h5E;
  wire          compressDataVec_hitReq_40_94 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h5E;
  wire          compressDataVec_hitReq_41_94 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h5E;
  wire          compressDataVec_hitReq_42_94 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h5E;
  wire          compressDataVec_hitReq_43_94 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h5E;
  wire          compressDataVec_hitReq_44_94 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h5E;
  wire          compressDataVec_hitReq_45_94 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h5E;
  wire          compressDataVec_hitReq_46_94 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h5E;
  wire          compressDataVec_hitReq_47_94 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h5E;
  wire          compressDataVec_hitReq_48_94 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h5E;
  wire          compressDataVec_hitReq_49_94 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h5E;
  wire          compressDataVec_hitReq_50_94 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h5E;
  wire          compressDataVec_hitReq_51_94 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h5E;
  wire          compressDataVec_hitReq_52_94 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h5E;
  wire          compressDataVec_hitReq_53_94 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h5E;
  wire          compressDataVec_hitReq_54_94 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h5E;
  wire          compressDataVec_hitReq_55_94 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h5E;
  wire          compressDataVec_hitReq_56_94 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h5E;
  wire          compressDataVec_hitReq_57_94 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h5E;
  wire          compressDataVec_hitReq_58_94 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h5E;
  wire          compressDataVec_hitReq_59_94 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h5E;
  wire          compressDataVec_hitReq_60_94 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h5E;
  wire          compressDataVec_hitReq_61_94 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h5E;
  wire          compressDataVec_hitReq_62_94 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h5E;
  wire          compressDataVec_hitReq_63_94 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h5E;
  wire [7:0]    compressDataVec_selectReqData_94 =
    (compressDataVec_hitReq_0_94 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_94 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_94 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_94 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_94 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_94 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_94 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_94 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_94 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_94 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_94 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_94 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_94 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_94 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_94 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_94 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_94 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_94 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_94 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_94 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_94 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_94 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_94 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_94 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_94 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_94 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_94 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_94 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_94 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_94 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_94 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_94 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_94 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_94 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_94 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_94 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_94 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_94 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_94 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_94 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_94 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_94 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_94 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_94 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_94 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_94 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_94 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_94 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_94 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_94 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_94 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_94 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_94 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_94 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_94 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_94 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_94 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_94 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_94 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_94 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_94 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_94 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_94 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_94 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_95 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h5F;
  wire          compressDataVec_hitReq_1_95 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h5F;
  wire          compressDataVec_hitReq_2_95 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h5F;
  wire          compressDataVec_hitReq_3_95 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h5F;
  wire          compressDataVec_hitReq_4_95 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h5F;
  wire          compressDataVec_hitReq_5_95 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h5F;
  wire          compressDataVec_hitReq_6_95 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h5F;
  wire          compressDataVec_hitReq_7_95 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h5F;
  wire          compressDataVec_hitReq_8_95 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h5F;
  wire          compressDataVec_hitReq_9_95 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h5F;
  wire          compressDataVec_hitReq_10_95 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h5F;
  wire          compressDataVec_hitReq_11_95 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h5F;
  wire          compressDataVec_hitReq_12_95 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h5F;
  wire          compressDataVec_hitReq_13_95 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h5F;
  wire          compressDataVec_hitReq_14_95 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h5F;
  wire          compressDataVec_hitReq_15_95 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h5F;
  wire          compressDataVec_hitReq_16_95 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h5F;
  wire          compressDataVec_hitReq_17_95 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h5F;
  wire          compressDataVec_hitReq_18_95 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h5F;
  wire          compressDataVec_hitReq_19_95 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h5F;
  wire          compressDataVec_hitReq_20_95 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h5F;
  wire          compressDataVec_hitReq_21_95 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h5F;
  wire          compressDataVec_hitReq_22_95 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h5F;
  wire          compressDataVec_hitReq_23_95 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h5F;
  wire          compressDataVec_hitReq_24_95 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h5F;
  wire          compressDataVec_hitReq_25_95 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h5F;
  wire          compressDataVec_hitReq_26_95 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h5F;
  wire          compressDataVec_hitReq_27_95 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h5F;
  wire          compressDataVec_hitReq_28_95 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h5F;
  wire          compressDataVec_hitReq_29_95 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h5F;
  wire          compressDataVec_hitReq_30_95 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h5F;
  wire          compressDataVec_hitReq_31_95 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h5F;
  wire          compressDataVec_hitReq_32_95 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h5F;
  wire          compressDataVec_hitReq_33_95 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h5F;
  wire          compressDataVec_hitReq_34_95 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h5F;
  wire          compressDataVec_hitReq_35_95 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h5F;
  wire          compressDataVec_hitReq_36_95 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h5F;
  wire          compressDataVec_hitReq_37_95 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h5F;
  wire          compressDataVec_hitReq_38_95 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h5F;
  wire          compressDataVec_hitReq_39_95 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h5F;
  wire          compressDataVec_hitReq_40_95 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h5F;
  wire          compressDataVec_hitReq_41_95 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h5F;
  wire          compressDataVec_hitReq_42_95 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h5F;
  wire          compressDataVec_hitReq_43_95 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h5F;
  wire          compressDataVec_hitReq_44_95 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h5F;
  wire          compressDataVec_hitReq_45_95 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h5F;
  wire          compressDataVec_hitReq_46_95 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h5F;
  wire          compressDataVec_hitReq_47_95 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h5F;
  wire          compressDataVec_hitReq_48_95 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h5F;
  wire          compressDataVec_hitReq_49_95 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h5F;
  wire          compressDataVec_hitReq_50_95 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h5F;
  wire          compressDataVec_hitReq_51_95 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h5F;
  wire          compressDataVec_hitReq_52_95 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h5F;
  wire          compressDataVec_hitReq_53_95 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h5F;
  wire          compressDataVec_hitReq_54_95 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h5F;
  wire          compressDataVec_hitReq_55_95 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h5F;
  wire          compressDataVec_hitReq_56_95 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h5F;
  wire          compressDataVec_hitReq_57_95 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h5F;
  wire          compressDataVec_hitReq_58_95 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h5F;
  wire          compressDataVec_hitReq_59_95 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h5F;
  wire          compressDataVec_hitReq_60_95 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h5F;
  wire          compressDataVec_hitReq_61_95 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h5F;
  wire          compressDataVec_hitReq_62_95 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h5F;
  wire          compressDataVec_hitReq_63_95 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h5F;
  wire [7:0]    compressDataVec_selectReqData_95 =
    (compressDataVec_hitReq_0_95 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_95 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_95 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_95 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_95 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_95 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_95 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_95 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_95 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_95 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_95 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_95 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_95 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_95 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_95 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_95 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_95 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_95 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_95 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_95 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_95 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_95 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_95 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_95 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_95 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_95 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_95 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_95 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_95 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_95 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_95 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_95 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_95 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_95 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_95 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_95 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_95 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_95 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_95 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_95 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_95 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_95 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_95 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_95 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_95 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_95 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_95 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_95 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_95 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_95 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_95 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_95 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_95 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_95 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_95 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_95 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_95 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_95 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_95 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_95 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_95 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_95 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_95 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_95 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_96 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h60;
  wire          compressDataVec_hitReq_1_96 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h60;
  wire          compressDataVec_hitReq_2_96 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h60;
  wire          compressDataVec_hitReq_3_96 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h60;
  wire          compressDataVec_hitReq_4_96 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h60;
  wire          compressDataVec_hitReq_5_96 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h60;
  wire          compressDataVec_hitReq_6_96 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h60;
  wire          compressDataVec_hitReq_7_96 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h60;
  wire          compressDataVec_hitReq_8_96 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h60;
  wire          compressDataVec_hitReq_9_96 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h60;
  wire          compressDataVec_hitReq_10_96 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h60;
  wire          compressDataVec_hitReq_11_96 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h60;
  wire          compressDataVec_hitReq_12_96 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h60;
  wire          compressDataVec_hitReq_13_96 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h60;
  wire          compressDataVec_hitReq_14_96 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h60;
  wire          compressDataVec_hitReq_15_96 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h60;
  wire          compressDataVec_hitReq_16_96 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h60;
  wire          compressDataVec_hitReq_17_96 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h60;
  wire          compressDataVec_hitReq_18_96 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h60;
  wire          compressDataVec_hitReq_19_96 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h60;
  wire          compressDataVec_hitReq_20_96 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h60;
  wire          compressDataVec_hitReq_21_96 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h60;
  wire          compressDataVec_hitReq_22_96 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h60;
  wire          compressDataVec_hitReq_23_96 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h60;
  wire          compressDataVec_hitReq_24_96 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h60;
  wire          compressDataVec_hitReq_25_96 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h60;
  wire          compressDataVec_hitReq_26_96 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h60;
  wire          compressDataVec_hitReq_27_96 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h60;
  wire          compressDataVec_hitReq_28_96 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h60;
  wire          compressDataVec_hitReq_29_96 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h60;
  wire          compressDataVec_hitReq_30_96 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h60;
  wire          compressDataVec_hitReq_31_96 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h60;
  wire          compressDataVec_hitReq_32_96 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h60;
  wire          compressDataVec_hitReq_33_96 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h60;
  wire          compressDataVec_hitReq_34_96 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h60;
  wire          compressDataVec_hitReq_35_96 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h60;
  wire          compressDataVec_hitReq_36_96 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h60;
  wire          compressDataVec_hitReq_37_96 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h60;
  wire          compressDataVec_hitReq_38_96 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h60;
  wire          compressDataVec_hitReq_39_96 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h60;
  wire          compressDataVec_hitReq_40_96 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h60;
  wire          compressDataVec_hitReq_41_96 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h60;
  wire          compressDataVec_hitReq_42_96 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h60;
  wire          compressDataVec_hitReq_43_96 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h60;
  wire          compressDataVec_hitReq_44_96 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h60;
  wire          compressDataVec_hitReq_45_96 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h60;
  wire          compressDataVec_hitReq_46_96 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h60;
  wire          compressDataVec_hitReq_47_96 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h60;
  wire          compressDataVec_hitReq_48_96 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h60;
  wire          compressDataVec_hitReq_49_96 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h60;
  wire          compressDataVec_hitReq_50_96 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h60;
  wire          compressDataVec_hitReq_51_96 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h60;
  wire          compressDataVec_hitReq_52_96 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h60;
  wire          compressDataVec_hitReq_53_96 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h60;
  wire          compressDataVec_hitReq_54_96 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h60;
  wire          compressDataVec_hitReq_55_96 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h60;
  wire          compressDataVec_hitReq_56_96 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h60;
  wire          compressDataVec_hitReq_57_96 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h60;
  wire          compressDataVec_hitReq_58_96 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h60;
  wire          compressDataVec_hitReq_59_96 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h60;
  wire          compressDataVec_hitReq_60_96 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h60;
  wire          compressDataVec_hitReq_61_96 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h60;
  wire          compressDataVec_hitReq_62_96 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h60;
  wire          compressDataVec_hitReq_63_96 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h60;
  wire [7:0]    compressDataVec_selectReqData_96 =
    (compressDataVec_hitReq_0_96 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_96 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_96 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_96 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_96 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_96 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_96 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_96 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_96 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_96 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_96 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_96 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_96 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_96 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_96 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_96 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_96 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_96 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_96 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_96 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_96 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_96 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_96 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_96 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_96 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_96 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_96 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_96 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_96 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_96 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_96 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_96 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_96 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_96 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_96 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_96 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_96 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_96 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_96 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_96 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_96 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_96 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_96 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_96 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_96 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_96 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_96 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_96 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_96 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_96 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_96 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_96 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_96 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_96 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_96 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_96 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_96 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_96 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_96 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_96 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_96 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_96 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_96 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_96 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_97 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h61;
  wire          compressDataVec_hitReq_1_97 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h61;
  wire          compressDataVec_hitReq_2_97 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h61;
  wire          compressDataVec_hitReq_3_97 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h61;
  wire          compressDataVec_hitReq_4_97 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h61;
  wire          compressDataVec_hitReq_5_97 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h61;
  wire          compressDataVec_hitReq_6_97 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h61;
  wire          compressDataVec_hitReq_7_97 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h61;
  wire          compressDataVec_hitReq_8_97 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h61;
  wire          compressDataVec_hitReq_9_97 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h61;
  wire          compressDataVec_hitReq_10_97 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h61;
  wire          compressDataVec_hitReq_11_97 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h61;
  wire          compressDataVec_hitReq_12_97 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h61;
  wire          compressDataVec_hitReq_13_97 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h61;
  wire          compressDataVec_hitReq_14_97 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h61;
  wire          compressDataVec_hitReq_15_97 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h61;
  wire          compressDataVec_hitReq_16_97 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h61;
  wire          compressDataVec_hitReq_17_97 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h61;
  wire          compressDataVec_hitReq_18_97 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h61;
  wire          compressDataVec_hitReq_19_97 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h61;
  wire          compressDataVec_hitReq_20_97 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h61;
  wire          compressDataVec_hitReq_21_97 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h61;
  wire          compressDataVec_hitReq_22_97 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h61;
  wire          compressDataVec_hitReq_23_97 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h61;
  wire          compressDataVec_hitReq_24_97 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h61;
  wire          compressDataVec_hitReq_25_97 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h61;
  wire          compressDataVec_hitReq_26_97 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h61;
  wire          compressDataVec_hitReq_27_97 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h61;
  wire          compressDataVec_hitReq_28_97 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h61;
  wire          compressDataVec_hitReq_29_97 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h61;
  wire          compressDataVec_hitReq_30_97 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h61;
  wire          compressDataVec_hitReq_31_97 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h61;
  wire          compressDataVec_hitReq_32_97 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h61;
  wire          compressDataVec_hitReq_33_97 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h61;
  wire          compressDataVec_hitReq_34_97 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h61;
  wire          compressDataVec_hitReq_35_97 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h61;
  wire          compressDataVec_hitReq_36_97 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h61;
  wire          compressDataVec_hitReq_37_97 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h61;
  wire          compressDataVec_hitReq_38_97 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h61;
  wire          compressDataVec_hitReq_39_97 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h61;
  wire          compressDataVec_hitReq_40_97 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h61;
  wire          compressDataVec_hitReq_41_97 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h61;
  wire          compressDataVec_hitReq_42_97 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h61;
  wire          compressDataVec_hitReq_43_97 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h61;
  wire          compressDataVec_hitReq_44_97 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h61;
  wire          compressDataVec_hitReq_45_97 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h61;
  wire          compressDataVec_hitReq_46_97 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h61;
  wire          compressDataVec_hitReq_47_97 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h61;
  wire          compressDataVec_hitReq_48_97 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h61;
  wire          compressDataVec_hitReq_49_97 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h61;
  wire          compressDataVec_hitReq_50_97 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h61;
  wire          compressDataVec_hitReq_51_97 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h61;
  wire          compressDataVec_hitReq_52_97 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h61;
  wire          compressDataVec_hitReq_53_97 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h61;
  wire          compressDataVec_hitReq_54_97 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h61;
  wire          compressDataVec_hitReq_55_97 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h61;
  wire          compressDataVec_hitReq_56_97 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h61;
  wire          compressDataVec_hitReq_57_97 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h61;
  wire          compressDataVec_hitReq_58_97 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h61;
  wire          compressDataVec_hitReq_59_97 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h61;
  wire          compressDataVec_hitReq_60_97 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h61;
  wire          compressDataVec_hitReq_61_97 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h61;
  wire          compressDataVec_hitReq_62_97 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h61;
  wire          compressDataVec_hitReq_63_97 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h61;
  wire [7:0]    compressDataVec_selectReqData_97 =
    (compressDataVec_hitReq_0_97 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_97 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_97 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_97 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_97 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_97 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_97 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_97 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_97 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_97 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_97 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_97 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_97 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_97 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_97 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_97 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_97 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_97 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_97 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_97 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_97 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_97 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_97 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_97 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_97 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_97 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_97 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_97 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_97 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_97 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_97 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_97 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_97 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_97 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_97 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_97 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_97 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_97 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_97 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_97 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_97 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_97 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_97 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_97 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_97 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_97 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_97 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_97 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_97 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_97 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_97 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_97 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_97 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_97 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_97 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_97 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_97 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_97 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_97 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_97 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_97 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_97 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_97 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_97 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_98 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h62;
  wire          compressDataVec_hitReq_1_98 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h62;
  wire          compressDataVec_hitReq_2_98 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h62;
  wire          compressDataVec_hitReq_3_98 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h62;
  wire          compressDataVec_hitReq_4_98 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h62;
  wire          compressDataVec_hitReq_5_98 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h62;
  wire          compressDataVec_hitReq_6_98 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h62;
  wire          compressDataVec_hitReq_7_98 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h62;
  wire          compressDataVec_hitReq_8_98 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h62;
  wire          compressDataVec_hitReq_9_98 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h62;
  wire          compressDataVec_hitReq_10_98 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h62;
  wire          compressDataVec_hitReq_11_98 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h62;
  wire          compressDataVec_hitReq_12_98 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h62;
  wire          compressDataVec_hitReq_13_98 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h62;
  wire          compressDataVec_hitReq_14_98 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h62;
  wire          compressDataVec_hitReq_15_98 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h62;
  wire          compressDataVec_hitReq_16_98 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h62;
  wire          compressDataVec_hitReq_17_98 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h62;
  wire          compressDataVec_hitReq_18_98 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h62;
  wire          compressDataVec_hitReq_19_98 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h62;
  wire          compressDataVec_hitReq_20_98 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h62;
  wire          compressDataVec_hitReq_21_98 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h62;
  wire          compressDataVec_hitReq_22_98 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h62;
  wire          compressDataVec_hitReq_23_98 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h62;
  wire          compressDataVec_hitReq_24_98 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h62;
  wire          compressDataVec_hitReq_25_98 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h62;
  wire          compressDataVec_hitReq_26_98 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h62;
  wire          compressDataVec_hitReq_27_98 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h62;
  wire          compressDataVec_hitReq_28_98 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h62;
  wire          compressDataVec_hitReq_29_98 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h62;
  wire          compressDataVec_hitReq_30_98 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h62;
  wire          compressDataVec_hitReq_31_98 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h62;
  wire          compressDataVec_hitReq_32_98 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h62;
  wire          compressDataVec_hitReq_33_98 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h62;
  wire          compressDataVec_hitReq_34_98 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h62;
  wire          compressDataVec_hitReq_35_98 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h62;
  wire          compressDataVec_hitReq_36_98 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h62;
  wire          compressDataVec_hitReq_37_98 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h62;
  wire          compressDataVec_hitReq_38_98 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h62;
  wire          compressDataVec_hitReq_39_98 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h62;
  wire          compressDataVec_hitReq_40_98 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h62;
  wire          compressDataVec_hitReq_41_98 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h62;
  wire          compressDataVec_hitReq_42_98 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h62;
  wire          compressDataVec_hitReq_43_98 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h62;
  wire          compressDataVec_hitReq_44_98 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h62;
  wire          compressDataVec_hitReq_45_98 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h62;
  wire          compressDataVec_hitReq_46_98 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h62;
  wire          compressDataVec_hitReq_47_98 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h62;
  wire          compressDataVec_hitReq_48_98 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h62;
  wire          compressDataVec_hitReq_49_98 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h62;
  wire          compressDataVec_hitReq_50_98 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h62;
  wire          compressDataVec_hitReq_51_98 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h62;
  wire          compressDataVec_hitReq_52_98 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h62;
  wire          compressDataVec_hitReq_53_98 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h62;
  wire          compressDataVec_hitReq_54_98 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h62;
  wire          compressDataVec_hitReq_55_98 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h62;
  wire          compressDataVec_hitReq_56_98 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h62;
  wire          compressDataVec_hitReq_57_98 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h62;
  wire          compressDataVec_hitReq_58_98 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h62;
  wire          compressDataVec_hitReq_59_98 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h62;
  wire          compressDataVec_hitReq_60_98 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h62;
  wire          compressDataVec_hitReq_61_98 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h62;
  wire          compressDataVec_hitReq_62_98 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h62;
  wire          compressDataVec_hitReq_63_98 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h62;
  wire [7:0]    compressDataVec_selectReqData_98 =
    (compressDataVec_hitReq_0_98 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_98 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_98 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_98 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_98 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_98 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_98 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_98 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_98 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_98 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_98 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_98 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_98 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_98 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_98 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_98 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_98 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_98 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_98 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_98 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_98 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_98 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_98 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_98 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_98 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_98 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_98 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_98 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_98 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_98 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_98 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_98 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_98 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_98 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_98 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_98 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_98 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_98 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_98 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_98 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_98 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_98 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_98 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_98 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_98 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_98 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_98 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_98 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_98 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_98 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_98 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_98 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_98 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_98 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_98 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_98 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_98 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_98 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_98 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_98 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_98 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_98 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_98 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_98 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_99 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h63;
  wire          compressDataVec_hitReq_1_99 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h63;
  wire          compressDataVec_hitReq_2_99 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h63;
  wire          compressDataVec_hitReq_3_99 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h63;
  wire          compressDataVec_hitReq_4_99 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h63;
  wire          compressDataVec_hitReq_5_99 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h63;
  wire          compressDataVec_hitReq_6_99 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h63;
  wire          compressDataVec_hitReq_7_99 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h63;
  wire          compressDataVec_hitReq_8_99 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h63;
  wire          compressDataVec_hitReq_9_99 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h63;
  wire          compressDataVec_hitReq_10_99 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h63;
  wire          compressDataVec_hitReq_11_99 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h63;
  wire          compressDataVec_hitReq_12_99 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h63;
  wire          compressDataVec_hitReq_13_99 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h63;
  wire          compressDataVec_hitReq_14_99 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h63;
  wire          compressDataVec_hitReq_15_99 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h63;
  wire          compressDataVec_hitReq_16_99 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h63;
  wire          compressDataVec_hitReq_17_99 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h63;
  wire          compressDataVec_hitReq_18_99 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h63;
  wire          compressDataVec_hitReq_19_99 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h63;
  wire          compressDataVec_hitReq_20_99 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h63;
  wire          compressDataVec_hitReq_21_99 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h63;
  wire          compressDataVec_hitReq_22_99 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h63;
  wire          compressDataVec_hitReq_23_99 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h63;
  wire          compressDataVec_hitReq_24_99 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h63;
  wire          compressDataVec_hitReq_25_99 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h63;
  wire          compressDataVec_hitReq_26_99 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h63;
  wire          compressDataVec_hitReq_27_99 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h63;
  wire          compressDataVec_hitReq_28_99 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h63;
  wire          compressDataVec_hitReq_29_99 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h63;
  wire          compressDataVec_hitReq_30_99 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h63;
  wire          compressDataVec_hitReq_31_99 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h63;
  wire          compressDataVec_hitReq_32_99 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h63;
  wire          compressDataVec_hitReq_33_99 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h63;
  wire          compressDataVec_hitReq_34_99 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h63;
  wire          compressDataVec_hitReq_35_99 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h63;
  wire          compressDataVec_hitReq_36_99 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h63;
  wire          compressDataVec_hitReq_37_99 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h63;
  wire          compressDataVec_hitReq_38_99 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h63;
  wire          compressDataVec_hitReq_39_99 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h63;
  wire          compressDataVec_hitReq_40_99 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h63;
  wire          compressDataVec_hitReq_41_99 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h63;
  wire          compressDataVec_hitReq_42_99 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h63;
  wire          compressDataVec_hitReq_43_99 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h63;
  wire          compressDataVec_hitReq_44_99 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h63;
  wire          compressDataVec_hitReq_45_99 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h63;
  wire          compressDataVec_hitReq_46_99 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h63;
  wire          compressDataVec_hitReq_47_99 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h63;
  wire          compressDataVec_hitReq_48_99 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h63;
  wire          compressDataVec_hitReq_49_99 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h63;
  wire          compressDataVec_hitReq_50_99 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h63;
  wire          compressDataVec_hitReq_51_99 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h63;
  wire          compressDataVec_hitReq_52_99 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h63;
  wire          compressDataVec_hitReq_53_99 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h63;
  wire          compressDataVec_hitReq_54_99 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h63;
  wire          compressDataVec_hitReq_55_99 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h63;
  wire          compressDataVec_hitReq_56_99 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h63;
  wire          compressDataVec_hitReq_57_99 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h63;
  wire          compressDataVec_hitReq_58_99 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h63;
  wire          compressDataVec_hitReq_59_99 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h63;
  wire          compressDataVec_hitReq_60_99 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h63;
  wire          compressDataVec_hitReq_61_99 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h63;
  wire          compressDataVec_hitReq_62_99 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h63;
  wire          compressDataVec_hitReq_63_99 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h63;
  wire [7:0]    compressDataVec_selectReqData_99 =
    (compressDataVec_hitReq_0_99 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_99 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_99 ? source2Pipe[23:16] : 8'h0) | (compressDataVec_hitReq_3_99 ? source2Pipe[31:24] : 8'h0)
    | (compressDataVec_hitReq_4_99 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_99 ? source2Pipe[47:40] : 8'h0) | (compressDataVec_hitReq_6_99 ? source2Pipe[55:48] : 8'h0)
    | (compressDataVec_hitReq_7_99 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_99 ? source2Pipe[71:64] : 8'h0) | (compressDataVec_hitReq_9_99 ? source2Pipe[79:72] : 8'h0)
    | (compressDataVec_hitReq_10_99 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_99 ? source2Pipe[95:88] : 8'h0) | (compressDataVec_hitReq_12_99 ? source2Pipe[103:96] : 8'h0)
    | (compressDataVec_hitReq_13_99 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_99 ? source2Pipe[119:112] : 8'h0) | (compressDataVec_hitReq_15_99 ? source2Pipe[127:120] : 8'h0)
    | (compressDataVec_hitReq_16_99 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_99 ? source2Pipe[143:136] : 8'h0) | (compressDataVec_hitReq_18_99 ? source2Pipe[151:144] : 8'h0)
    | (compressDataVec_hitReq_19_99 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_99 ? source2Pipe[167:160] : 8'h0) | (compressDataVec_hitReq_21_99 ? source2Pipe[175:168] : 8'h0)
    | (compressDataVec_hitReq_22_99 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_99 ? source2Pipe[191:184] : 8'h0) | (compressDataVec_hitReq_24_99 ? source2Pipe[199:192] : 8'h0)
    | (compressDataVec_hitReq_25_99 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_99 ? source2Pipe[215:208] : 8'h0) | (compressDataVec_hitReq_27_99 ? source2Pipe[223:216] : 8'h0)
    | (compressDataVec_hitReq_28_99 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_99 ? source2Pipe[239:232] : 8'h0) | (compressDataVec_hitReq_30_99 ? source2Pipe[247:240] : 8'h0)
    | (compressDataVec_hitReq_31_99 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_99 ? source2Pipe[263:256] : 8'h0) | (compressDataVec_hitReq_33_99 ? source2Pipe[271:264] : 8'h0)
    | (compressDataVec_hitReq_34_99 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_99 ? source2Pipe[287:280] : 8'h0) | (compressDataVec_hitReq_36_99 ? source2Pipe[295:288] : 8'h0)
    | (compressDataVec_hitReq_37_99 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_99 ? source2Pipe[311:304] : 8'h0) | (compressDataVec_hitReq_39_99 ? source2Pipe[319:312] : 8'h0)
    | (compressDataVec_hitReq_40_99 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_99 ? source2Pipe[335:328] : 8'h0) | (compressDataVec_hitReq_42_99 ? source2Pipe[343:336] : 8'h0)
    | (compressDataVec_hitReq_43_99 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_99 ? source2Pipe[359:352] : 8'h0) | (compressDataVec_hitReq_45_99 ? source2Pipe[367:360] : 8'h0)
    | (compressDataVec_hitReq_46_99 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_99 ? source2Pipe[383:376] : 8'h0) | (compressDataVec_hitReq_48_99 ? source2Pipe[391:384] : 8'h0)
    | (compressDataVec_hitReq_49_99 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_99 ? source2Pipe[407:400] : 8'h0) | (compressDataVec_hitReq_51_99 ? source2Pipe[415:408] : 8'h0)
    | (compressDataVec_hitReq_52_99 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_99 ? source2Pipe[431:424] : 8'h0) | (compressDataVec_hitReq_54_99 ? source2Pipe[439:432] : 8'h0)
    | (compressDataVec_hitReq_55_99 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_99 ? source2Pipe[455:448] : 8'h0) | (compressDataVec_hitReq_57_99 ? source2Pipe[463:456] : 8'h0)
    | (compressDataVec_hitReq_58_99 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_99 ? source2Pipe[479:472] : 8'h0) | (compressDataVec_hitReq_60_99 ? source2Pipe[487:480] : 8'h0)
    | (compressDataVec_hitReq_61_99 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_99 ? source2Pipe[503:496] : 8'h0) | (compressDataVec_hitReq_63_99 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_100 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h64;
  wire          compressDataVec_hitReq_1_100 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h64;
  wire          compressDataVec_hitReq_2_100 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h64;
  wire          compressDataVec_hitReq_3_100 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h64;
  wire          compressDataVec_hitReq_4_100 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h64;
  wire          compressDataVec_hitReq_5_100 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h64;
  wire          compressDataVec_hitReq_6_100 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h64;
  wire          compressDataVec_hitReq_7_100 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h64;
  wire          compressDataVec_hitReq_8_100 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h64;
  wire          compressDataVec_hitReq_9_100 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h64;
  wire          compressDataVec_hitReq_10_100 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h64;
  wire          compressDataVec_hitReq_11_100 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h64;
  wire          compressDataVec_hitReq_12_100 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h64;
  wire          compressDataVec_hitReq_13_100 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h64;
  wire          compressDataVec_hitReq_14_100 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h64;
  wire          compressDataVec_hitReq_15_100 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h64;
  wire          compressDataVec_hitReq_16_100 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h64;
  wire          compressDataVec_hitReq_17_100 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h64;
  wire          compressDataVec_hitReq_18_100 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h64;
  wire          compressDataVec_hitReq_19_100 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h64;
  wire          compressDataVec_hitReq_20_100 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h64;
  wire          compressDataVec_hitReq_21_100 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h64;
  wire          compressDataVec_hitReq_22_100 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h64;
  wire          compressDataVec_hitReq_23_100 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h64;
  wire          compressDataVec_hitReq_24_100 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h64;
  wire          compressDataVec_hitReq_25_100 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h64;
  wire          compressDataVec_hitReq_26_100 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h64;
  wire          compressDataVec_hitReq_27_100 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h64;
  wire          compressDataVec_hitReq_28_100 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h64;
  wire          compressDataVec_hitReq_29_100 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h64;
  wire          compressDataVec_hitReq_30_100 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h64;
  wire          compressDataVec_hitReq_31_100 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h64;
  wire          compressDataVec_hitReq_32_100 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h64;
  wire          compressDataVec_hitReq_33_100 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h64;
  wire          compressDataVec_hitReq_34_100 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h64;
  wire          compressDataVec_hitReq_35_100 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h64;
  wire          compressDataVec_hitReq_36_100 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h64;
  wire          compressDataVec_hitReq_37_100 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h64;
  wire          compressDataVec_hitReq_38_100 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h64;
  wire          compressDataVec_hitReq_39_100 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h64;
  wire          compressDataVec_hitReq_40_100 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h64;
  wire          compressDataVec_hitReq_41_100 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h64;
  wire          compressDataVec_hitReq_42_100 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h64;
  wire          compressDataVec_hitReq_43_100 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h64;
  wire          compressDataVec_hitReq_44_100 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h64;
  wire          compressDataVec_hitReq_45_100 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h64;
  wire          compressDataVec_hitReq_46_100 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h64;
  wire          compressDataVec_hitReq_47_100 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h64;
  wire          compressDataVec_hitReq_48_100 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h64;
  wire          compressDataVec_hitReq_49_100 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h64;
  wire          compressDataVec_hitReq_50_100 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h64;
  wire          compressDataVec_hitReq_51_100 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h64;
  wire          compressDataVec_hitReq_52_100 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h64;
  wire          compressDataVec_hitReq_53_100 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h64;
  wire          compressDataVec_hitReq_54_100 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h64;
  wire          compressDataVec_hitReq_55_100 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h64;
  wire          compressDataVec_hitReq_56_100 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h64;
  wire          compressDataVec_hitReq_57_100 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h64;
  wire          compressDataVec_hitReq_58_100 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h64;
  wire          compressDataVec_hitReq_59_100 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h64;
  wire          compressDataVec_hitReq_60_100 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h64;
  wire          compressDataVec_hitReq_61_100 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h64;
  wire          compressDataVec_hitReq_62_100 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h64;
  wire          compressDataVec_hitReq_63_100 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h64;
  wire [7:0]    compressDataVec_selectReqData_100 =
    (compressDataVec_hitReq_0_100 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_100 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_100 ? source2Pipe[23:16] : 8'h0)
    | (compressDataVec_hitReq_3_100 ? source2Pipe[31:24] : 8'h0) | (compressDataVec_hitReq_4_100 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_100 ? source2Pipe[47:40] : 8'h0)
    | (compressDataVec_hitReq_6_100 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_100 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_100 ? source2Pipe[71:64] : 8'h0)
    | (compressDataVec_hitReq_9_100 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_100 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_100 ? source2Pipe[95:88] : 8'h0)
    | (compressDataVec_hitReq_12_100 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_100 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_100 ? source2Pipe[119:112] : 8'h0)
    | (compressDataVec_hitReq_15_100 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_100 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_100 ? source2Pipe[143:136] : 8'h0)
    | (compressDataVec_hitReq_18_100 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_100 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_100 ? source2Pipe[167:160] : 8'h0)
    | (compressDataVec_hitReq_21_100 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_100 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_100 ? source2Pipe[191:184] : 8'h0)
    | (compressDataVec_hitReq_24_100 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_100 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_100 ? source2Pipe[215:208] : 8'h0)
    | (compressDataVec_hitReq_27_100 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_100 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_100 ? source2Pipe[239:232] : 8'h0)
    | (compressDataVec_hitReq_30_100 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_100 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_100 ? source2Pipe[263:256] : 8'h0)
    | (compressDataVec_hitReq_33_100 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_100 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_100 ? source2Pipe[287:280] : 8'h0)
    | (compressDataVec_hitReq_36_100 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_100 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_100 ? source2Pipe[311:304] : 8'h0)
    | (compressDataVec_hitReq_39_100 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_100 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_100 ? source2Pipe[335:328] : 8'h0)
    | (compressDataVec_hitReq_42_100 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_100 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_100 ? source2Pipe[359:352] : 8'h0)
    | (compressDataVec_hitReq_45_100 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_100 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_100 ? source2Pipe[383:376] : 8'h0)
    | (compressDataVec_hitReq_48_100 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_100 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_100 ? source2Pipe[407:400] : 8'h0)
    | (compressDataVec_hitReq_51_100 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_100 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_100 ? source2Pipe[431:424] : 8'h0)
    | (compressDataVec_hitReq_54_100 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_100 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_100 ? source2Pipe[455:448] : 8'h0)
    | (compressDataVec_hitReq_57_100 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_100 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_100 ? source2Pipe[479:472] : 8'h0)
    | (compressDataVec_hitReq_60_100 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_100 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_100 ? source2Pipe[503:496] : 8'h0)
    | (compressDataVec_hitReq_63_100 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_101 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h65;
  wire          compressDataVec_hitReq_1_101 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h65;
  wire          compressDataVec_hitReq_2_101 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h65;
  wire          compressDataVec_hitReq_3_101 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h65;
  wire          compressDataVec_hitReq_4_101 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h65;
  wire          compressDataVec_hitReq_5_101 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h65;
  wire          compressDataVec_hitReq_6_101 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h65;
  wire          compressDataVec_hitReq_7_101 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h65;
  wire          compressDataVec_hitReq_8_101 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h65;
  wire          compressDataVec_hitReq_9_101 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h65;
  wire          compressDataVec_hitReq_10_101 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h65;
  wire          compressDataVec_hitReq_11_101 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h65;
  wire          compressDataVec_hitReq_12_101 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h65;
  wire          compressDataVec_hitReq_13_101 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h65;
  wire          compressDataVec_hitReq_14_101 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h65;
  wire          compressDataVec_hitReq_15_101 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h65;
  wire          compressDataVec_hitReq_16_101 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h65;
  wire          compressDataVec_hitReq_17_101 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h65;
  wire          compressDataVec_hitReq_18_101 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h65;
  wire          compressDataVec_hitReq_19_101 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h65;
  wire          compressDataVec_hitReq_20_101 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h65;
  wire          compressDataVec_hitReq_21_101 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h65;
  wire          compressDataVec_hitReq_22_101 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h65;
  wire          compressDataVec_hitReq_23_101 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h65;
  wire          compressDataVec_hitReq_24_101 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h65;
  wire          compressDataVec_hitReq_25_101 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h65;
  wire          compressDataVec_hitReq_26_101 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h65;
  wire          compressDataVec_hitReq_27_101 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h65;
  wire          compressDataVec_hitReq_28_101 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h65;
  wire          compressDataVec_hitReq_29_101 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h65;
  wire          compressDataVec_hitReq_30_101 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h65;
  wire          compressDataVec_hitReq_31_101 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h65;
  wire          compressDataVec_hitReq_32_101 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h65;
  wire          compressDataVec_hitReq_33_101 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h65;
  wire          compressDataVec_hitReq_34_101 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h65;
  wire          compressDataVec_hitReq_35_101 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h65;
  wire          compressDataVec_hitReq_36_101 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h65;
  wire          compressDataVec_hitReq_37_101 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h65;
  wire          compressDataVec_hitReq_38_101 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h65;
  wire          compressDataVec_hitReq_39_101 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h65;
  wire          compressDataVec_hitReq_40_101 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h65;
  wire          compressDataVec_hitReq_41_101 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h65;
  wire          compressDataVec_hitReq_42_101 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h65;
  wire          compressDataVec_hitReq_43_101 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h65;
  wire          compressDataVec_hitReq_44_101 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h65;
  wire          compressDataVec_hitReq_45_101 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h65;
  wire          compressDataVec_hitReq_46_101 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h65;
  wire          compressDataVec_hitReq_47_101 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h65;
  wire          compressDataVec_hitReq_48_101 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h65;
  wire          compressDataVec_hitReq_49_101 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h65;
  wire          compressDataVec_hitReq_50_101 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h65;
  wire          compressDataVec_hitReq_51_101 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h65;
  wire          compressDataVec_hitReq_52_101 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h65;
  wire          compressDataVec_hitReq_53_101 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h65;
  wire          compressDataVec_hitReq_54_101 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h65;
  wire          compressDataVec_hitReq_55_101 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h65;
  wire          compressDataVec_hitReq_56_101 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h65;
  wire          compressDataVec_hitReq_57_101 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h65;
  wire          compressDataVec_hitReq_58_101 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h65;
  wire          compressDataVec_hitReq_59_101 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h65;
  wire          compressDataVec_hitReq_60_101 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h65;
  wire          compressDataVec_hitReq_61_101 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h65;
  wire          compressDataVec_hitReq_62_101 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h65;
  wire          compressDataVec_hitReq_63_101 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h65;
  wire [7:0]    compressDataVec_selectReqData_101 =
    (compressDataVec_hitReq_0_101 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_101 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_101 ? source2Pipe[23:16] : 8'h0)
    | (compressDataVec_hitReq_3_101 ? source2Pipe[31:24] : 8'h0) | (compressDataVec_hitReq_4_101 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_101 ? source2Pipe[47:40] : 8'h0)
    | (compressDataVec_hitReq_6_101 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_101 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_101 ? source2Pipe[71:64] : 8'h0)
    | (compressDataVec_hitReq_9_101 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_101 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_101 ? source2Pipe[95:88] : 8'h0)
    | (compressDataVec_hitReq_12_101 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_101 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_101 ? source2Pipe[119:112] : 8'h0)
    | (compressDataVec_hitReq_15_101 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_101 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_101 ? source2Pipe[143:136] : 8'h0)
    | (compressDataVec_hitReq_18_101 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_101 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_101 ? source2Pipe[167:160] : 8'h0)
    | (compressDataVec_hitReq_21_101 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_101 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_101 ? source2Pipe[191:184] : 8'h0)
    | (compressDataVec_hitReq_24_101 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_101 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_101 ? source2Pipe[215:208] : 8'h0)
    | (compressDataVec_hitReq_27_101 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_101 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_101 ? source2Pipe[239:232] : 8'h0)
    | (compressDataVec_hitReq_30_101 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_101 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_101 ? source2Pipe[263:256] : 8'h0)
    | (compressDataVec_hitReq_33_101 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_101 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_101 ? source2Pipe[287:280] : 8'h0)
    | (compressDataVec_hitReq_36_101 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_101 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_101 ? source2Pipe[311:304] : 8'h0)
    | (compressDataVec_hitReq_39_101 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_101 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_101 ? source2Pipe[335:328] : 8'h0)
    | (compressDataVec_hitReq_42_101 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_101 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_101 ? source2Pipe[359:352] : 8'h0)
    | (compressDataVec_hitReq_45_101 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_101 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_101 ? source2Pipe[383:376] : 8'h0)
    | (compressDataVec_hitReq_48_101 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_101 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_101 ? source2Pipe[407:400] : 8'h0)
    | (compressDataVec_hitReq_51_101 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_101 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_101 ? source2Pipe[431:424] : 8'h0)
    | (compressDataVec_hitReq_54_101 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_101 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_101 ? source2Pipe[455:448] : 8'h0)
    | (compressDataVec_hitReq_57_101 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_101 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_101 ? source2Pipe[479:472] : 8'h0)
    | (compressDataVec_hitReq_60_101 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_101 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_101 ? source2Pipe[503:496] : 8'h0)
    | (compressDataVec_hitReq_63_101 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_102 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h66;
  wire          compressDataVec_hitReq_1_102 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h66;
  wire          compressDataVec_hitReq_2_102 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h66;
  wire          compressDataVec_hitReq_3_102 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h66;
  wire          compressDataVec_hitReq_4_102 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h66;
  wire          compressDataVec_hitReq_5_102 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h66;
  wire          compressDataVec_hitReq_6_102 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h66;
  wire          compressDataVec_hitReq_7_102 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h66;
  wire          compressDataVec_hitReq_8_102 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h66;
  wire          compressDataVec_hitReq_9_102 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h66;
  wire          compressDataVec_hitReq_10_102 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h66;
  wire          compressDataVec_hitReq_11_102 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h66;
  wire          compressDataVec_hitReq_12_102 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h66;
  wire          compressDataVec_hitReq_13_102 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h66;
  wire          compressDataVec_hitReq_14_102 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h66;
  wire          compressDataVec_hitReq_15_102 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h66;
  wire          compressDataVec_hitReq_16_102 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h66;
  wire          compressDataVec_hitReq_17_102 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h66;
  wire          compressDataVec_hitReq_18_102 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h66;
  wire          compressDataVec_hitReq_19_102 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h66;
  wire          compressDataVec_hitReq_20_102 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h66;
  wire          compressDataVec_hitReq_21_102 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h66;
  wire          compressDataVec_hitReq_22_102 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h66;
  wire          compressDataVec_hitReq_23_102 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h66;
  wire          compressDataVec_hitReq_24_102 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h66;
  wire          compressDataVec_hitReq_25_102 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h66;
  wire          compressDataVec_hitReq_26_102 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h66;
  wire          compressDataVec_hitReq_27_102 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h66;
  wire          compressDataVec_hitReq_28_102 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h66;
  wire          compressDataVec_hitReq_29_102 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h66;
  wire          compressDataVec_hitReq_30_102 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h66;
  wire          compressDataVec_hitReq_31_102 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h66;
  wire          compressDataVec_hitReq_32_102 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h66;
  wire          compressDataVec_hitReq_33_102 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h66;
  wire          compressDataVec_hitReq_34_102 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h66;
  wire          compressDataVec_hitReq_35_102 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h66;
  wire          compressDataVec_hitReq_36_102 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h66;
  wire          compressDataVec_hitReq_37_102 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h66;
  wire          compressDataVec_hitReq_38_102 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h66;
  wire          compressDataVec_hitReq_39_102 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h66;
  wire          compressDataVec_hitReq_40_102 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h66;
  wire          compressDataVec_hitReq_41_102 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h66;
  wire          compressDataVec_hitReq_42_102 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h66;
  wire          compressDataVec_hitReq_43_102 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h66;
  wire          compressDataVec_hitReq_44_102 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h66;
  wire          compressDataVec_hitReq_45_102 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h66;
  wire          compressDataVec_hitReq_46_102 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h66;
  wire          compressDataVec_hitReq_47_102 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h66;
  wire          compressDataVec_hitReq_48_102 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h66;
  wire          compressDataVec_hitReq_49_102 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h66;
  wire          compressDataVec_hitReq_50_102 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h66;
  wire          compressDataVec_hitReq_51_102 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h66;
  wire          compressDataVec_hitReq_52_102 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h66;
  wire          compressDataVec_hitReq_53_102 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h66;
  wire          compressDataVec_hitReq_54_102 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h66;
  wire          compressDataVec_hitReq_55_102 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h66;
  wire          compressDataVec_hitReq_56_102 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h66;
  wire          compressDataVec_hitReq_57_102 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h66;
  wire          compressDataVec_hitReq_58_102 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h66;
  wire          compressDataVec_hitReq_59_102 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h66;
  wire          compressDataVec_hitReq_60_102 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h66;
  wire          compressDataVec_hitReq_61_102 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h66;
  wire          compressDataVec_hitReq_62_102 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h66;
  wire          compressDataVec_hitReq_63_102 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h66;
  wire [7:0]    compressDataVec_selectReqData_102 =
    (compressDataVec_hitReq_0_102 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_102 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_102 ? source2Pipe[23:16] : 8'h0)
    | (compressDataVec_hitReq_3_102 ? source2Pipe[31:24] : 8'h0) | (compressDataVec_hitReq_4_102 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_102 ? source2Pipe[47:40] : 8'h0)
    | (compressDataVec_hitReq_6_102 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_102 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_102 ? source2Pipe[71:64] : 8'h0)
    | (compressDataVec_hitReq_9_102 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_102 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_102 ? source2Pipe[95:88] : 8'h0)
    | (compressDataVec_hitReq_12_102 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_102 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_102 ? source2Pipe[119:112] : 8'h0)
    | (compressDataVec_hitReq_15_102 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_102 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_102 ? source2Pipe[143:136] : 8'h0)
    | (compressDataVec_hitReq_18_102 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_102 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_102 ? source2Pipe[167:160] : 8'h0)
    | (compressDataVec_hitReq_21_102 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_102 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_102 ? source2Pipe[191:184] : 8'h0)
    | (compressDataVec_hitReq_24_102 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_102 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_102 ? source2Pipe[215:208] : 8'h0)
    | (compressDataVec_hitReq_27_102 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_102 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_102 ? source2Pipe[239:232] : 8'h0)
    | (compressDataVec_hitReq_30_102 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_102 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_102 ? source2Pipe[263:256] : 8'h0)
    | (compressDataVec_hitReq_33_102 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_102 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_102 ? source2Pipe[287:280] : 8'h0)
    | (compressDataVec_hitReq_36_102 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_102 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_102 ? source2Pipe[311:304] : 8'h0)
    | (compressDataVec_hitReq_39_102 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_102 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_102 ? source2Pipe[335:328] : 8'h0)
    | (compressDataVec_hitReq_42_102 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_102 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_102 ? source2Pipe[359:352] : 8'h0)
    | (compressDataVec_hitReq_45_102 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_102 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_102 ? source2Pipe[383:376] : 8'h0)
    | (compressDataVec_hitReq_48_102 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_102 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_102 ? source2Pipe[407:400] : 8'h0)
    | (compressDataVec_hitReq_51_102 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_102 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_102 ? source2Pipe[431:424] : 8'h0)
    | (compressDataVec_hitReq_54_102 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_102 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_102 ? source2Pipe[455:448] : 8'h0)
    | (compressDataVec_hitReq_57_102 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_102 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_102 ? source2Pipe[479:472] : 8'h0)
    | (compressDataVec_hitReq_60_102 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_102 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_102 ? source2Pipe[503:496] : 8'h0)
    | (compressDataVec_hitReq_63_102 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_103 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h67;
  wire          compressDataVec_hitReq_1_103 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h67;
  wire          compressDataVec_hitReq_2_103 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h67;
  wire          compressDataVec_hitReq_3_103 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h67;
  wire          compressDataVec_hitReq_4_103 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h67;
  wire          compressDataVec_hitReq_5_103 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h67;
  wire          compressDataVec_hitReq_6_103 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h67;
  wire          compressDataVec_hitReq_7_103 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h67;
  wire          compressDataVec_hitReq_8_103 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h67;
  wire          compressDataVec_hitReq_9_103 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h67;
  wire          compressDataVec_hitReq_10_103 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h67;
  wire          compressDataVec_hitReq_11_103 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h67;
  wire          compressDataVec_hitReq_12_103 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h67;
  wire          compressDataVec_hitReq_13_103 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h67;
  wire          compressDataVec_hitReq_14_103 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h67;
  wire          compressDataVec_hitReq_15_103 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h67;
  wire          compressDataVec_hitReq_16_103 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h67;
  wire          compressDataVec_hitReq_17_103 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h67;
  wire          compressDataVec_hitReq_18_103 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h67;
  wire          compressDataVec_hitReq_19_103 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h67;
  wire          compressDataVec_hitReq_20_103 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h67;
  wire          compressDataVec_hitReq_21_103 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h67;
  wire          compressDataVec_hitReq_22_103 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h67;
  wire          compressDataVec_hitReq_23_103 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h67;
  wire          compressDataVec_hitReq_24_103 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h67;
  wire          compressDataVec_hitReq_25_103 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h67;
  wire          compressDataVec_hitReq_26_103 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h67;
  wire          compressDataVec_hitReq_27_103 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h67;
  wire          compressDataVec_hitReq_28_103 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h67;
  wire          compressDataVec_hitReq_29_103 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h67;
  wire          compressDataVec_hitReq_30_103 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h67;
  wire          compressDataVec_hitReq_31_103 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h67;
  wire          compressDataVec_hitReq_32_103 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h67;
  wire          compressDataVec_hitReq_33_103 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h67;
  wire          compressDataVec_hitReq_34_103 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h67;
  wire          compressDataVec_hitReq_35_103 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h67;
  wire          compressDataVec_hitReq_36_103 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h67;
  wire          compressDataVec_hitReq_37_103 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h67;
  wire          compressDataVec_hitReq_38_103 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h67;
  wire          compressDataVec_hitReq_39_103 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h67;
  wire          compressDataVec_hitReq_40_103 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h67;
  wire          compressDataVec_hitReq_41_103 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h67;
  wire          compressDataVec_hitReq_42_103 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h67;
  wire          compressDataVec_hitReq_43_103 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h67;
  wire          compressDataVec_hitReq_44_103 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h67;
  wire          compressDataVec_hitReq_45_103 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h67;
  wire          compressDataVec_hitReq_46_103 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h67;
  wire          compressDataVec_hitReq_47_103 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h67;
  wire          compressDataVec_hitReq_48_103 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h67;
  wire          compressDataVec_hitReq_49_103 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h67;
  wire          compressDataVec_hitReq_50_103 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h67;
  wire          compressDataVec_hitReq_51_103 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h67;
  wire          compressDataVec_hitReq_52_103 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h67;
  wire          compressDataVec_hitReq_53_103 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h67;
  wire          compressDataVec_hitReq_54_103 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h67;
  wire          compressDataVec_hitReq_55_103 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h67;
  wire          compressDataVec_hitReq_56_103 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h67;
  wire          compressDataVec_hitReq_57_103 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h67;
  wire          compressDataVec_hitReq_58_103 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h67;
  wire          compressDataVec_hitReq_59_103 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h67;
  wire          compressDataVec_hitReq_60_103 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h67;
  wire          compressDataVec_hitReq_61_103 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h67;
  wire          compressDataVec_hitReq_62_103 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h67;
  wire          compressDataVec_hitReq_63_103 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h67;
  wire [7:0]    compressDataVec_selectReqData_103 =
    (compressDataVec_hitReq_0_103 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_103 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_103 ? source2Pipe[23:16] : 8'h0)
    | (compressDataVec_hitReq_3_103 ? source2Pipe[31:24] : 8'h0) | (compressDataVec_hitReq_4_103 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_103 ? source2Pipe[47:40] : 8'h0)
    | (compressDataVec_hitReq_6_103 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_103 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_103 ? source2Pipe[71:64] : 8'h0)
    | (compressDataVec_hitReq_9_103 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_103 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_103 ? source2Pipe[95:88] : 8'h0)
    | (compressDataVec_hitReq_12_103 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_103 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_103 ? source2Pipe[119:112] : 8'h0)
    | (compressDataVec_hitReq_15_103 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_103 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_103 ? source2Pipe[143:136] : 8'h0)
    | (compressDataVec_hitReq_18_103 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_103 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_103 ? source2Pipe[167:160] : 8'h0)
    | (compressDataVec_hitReq_21_103 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_103 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_103 ? source2Pipe[191:184] : 8'h0)
    | (compressDataVec_hitReq_24_103 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_103 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_103 ? source2Pipe[215:208] : 8'h0)
    | (compressDataVec_hitReq_27_103 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_103 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_103 ? source2Pipe[239:232] : 8'h0)
    | (compressDataVec_hitReq_30_103 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_103 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_103 ? source2Pipe[263:256] : 8'h0)
    | (compressDataVec_hitReq_33_103 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_103 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_103 ? source2Pipe[287:280] : 8'h0)
    | (compressDataVec_hitReq_36_103 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_103 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_103 ? source2Pipe[311:304] : 8'h0)
    | (compressDataVec_hitReq_39_103 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_103 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_103 ? source2Pipe[335:328] : 8'h0)
    | (compressDataVec_hitReq_42_103 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_103 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_103 ? source2Pipe[359:352] : 8'h0)
    | (compressDataVec_hitReq_45_103 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_103 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_103 ? source2Pipe[383:376] : 8'h0)
    | (compressDataVec_hitReq_48_103 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_103 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_103 ? source2Pipe[407:400] : 8'h0)
    | (compressDataVec_hitReq_51_103 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_103 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_103 ? source2Pipe[431:424] : 8'h0)
    | (compressDataVec_hitReq_54_103 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_103 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_103 ? source2Pipe[455:448] : 8'h0)
    | (compressDataVec_hitReq_57_103 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_103 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_103 ? source2Pipe[479:472] : 8'h0)
    | (compressDataVec_hitReq_60_103 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_103 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_103 ? source2Pipe[503:496] : 8'h0)
    | (compressDataVec_hitReq_63_103 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_104 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h68;
  wire          compressDataVec_hitReq_1_104 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h68;
  wire          compressDataVec_hitReq_2_104 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h68;
  wire          compressDataVec_hitReq_3_104 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h68;
  wire          compressDataVec_hitReq_4_104 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h68;
  wire          compressDataVec_hitReq_5_104 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h68;
  wire          compressDataVec_hitReq_6_104 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h68;
  wire          compressDataVec_hitReq_7_104 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h68;
  wire          compressDataVec_hitReq_8_104 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h68;
  wire          compressDataVec_hitReq_9_104 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h68;
  wire          compressDataVec_hitReq_10_104 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h68;
  wire          compressDataVec_hitReq_11_104 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h68;
  wire          compressDataVec_hitReq_12_104 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h68;
  wire          compressDataVec_hitReq_13_104 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h68;
  wire          compressDataVec_hitReq_14_104 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h68;
  wire          compressDataVec_hitReq_15_104 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h68;
  wire          compressDataVec_hitReq_16_104 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h68;
  wire          compressDataVec_hitReq_17_104 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h68;
  wire          compressDataVec_hitReq_18_104 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h68;
  wire          compressDataVec_hitReq_19_104 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h68;
  wire          compressDataVec_hitReq_20_104 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h68;
  wire          compressDataVec_hitReq_21_104 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h68;
  wire          compressDataVec_hitReq_22_104 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h68;
  wire          compressDataVec_hitReq_23_104 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h68;
  wire          compressDataVec_hitReq_24_104 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h68;
  wire          compressDataVec_hitReq_25_104 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h68;
  wire          compressDataVec_hitReq_26_104 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h68;
  wire          compressDataVec_hitReq_27_104 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h68;
  wire          compressDataVec_hitReq_28_104 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h68;
  wire          compressDataVec_hitReq_29_104 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h68;
  wire          compressDataVec_hitReq_30_104 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h68;
  wire          compressDataVec_hitReq_31_104 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h68;
  wire          compressDataVec_hitReq_32_104 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h68;
  wire          compressDataVec_hitReq_33_104 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h68;
  wire          compressDataVec_hitReq_34_104 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h68;
  wire          compressDataVec_hitReq_35_104 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h68;
  wire          compressDataVec_hitReq_36_104 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h68;
  wire          compressDataVec_hitReq_37_104 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h68;
  wire          compressDataVec_hitReq_38_104 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h68;
  wire          compressDataVec_hitReq_39_104 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h68;
  wire          compressDataVec_hitReq_40_104 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h68;
  wire          compressDataVec_hitReq_41_104 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h68;
  wire          compressDataVec_hitReq_42_104 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h68;
  wire          compressDataVec_hitReq_43_104 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h68;
  wire          compressDataVec_hitReq_44_104 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h68;
  wire          compressDataVec_hitReq_45_104 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h68;
  wire          compressDataVec_hitReq_46_104 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h68;
  wire          compressDataVec_hitReq_47_104 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h68;
  wire          compressDataVec_hitReq_48_104 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h68;
  wire          compressDataVec_hitReq_49_104 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h68;
  wire          compressDataVec_hitReq_50_104 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h68;
  wire          compressDataVec_hitReq_51_104 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h68;
  wire          compressDataVec_hitReq_52_104 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h68;
  wire          compressDataVec_hitReq_53_104 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h68;
  wire          compressDataVec_hitReq_54_104 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h68;
  wire          compressDataVec_hitReq_55_104 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h68;
  wire          compressDataVec_hitReq_56_104 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h68;
  wire          compressDataVec_hitReq_57_104 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h68;
  wire          compressDataVec_hitReq_58_104 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h68;
  wire          compressDataVec_hitReq_59_104 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h68;
  wire          compressDataVec_hitReq_60_104 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h68;
  wire          compressDataVec_hitReq_61_104 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h68;
  wire          compressDataVec_hitReq_62_104 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h68;
  wire          compressDataVec_hitReq_63_104 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h68;
  wire [7:0]    compressDataVec_selectReqData_104 =
    (compressDataVec_hitReq_0_104 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_104 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_104 ? source2Pipe[23:16] : 8'h0)
    | (compressDataVec_hitReq_3_104 ? source2Pipe[31:24] : 8'h0) | (compressDataVec_hitReq_4_104 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_104 ? source2Pipe[47:40] : 8'h0)
    | (compressDataVec_hitReq_6_104 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_104 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_104 ? source2Pipe[71:64] : 8'h0)
    | (compressDataVec_hitReq_9_104 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_104 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_104 ? source2Pipe[95:88] : 8'h0)
    | (compressDataVec_hitReq_12_104 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_104 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_104 ? source2Pipe[119:112] : 8'h0)
    | (compressDataVec_hitReq_15_104 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_104 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_104 ? source2Pipe[143:136] : 8'h0)
    | (compressDataVec_hitReq_18_104 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_104 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_104 ? source2Pipe[167:160] : 8'h0)
    | (compressDataVec_hitReq_21_104 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_104 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_104 ? source2Pipe[191:184] : 8'h0)
    | (compressDataVec_hitReq_24_104 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_104 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_104 ? source2Pipe[215:208] : 8'h0)
    | (compressDataVec_hitReq_27_104 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_104 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_104 ? source2Pipe[239:232] : 8'h0)
    | (compressDataVec_hitReq_30_104 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_104 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_104 ? source2Pipe[263:256] : 8'h0)
    | (compressDataVec_hitReq_33_104 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_104 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_104 ? source2Pipe[287:280] : 8'h0)
    | (compressDataVec_hitReq_36_104 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_104 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_104 ? source2Pipe[311:304] : 8'h0)
    | (compressDataVec_hitReq_39_104 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_104 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_104 ? source2Pipe[335:328] : 8'h0)
    | (compressDataVec_hitReq_42_104 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_104 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_104 ? source2Pipe[359:352] : 8'h0)
    | (compressDataVec_hitReq_45_104 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_104 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_104 ? source2Pipe[383:376] : 8'h0)
    | (compressDataVec_hitReq_48_104 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_104 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_104 ? source2Pipe[407:400] : 8'h0)
    | (compressDataVec_hitReq_51_104 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_104 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_104 ? source2Pipe[431:424] : 8'h0)
    | (compressDataVec_hitReq_54_104 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_104 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_104 ? source2Pipe[455:448] : 8'h0)
    | (compressDataVec_hitReq_57_104 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_104 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_104 ? source2Pipe[479:472] : 8'h0)
    | (compressDataVec_hitReq_60_104 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_104 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_104 ? source2Pipe[503:496] : 8'h0)
    | (compressDataVec_hitReq_63_104 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_105 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h69;
  wire          compressDataVec_hitReq_1_105 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h69;
  wire          compressDataVec_hitReq_2_105 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h69;
  wire          compressDataVec_hitReq_3_105 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h69;
  wire          compressDataVec_hitReq_4_105 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h69;
  wire          compressDataVec_hitReq_5_105 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h69;
  wire          compressDataVec_hitReq_6_105 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h69;
  wire          compressDataVec_hitReq_7_105 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h69;
  wire          compressDataVec_hitReq_8_105 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h69;
  wire          compressDataVec_hitReq_9_105 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h69;
  wire          compressDataVec_hitReq_10_105 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h69;
  wire          compressDataVec_hitReq_11_105 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h69;
  wire          compressDataVec_hitReq_12_105 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h69;
  wire          compressDataVec_hitReq_13_105 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h69;
  wire          compressDataVec_hitReq_14_105 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h69;
  wire          compressDataVec_hitReq_15_105 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h69;
  wire          compressDataVec_hitReq_16_105 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h69;
  wire          compressDataVec_hitReq_17_105 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h69;
  wire          compressDataVec_hitReq_18_105 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h69;
  wire          compressDataVec_hitReq_19_105 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h69;
  wire          compressDataVec_hitReq_20_105 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h69;
  wire          compressDataVec_hitReq_21_105 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h69;
  wire          compressDataVec_hitReq_22_105 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h69;
  wire          compressDataVec_hitReq_23_105 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h69;
  wire          compressDataVec_hitReq_24_105 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h69;
  wire          compressDataVec_hitReq_25_105 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h69;
  wire          compressDataVec_hitReq_26_105 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h69;
  wire          compressDataVec_hitReq_27_105 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h69;
  wire          compressDataVec_hitReq_28_105 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h69;
  wire          compressDataVec_hitReq_29_105 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h69;
  wire          compressDataVec_hitReq_30_105 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h69;
  wire          compressDataVec_hitReq_31_105 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h69;
  wire          compressDataVec_hitReq_32_105 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h69;
  wire          compressDataVec_hitReq_33_105 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h69;
  wire          compressDataVec_hitReq_34_105 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h69;
  wire          compressDataVec_hitReq_35_105 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h69;
  wire          compressDataVec_hitReq_36_105 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h69;
  wire          compressDataVec_hitReq_37_105 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h69;
  wire          compressDataVec_hitReq_38_105 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h69;
  wire          compressDataVec_hitReq_39_105 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h69;
  wire          compressDataVec_hitReq_40_105 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h69;
  wire          compressDataVec_hitReq_41_105 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h69;
  wire          compressDataVec_hitReq_42_105 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h69;
  wire          compressDataVec_hitReq_43_105 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h69;
  wire          compressDataVec_hitReq_44_105 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h69;
  wire          compressDataVec_hitReq_45_105 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h69;
  wire          compressDataVec_hitReq_46_105 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h69;
  wire          compressDataVec_hitReq_47_105 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h69;
  wire          compressDataVec_hitReq_48_105 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h69;
  wire          compressDataVec_hitReq_49_105 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h69;
  wire          compressDataVec_hitReq_50_105 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h69;
  wire          compressDataVec_hitReq_51_105 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h69;
  wire          compressDataVec_hitReq_52_105 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h69;
  wire          compressDataVec_hitReq_53_105 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h69;
  wire          compressDataVec_hitReq_54_105 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h69;
  wire          compressDataVec_hitReq_55_105 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h69;
  wire          compressDataVec_hitReq_56_105 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h69;
  wire          compressDataVec_hitReq_57_105 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h69;
  wire          compressDataVec_hitReq_58_105 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h69;
  wire          compressDataVec_hitReq_59_105 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h69;
  wire          compressDataVec_hitReq_60_105 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h69;
  wire          compressDataVec_hitReq_61_105 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h69;
  wire          compressDataVec_hitReq_62_105 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h69;
  wire          compressDataVec_hitReq_63_105 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h69;
  wire [7:0]    compressDataVec_selectReqData_105 =
    (compressDataVec_hitReq_0_105 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_105 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_105 ? source2Pipe[23:16] : 8'h0)
    | (compressDataVec_hitReq_3_105 ? source2Pipe[31:24] : 8'h0) | (compressDataVec_hitReq_4_105 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_105 ? source2Pipe[47:40] : 8'h0)
    | (compressDataVec_hitReq_6_105 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_105 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_105 ? source2Pipe[71:64] : 8'h0)
    | (compressDataVec_hitReq_9_105 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_105 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_105 ? source2Pipe[95:88] : 8'h0)
    | (compressDataVec_hitReq_12_105 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_105 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_105 ? source2Pipe[119:112] : 8'h0)
    | (compressDataVec_hitReq_15_105 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_105 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_105 ? source2Pipe[143:136] : 8'h0)
    | (compressDataVec_hitReq_18_105 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_105 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_105 ? source2Pipe[167:160] : 8'h0)
    | (compressDataVec_hitReq_21_105 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_105 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_105 ? source2Pipe[191:184] : 8'h0)
    | (compressDataVec_hitReq_24_105 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_105 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_105 ? source2Pipe[215:208] : 8'h0)
    | (compressDataVec_hitReq_27_105 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_105 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_105 ? source2Pipe[239:232] : 8'h0)
    | (compressDataVec_hitReq_30_105 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_105 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_105 ? source2Pipe[263:256] : 8'h0)
    | (compressDataVec_hitReq_33_105 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_105 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_105 ? source2Pipe[287:280] : 8'h0)
    | (compressDataVec_hitReq_36_105 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_105 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_105 ? source2Pipe[311:304] : 8'h0)
    | (compressDataVec_hitReq_39_105 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_105 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_105 ? source2Pipe[335:328] : 8'h0)
    | (compressDataVec_hitReq_42_105 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_105 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_105 ? source2Pipe[359:352] : 8'h0)
    | (compressDataVec_hitReq_45_105 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_105 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_105 ? source2Pipe[383:376] : 8'h0)
    | (compressDataVec_hitReq_48_105 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_105 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_105 ? source2Pipe[407:400] : 8'h0)
    | (compressDataVec_hitReq_51_105 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_105 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_105 ? source2Pipe[431:424] : 8'h0)
    | (compressDataVec_hitReq_54_105 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_105 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_105 ? source2Pipe[455:448] : 8'h0)
    | (compressDataVec_hitReq_57_105 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_105 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_105 ? source2Pipe[479:472] : 8'h0)
    | (compressDataVec_hitReq_60_105 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_105 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_105 ? source2Pipe[503:496] : 8'h0)
    | (compressDataVec_hitReq_63_105 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_106 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h6A;
  wire          compressDataVec_hitReq_1_106 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h6A;
  wire          compressDataVec_hitReq_2_106 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h6A;
  wire          compressDataVec_hitReq_3_106 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h6A;
  wire          compressDataVec_hitReq_4_106 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h6A;
  wire          compressDataVec_hitReq_5_106 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h6A;
  wire          compressDataVec_hitReq_6_106 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h6A;
  wire          compressDataVec_hitReq_7_106 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h6A;
  wire          compressDataVec_hitReq_8_106 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h6A;
  wire          compressDataVec_hitReq_9_106 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h6A;
  wire          compressDataVec_hitReq_10_106 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h6A;
  wire          compressDataVec_hitReq_11_106 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h6A;
  wire          compressDataVec_hitReq_12_106 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h6A;
  wire          compressDataVec_hitReq_13_106 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h6A;
  wire          compressDataVec_hitReq_14_106 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h6A;
  wire          compressDataVec_hitReq_15_106 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h6A;
  wire          compressDataVec_hitReq_16_106 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h6A;
  wire          compressDataVec_hitReq_17_106 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h6A;
  wire          compressDataVec_hitReq_18_106 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h6A;
  wire          compressDataVec_hitReq_19_106 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h6A;
  wire          compressDataVec_hitReq_20_106 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h6A;
  wire          compressDataVec_hitReq_21_106 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h6A;
  wire          compressDataVec_hitReq_22_106 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h6A;
  wire          compressDataVec_hitReq_23_106 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h6A;
  wire          compressDataVec_hitReq_24_106 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h6A;
  wire          compressDataVec_hitReq_25_106 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h6A;
  wire          compressDataVec_hitReq_26_106 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h6A;
  wire          compressDataVec_hitReq_27_106 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h6A;
  wire          compressDataVec_hitReq_28_106 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h6A;
  wire          compressDataVec_hitReq_29_106 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h6A;
  wire          compressDataVec_hitReq_30_106 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h6A;
  wire          compressDataVec_hitReq_31_106 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h6A;
  wire          compressDataVec_hitReq_32_106 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h6A;
  wire          compressDataVec_hitReq_33_106 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h6A;
  wire          compressDataVec_hitReq_34_106 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h6A;
  wire          compressDataVec_hitReq_35_106 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h6A;
  wire          compressDataVec_hitReq_36_106 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h6A;
  wire          compressDataVec_hitReq_37_106 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h6A;
  wire          compressDataVec_hitReq_38_106 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h6A;
  wire          compressDataVec_hitReq_39_106 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h6A;
  wire          compressDataVec_hitReq_40_106 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h6A;
  wire          compressDataVec_hitReq_41_106 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h6A;
  wire          compressDataVec_hitReq_42_106 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h6A;
  wire          compressDataVec_hitReq_43_106 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h6A;
  wire          compressDataVec_hitReq_44_106 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h6A;
  wire          compressDataVec_hitReq_45_106 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h6A;
  wire          compressDataVec_hitReq_46_106 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h6A;
  wire          compressDataVec_hitReq_47_106 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h6A;
  wire          compressDataVec_hitReq_48_106 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h6A;
  wire          compressDataVec_hitReq_49_106 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h6A;
  wire          compressDataVec_hitReq_50_106 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h6A;
  wire          compressDataVec_hitReq_51_106 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h6A;
  wire          compressDataVec_hitReq_52_106 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h6A;
  wire          compressDataVec_hitReq_53_106 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h6A;
  wire          compressDataVec_hitReq_54_106 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h6A;
  wire          compressDataVec_hitReq_55_106 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h6A;
  wire          compressDataVec_hitReq_56_106 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h6A;
  wire          compressDataVec_hitReq_57_106 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h6A;
  wire          compressDataVec_hitReq_58_106 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h6A;
  wire          compressDataVec_hitReq_59_106 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h6A;
  wire          compressDataVec_hitReq_60_106 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h6A;
  wire          compressDataVec_hitReq_61_106 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h6A;
  wire          compressDataVec_hitReq_62_106 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h6A;
  wire          compressDataVec_hitReq_63_106 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h6A;
  wire [7:0]    compressDataVec_selectReqData_106 =
    (compressDataVec_hitReq_0_106 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_106 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_106 ? source2Pipe[23:16] : 8'h0)
    | (compressDataVec_hitReq_3_106 ? source2Pipe[31:24] : 8'h0) | (compressDataVec_hitReq_4_106 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_106 ? source2Pipe[47:40] : 8'h0)
    | (compressDataVec_hitReq_6_106 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_106 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_106 ? source2Pipe[71:64] : 8'h0)
    | (compressDataVec_hitReq_9_106 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_106 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_106 ? source2Pipe[95:88] : 8'h0)
    | (compressDataVec_hitReq_12_106 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_106 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_106 ? source2Pipe[119:112] : 8'h0)
    | (compressDataVec_hitReq_15_106 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_106 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_106 ? source2Pipe[143:136] : 8'h0)
    | (compressDataVec_hitReq_18_106 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_106 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_106 ? source2Pipe[167:160] : 8'h0)
    | (compressDataVec_hitReq_21_106 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_106 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_106 ? source2Pipe[191:184] : 8'h0)
    | (compressDataVec_hitReq_24_106 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_106 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_106 ? source2Pipe[215:208] : 8'h0)
    | (compressDataVec_hitReq_27_106 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_106 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_106 ? source2Pipe[239:232] : 8'h0)
    | (compressDataVec_hitReq_30_106 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_106 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_106 ? source2Pipe[263:256] : 8'h0)
    | (compressDataVec_hitReq_33_106 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_106 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_106 ? source2Pipe[287:280] : 8'h0)
    | (compressDataVec_hitReq_36_106 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_106 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_106 ? source2Pipe[311:304] : 8'h0)
    | (compressDataVec_hitReq_39_106 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_106 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_106 ? source2Pipe[335:328] : 8'h0)
    | (compressDataVec_hitReq_42_106 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_106 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_106 ? source2Pipe[359:352] : 8'h0)
    | (compressDataVec_hitReq_45_106 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_106 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_106 ? source2Pipe[383:376] : 8'h0)
    | (compressDataVec_hitReq_48_106 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_106 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_106 ? source2Pipe[407:400] : 8'h0)
    | (compressDataVec_hitReq_51_106 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_106 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_106 ? source2Pipe[431:424] : 8'h0)
    | (compressDataVec_hitReq_54_106 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_106 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_106 ? source2Pipe[455:448] : 8'h0)
    | (compressDataVec_hitReq_57_106 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_106 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_106 ? source2Pipe[479:472] : 8'h0)
    | (compressDataVec_hitReq_60_106 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_106 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_106 ? source2Pipe[503:496] : 8'h0)
    | (compressDataVec_hitReq_63_106 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_107 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h6B;
  wire          compressDataVec_hitReq_1_107 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h6B;
  wire          compressDataVec_hitReq_2_107 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h6B;
  wire          compressDataVec_hitReq_3_107 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h6B;
  wire          compressDataVec_hitReq_4_107 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h6B;
  wire          compressDataVec_hitReq_5_107 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h6B;
  wire          compressDataVec_hitReq_6_107 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h6B;
  wire          compressDataVec_hitReq_7_107 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h6B;
  wire          compressDataVec_hitReq_8_107 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h6B;
  wire          compressDataVec_hitReq_9_107 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h6B;
  wire          compressDataVec_hitReq_10_107 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h6B;
  wire          compressDataVec_hitReq_11_107 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h6B;
  wire          compressDataVec_hitReq_12_107 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h6B;
  wire          compressDataVec_hitReq_13_107 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h6B;
  wire          compressDataVec_hitReq_14_107 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h6B;
  wire          compressDataVec_hitReq_15_107 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h6B;
  wire          compressDataVec_hitReq_16_107 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h6B;
  wire          compressDataVec_hitReq_17_107 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h6B;
  wire          compressDataVec_hitReq_18_107 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h6B;
  wire          compressDataVec_hitReq_19_107 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h6B;
  wire          compressDataVec_hitReq_20_107 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h6B;
  wire          compressDataVec_hitReq_21_107 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h6B;
  wire          compressDataVec_hitReq_22_107 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h6B;
  wire          compressDataVec_hitReq_23_107 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h6B;
  wire          compressDataVec_hitReq_24_107 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h6B;
  wire          compressDataVec_hitReq_25_107 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h6B;
  wire          compressDataVec_hitReq_26_107 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h6B;
  wire          compressDataVec_hitReq_27_107 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h6B;
  wire          compressDataVec_hitReq_28_107 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h6B;
  wire          compressDataVec_hitReq_29_107 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h6B;
  wire          compressDataVec_hitReq_30_107 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h6B;
  wire          compressDataVec_hitReq_31_107 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h6B;
  wire          compressDataVec_hitReq_32_107 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h6B;
  wire          compressDataVec_hitReq_33_107 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h6B;
  wire          compressDataVec_hitReq_34_107 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h6B;
  wire          compressDataVec_hitReq_35_107 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h6B;
  wire          compressDataVec_hitReq_36_107 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h6B;
  wire          compressDataVec_hitReq_37_107 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h6B;
  wire          compressDataVec_hitReq_38_107 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h6B;
  wire          compressDataVec_hitReq_39_107 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h6B;
  wire          compressDataVec_hitReq_40_107 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h6B;
  wire          compressDataVec_hitReq_41_107 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h6B;
  wire          compressDataVec_hitReq_42_107 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h6B;
  wire          compressDataVec_hitReq_43_107 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h6B;
  wire          compressDataVec_hitReq_44_107 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h6B;
  wire          compressDataVec_hitReq_45_107 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h6B;
  wire          compressDataVec_hitReq_46_107 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h6B;
  wire          compressDataVec_hitReq_47_107 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h6B;
  wire          compressDataVec_hitReq_48_107 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h6B;
  wire          compressDataVec_hitReq_49_107 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h6B;
  wire          compressDataVec_hitReq_50_107 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h6B;
  wire          compressDataVec_hitReq_51_107 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h6B;
  wire          compressDataVec_hitReq_52_107 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h6B;
  wire          compressDataVec_hitReq_53_107 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h6B;
  wire          compressDataVec_hitReq_54_107 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h6B;
  wire          compressDataVec_hitReq_55_107 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h6B;
  wire          compressDataVec_hitReq_56_107 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h6B;
  wire          compressDataVec_hitReq_57_107 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h6B;
  wire          compressDataVec_hitReq_58_107 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h6B;
  wire          compressDataVec_hitReq_59_107 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h6B;
  wire          compressDataVec_hitReq_60_107 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h6B;
  wire          compressDataVec_hitReq_61_107 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h6B;
  wire          compressDataVec_hitReq_62_107 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h6B;
  wire          compressDataVec_hitReq_63_107 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h6B;
  wire [7:0]    compressDataVec_selectReqData_107 =
    (compressDataVec_hitReq_0_107 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_107 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_107 ? source2Pipe[23:16] : 8'h0)
    | (compressDataVec_hitReq_3_107 ? source2Pipe[31:24] : 8'h0) | (compressDataVec_hitReq_4_107 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_107 ? source2Pipe[47:40] : 8'h0)
    | (compressDataVec_hitReq_6_107 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_107 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_107 ? source2Pipe[71:64] : 8'h0)
    | (compressDataVec_hitReq_9_107 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_107 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_107 ? source2Pipe[95:88] : 8'h0)
    | (compressDataVec_hitReq_12_107 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_107 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_107 ? source2Pipe[119:112] : 8'h0)
    | (compressDataVec_hitReq_15_107 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_107 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_107 ? source2Pipe[143:136] : 8'h0)
    | (compressDataVec_hitReq_18_107 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_107 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_107 ? source2Pipe[167:160] : 8'h0)
    | (compressDataVec_hitReq_21_107 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_107 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_107 ? source2Pipe[191:184] : 8'h0)
    | (compressDataVec_hitReq_24_107 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_107 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_107 ? source2Pipe[215:208] : 8'h0)
    | (compressDataVec_hitReq_27_107 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_107 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_107 ? source2Pipe[239:232] : 8'h0)
    | (compressDataVec_hitReq_30_107 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_107 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_107 ? source2Pipe[263:256] : 8'h0)
    | (compressDataVec_hitReq_33_107 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_107 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_107 ? source2Pipe[287:280] : 8'h0)
    | (compressDataVec_hitReq_36_107 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_107 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_107 ? source2Pipe[311:304] : 8'h0)
    | (compressDataVec_hitReq_39_107 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_107 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_107 ? source2Pipe[335:328] : 8'h0)
    | (compressDataVec_hitReq_42_107 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_107 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_107 ? source2Pipe[359:352] : 8'h0)
    | (compressDataVec_hitReq_45_107 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_107 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_107 ? source2Pipe[383:376] : 8'h0)
    | (compressDataVec_hitReq_48_107 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_107 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_107 ? source2Pipe[407:400] : 8'h0)
    | (compressDataVec_hitReq_51_107 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_107 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_107 ? source2Pipe[431:424] : 8'h0)
    | (compressDataVec_hitReq_54_107 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_107 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_107 ? source2Pipe[455:448] : 8'h0)
    | (compressDataVec_hitReq_57_107 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_107 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_107 ? source2Pipe[479:472] : 8'h0)
    | (compressDataVec_hitReq_60_107 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_107 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_107 ? source2Pipe[503:496] : 8'h0)
    | (compressDataVec_hitReq_63_107 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_108 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h6C;
  wire          compressDataVec_hitReq_1_108 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h6C;
  wire          compressDataVec_hitReq_2_108 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h6C;
  wire          compressDataVec_hitReq_3_108 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h6C;
  wire          compressDataVec_hitReq_4_108 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h6C;
  wire          compressDataVec_hitReq_5_108 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h6C;
  wire          compressDataVec_hitReq_6_108 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h6C;
  wire          compressDataVec_hitReq_7_108 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h6C;
  wire          compressDataVec_hitReq_8_108 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h6C;
  wire          compressDataVec_hitReq_9_108 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h6C;
  wire          compressDataVec_hitReq_10_108 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h6C;
  wire          compressDataVec_hitReq_11_108 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h6C;
  wire          compressDataVec_hitReq_12_108 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h6C;
  wire          compressDataVec_hitReq_13_108 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h6C;
  wire          compressDataVec_hitReq_14_108 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h6C;
  wire          compressDataVec_hitReq_15_108 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h6C;
  wire          compressDataVec_hitReq_16_108 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h6C;
  wire          compressDataVec_hitReq_17_108 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h6C;
  wire          compressDataVec_hitReq_18_108 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h6C;
  wire          compressDataVec_hitReq_19_108 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h6C;
  wire          compressDataVec_hitReq_20_108 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h6C;
  wire          compressDataVec_hitReq_21_108 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h6C;
  wire          compressDataVec_hitReq_22_108 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h6C;
  wire          compressDataVec_hitReq_23_108 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h6C;
  wire          compressDataVec_hitReq_24_108 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h6C;
  wire          compressDataVec_hitReq_25_108 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h6C;
  wire          compressDataVec_hitReq_26_108 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h6C;
  wire          compressDataVec_hitReq_27_108 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h6C;
  wire          compressDataVec_hitReq_28_108 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h6C;
  wire          compressDataVec_hitReq_29_108 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h6C;
  wire          compressDataVec_hitReq_30_108 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h6C;
  wire          compressDataVec_hitReq_31_108 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h6C;
  wire          compressDataVec_hitReq_32_108 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h6C;
  wire          compressDataVec_hitReq_33_108 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h6C;
  wire          compressDataVec_hitReq_34_108 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h6C;
  wire          compressDataVec_hitReq_35_108 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h6C;
  wire          compressDataVec_hitReq_36_108 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h6C;
  wire          compressDataVec_hitReq_37_108 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h6C;
  wire          compressDataVec_hitReq_38_108 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h6C;
  wire          compressDataVec_hitReq_39_108 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h6C;
  wire          compressDataVec_hitReq_40_108 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h6C;
  wire          compressDataVec_hitReq_41_108 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h6C;
  wire          compressDataVec_hitReq_42_108 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h6C;
  wire          compressDataVec_hitReq_43_108 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h6C;
  wire          compressDataVec_hitReq_44_108 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h6C;
  wire          compressDataVec_hitReq_45_108 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h6C;
  wire          compressDataVec_hitReq_46_108 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h6C;
  wire          compressDataVec_hitReq_47_108 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h6C;
  wire          compressDataVec_hitReq_48_108 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h6C;
  wire          compressDataVec_hitReq_49_108 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h6C;
  wire          compressDataVec_hitReq_50_108 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h6C;
  wire          compressDataVec_hitReq_51_108 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h6C;
  wire          compressDataVec_hitReq_52_108 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h6C;
  wire          compressDataVec_hitReq_53_108 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h6C;
  wire          compressDataVec_hitReq_54_108 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h6C;
  wire          compressDataVec_hitReq_55_108 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h6C;
  wire          compressDataVec_hitReq_56_108 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h6C;
  wire          compressDataVec_hitReq_57_108 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h6C;
  wire          compressDataVec_hitReq_58_108 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h6C;
  wire          compressDataVec_hitReq_59_108 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h6C;
  wire          compressDataVec_hitReq_60_108 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h6C;
  wire          compressDataVec_hitReq_61_108 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h6C;
  wire          compressDataVec_hitReq_62_108 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h6C;
  wire          compressDataVec_hitReq_63_108 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h6C;
  wire [7:0]    compressDataVec_selectReqData_108 =
    (compressDataVec_hitReq_0_108 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_108 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_108 ? source2Pipe[23:16] : 8'h0)
    | (compressDataVec_hitReq_3_108 ? source2Pipe[31:24] : 8'h0) | (compressDataVec_hitReq_4_108 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_108 ? source2Pipe[47:40] : 8'h0)
    | (compressDataVec_hitReq_6_108 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_108 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_108 ? source2Pipe[71:64] : 8'h0)
    | (compressDataVec_hitReq_9_108 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_108 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_108 ? source2Pipe[95:88] : 8'h0)
    | (compressDataVec_hitReq_12_108 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_108 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_108 ? source2Pipe[119:112] : 8'h0)
    | (compressDataVec_hitReq_15_108 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_108 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_108 ? source2Pipe[143:136] : 8'h0)
    | (compressDataVec_hitReq_18_108 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_108 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_108 ? source2Pipe[167:160] : 8'h0)
    | (compressDataVec_hitReq_21_108 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_108 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_108 ? source2Pipe[191:184] : 8'h0)
    | (compressDataVec_hitReq_24_108 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_108 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_108 ? source2Pipe[215:208] : 8'h0)
    | (compressDataVec_hitReq_27_108 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_108 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_108 ? source2Pipe[239:232] : 8'h0)
    | (compressDataVec_hitReq_30_108 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_108 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_108 ? source2Pipe[263:256] : 8'h0)
    | (compressDataVec_hitReq_33_108 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_108 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_108 ? source2Pipe[287:280] : 8'h0)
    | (compressDataVec_hitReq_36_108 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_108 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_108 ? source2Pipe[311:304] : 8'h0)
    | (compressDataVec_hitReq_39_108 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_108 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_108 ? source2Pipe[335:328] : 8'h0)
    | (compressDataVec_hitReq_42_108 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_108 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_108 ? source2Pipe[359:352] : 8'h0)
    | (compressDataVec_hitReq_45_108 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_108 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_108 ? source2Pipe[383:376] : 8'h0)
    | (compressDataVec_hitReq_48_108 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_108 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_108 ? source2Pipe[407:400] : 8'h0)
    | (compressDataVec_hitReq_51_108 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_108 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_108 ? source2Pipe[431:424] : 8'h0)
    | (compressDataVec_hitReq_54_108 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_108 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_108 ? source2Pipe[455:448] : 8'h0)
    | (compressDataVec_hitReq_57_108 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_108 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_108 ? source2Pipe[479:472] : 8'h0)
    | (compressDataVec_hitReq_60_108 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_108 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_108 ? source2Pipe[503:496] : 8'h0)
    | (compressDataVec_hitReq_63_108 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_109 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h6D;
  wire          compressDataVec_hitReq_1_109 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h6D;
  wire          compressDataVec_hitReq_2_109 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h6D;
  wire          compressDataVec_hitReq_3_109 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h6D;
  wire          compressDataVec_hitReq_4_109 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h6D;
  wire          compressDataVec_hitReq_5_109 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h6D;
  wire          compressDataVec_hitReq_6_109 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h6D;
  wire          compressDataVec_hitReq_7_109 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h6D;
  wire          compressDataVec_hitReq_8_109 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h6D;
  wire          compressDataVec_hitReq_9_109 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h6D;
  wire          compressDataVec_hitReq_10_109 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h6D;
  wire          compressDataVec_hitReq_11_109 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h6D;
  wire          compressDataVec_hitReq_12_109 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h6D;
  wire          compressDataVec_hitReq_13_109 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h6D;
  wire          compressDataVec_hitReq_14_109 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h6D;
  wire          compressDataVec_hitReq_15_109 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h6D;
  wire          compressDataVec_hitReq_16_109 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h6D;
  wire          compressDataVec_hitReq_17_109 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h6D;
  wire          compressDataVec_hitReq_18_109 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h6D;
  wire          compressDataVec_hitReq_19_109 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h6D;
  wire          compressDataVec_hitReq_20_109 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h6D;
  wire          compressDataVec_hitReq_21_109 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h6D;
  wire          compressDataVec_hitReq_22_109 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h6D;
  wire          compressDataVec_hitReq_23_109 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h6D;
  wire          compressDataVec_hitReq_24_109 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h6D;
  wire          compressDataVec_hitReq_25_109 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h6D;
  wire          compressDataVec_hitReq_26_109 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h6D;
  wire          compressDataVec_hitReq_27_109 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h6D;
  wire          compressDataVec_hitReq_28_109 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h6D;
  wire          compressDataVec_hitReq_29_109 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h6D;
  wire          compressDataVec_hitReq_30_109 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h6D;
  wire          compressDataVec_hitReq_31_109 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h6D;
  wire          compressDataVec_hitReq_32_109 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h6D;
  wire          compressDataVec_hitReq_33_109 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h6D;
  wire          compressDataVec_hitReq_34_109 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h6D;
  wire          compressDataVec_hitReq_35_109 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h6D;
  wire          compressDataVec_hitReq_36_109 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h6D;
  wire          compressDataVec_hitReq_37_109 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h6D;
  wire          compressDataVec_hitReq_38_109 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h6D;
  wire          compressDataVec_hitReq_39_109 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h6D;
  wire          compressDataVec_hitReq_40_109 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h6D;
  wire          compressDataVec_hitReq_41_109 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h6D;
  wire          compressDataVec_hitReq_42_109 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h6D;
  wire          compressDataVec_hitReq_43_109 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h6D;
  wire          compressDataVec_hitReq_44_109 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h6D;
  wire          compressDataVec_hitReq_45_109 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h6D;
  wire          compressDataVec_hitReq_46_109 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h6D;
  wire          compressDataVec_hitReq_47_109 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h6D;
  wire          compressDataVec_hitReq_48_109 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h6D;
  wire          compressDataVec_hitReq_49_109 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h6D;
  wire          compressDataVec_hitReq_50_109 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h6D;
  wire          compressDataVec_hitReq_51_109 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h6D;
  wire          compressDataVec_hitReq_52_109 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h6D;
  wire          compressDataVec_hitReq_53_109 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h6D;
  wire          compressDataVec_hitReq_54_109 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h6D;
  wire          compressDataVec_hitReq_55_109 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h6D;
  wire          compressDataVec_hitReq_56_109 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h6D;
  wire          compressDataVec_hitReq_57_109 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h6D;
  wire          compressDataVec_hitReq_58_109 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h6D;
  wire          compressDataVec_hitReq_59_109 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h6D;
  wire          compressDataVec_hitReq_60_109 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h6D;
  wire          compressDataVec_hitReq_61_109 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h6D;
  wire          compressDataVec_hitReq_62_109 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h6D;
  wire          compressDataVec_hitReq_63_109 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h6D;
  wire [7:0]    compressDataVec_selectReqData_109 =
    (compressDataVec_hitReq_0_109 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_109 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_109 ? source2Pipe[23:16] : 8'h0)
    | (compressDataVec_hitReq_3_109 ? source2Pipe[31:24] : 8'h0) | (compressDataVec_hitReq_4_109 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_109 ? source2Pipe[47:40] : 8'h0)
    | (compressDataVec_hitReq_6_109 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_109 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_109 ? source2Pipe[71:64] : 8'h0)
    | (compressDataVec_hitReq_9_109 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_109 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_109 ? source2Pipe[95:88] : 8'h0)
    | (compressDataVec_hitReq_12_109 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_109 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_109 ? source2Pipe[119:112] : 8'h0)
    | (compressDataVec_hitReq_15_109 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_109 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_109 ? source2Pipe[143:136] : 8'h0)
    | (compressDataVec_hitReq_18_109 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_109 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_109 ? source2Pipe[167:160] : 8'h0)
    | (compressDataVec_hitReq_21_109 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_109 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_109 ? source2Pipe[191:184] : 8'h0)
    | (compressDataVec_hitReq_24_109 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_109 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_109 ? source2Pipe[215:208] : 8'h0)
    | (compressDataVec_hitReq_27_109 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_109 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_109 ? source2Pipe[239:232] : 8'h0)
    | (compressDataVec_hitReq_30_109 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_109 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_109 ? source2Pipe[263:256] : 8'h0)
    | (compressDataVec_hitReq_33_109 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_109 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_109 ? source2Pipe[287:280] : 8'h0)
    | (compressDataVec_hitReq_36_109 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_109 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_109 ? source2Pipe[311:304] : 8'h0)
    | (compressDataVec_hitReq_39_109 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_109 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_109 ? source2Pipe[335:328] : 8'h0)
    | (compressDataVec_hitReq_42_109 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_109 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_109 ? source2Pipe[359:352] : 8'h0)
    | (compressDataVec_hitReq_45_109 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_109 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_109 ? source2Pipe[383:376] : 8'h0)
    | (compressDataVec_hitReq_48_109 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_109 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_109 ? source2Pipe[407:400] : 8'h0)
    | (compressDataVec_hitReq_51_109 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_109 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_109 ? source2Pipe[431:424] : 8'h0)
    | (compressDataVec_hitReq_54_109 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_109 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_109 ? source2Pipe[455:448] : 8'h0)
    | (compressDataVec_hitReq_57_109 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_109 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_109 ? source2Pipe[479:472] : 8'h0)
    | (compressDataVec_hitReq_60_109 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_109 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_109 ? source2Pipe[503:496] : 8'h0)
    | (compressDataVec_hitReq_63_109 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_110 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h6E;
  wire          compressDataVec_hitReq_1_110 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h6E;
  wire          compressDataVec_hitReq_2_110 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h6E;
  wire          compressDataVec_hitReq_3_110 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h6E;
  wire          compressDataVec_hitReq_4_110 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h6E;
  wire          compressDataVec_hitReq_5_110 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h6E;
  wire          compressDataVec_hitReq_6_110 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h6E;
  wire          compressDataVec_hitReq_7_110 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h6E;
  wire          compressDataVec_hitReq_8_110 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h6E;
  wire          compressDataVec_hitReq_9_110 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h6E;
  wire          compressDataVec_hitReq_10_110 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h6E;
  wire          compressDataVec_hitReq_11_110 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h6E;
  wire          compressDataVec_hitReq_12_110 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h6E;
  wire          compressDataVec_hitReq_13_110 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h6E;
  wire          compressDataVec_hitReq_14_110 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h6E;
  wire          compressDataVec_hitReq_15_110 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h6E;
  wire          compressDataVec_hitReq_16_110 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h6E;
  wire          compressDataVec_hitReq_17_110 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h6E;
  wire          compressDataVec_hitReq_18_110 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h6E;
  wire          compressDataVec_hitReq_19_110 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h6E;
  wire          compressDataVec_hitReq_20_110 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h6E;
  wire          compressDataVec_hitReq_21_110 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h6E;
  wire          compressDataVec_hitReq_22_110 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h6E;
  wire          compressDataVec_hitReq_23_110 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h6E;
  wire          compressDataVec_hitReq_24_110 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h6E;
  wire          compressDataVec_hitReq_25_110 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h6E;
  wire          compressDataVec_hitReq_26_110 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h6E;
  wire          compressDataVec_hitReq_27_110 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h6E;
  wire          compressDataVec_hitReq_28_110 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h6E;
  wire          compressDataVec_hitReq_29_110 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h6E;
  wire          compressDataVec_hitReq_30_110 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h6E;
  wire          compressDataVec_hitReq_31_110 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h6E;
  wire          compressDataVec_hitReq_32_110 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h6E;
  wire          compressDataVec_hitReq_33_110 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h6E;
  wire          compressDataVec_hitReq_34_110 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h6E;
  wire          compressDataVec_hitReq_35_110 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h6E;
  wire          compressDataVec_hitReq_36_110 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h6E;
  wire          compressDataVec_hitReq_37_110 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h6E;
  wire          compressDataVec_hitReq_38_110 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h6E;
  wire          compressDataVec_hitReq_39_110 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h6E;
  wire          compressDataVec_hitReq_40_110 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h6E;
  wire          compressDataVec_hitReq_41_110 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h6E;
  wire          compressDataVec_hitReq_42_110 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h6E;
  wire          compressDataVec_hitReq_43_110 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h6E;
  wire          compressDataVec_hitReq_44_110 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h6E;
  wire          compressDataVec_hitReq_45_110 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h6E;
  wire          compressDataVec_hitReq_46_110 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h6E;
  wire          compressDataVec_hitReq_47_110 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h6E;
  wire          compressDataVec_hitReq_48_110 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h6E;
  wire          compressDataVec_hitReq_49_110 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h6E;
  wire          compressDataVec_hitReq_50_110 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h6E;
  wire          compressDataVec_hitReq_51_110 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h6E;
  wire          compressDataVec_hitReq_52_110 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h6E;
  wire          compressDataVec_hitReq_53_110 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h6E;
  wire          compressDataVec_hitReq_54_110 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h6E;
  wire          compressDataVec_hitReq_55_110 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h6E;
  wire          compressDataVec_hitReq_56_110 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h6E;
  wire          compressDataVec_hitReq_57_110 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h6E;
  wire          compressDataVec_hitReq_58_110 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h6E;
  wire          compressDataVec_hitReq_59_110 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h6E;
  wire          compressDataVec_hitReq_60_110 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h6E;
  wire          compressDataVec_hitReq_61_110 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h6E;
  wire          compressDataVec_hitReq_62_110 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h6E;
  wire          compressDataVec_hitReq_63_110 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h6E;
  wire [7:0]    compressDataVec_selectReqData_110 =
    (compressDataVec_hitReq_0_110 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_110 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_110 ? source2Pipe[23:16] : 8'h0)
    | (compressDataVec_hitReq_3_110 ? source2Pipe[31:24] : 8'h0) | (compressDataVec_hitReq_4_110 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_110 ? source2Pipe[47:40] : 8'h0)
    | (compressDataVec_hitReq_6_110 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_110 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_110 ? source2Pipe[71:64] : 8'h0)
    | (compressDataVec_hitReq_9_110 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_110 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_110 ? source2Pipe[95:88] : 8'h0)
    | (compressDataVec_hitReq_12_110 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_110 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_110 ? source2Pipe[119:112] : 8'h0)
    | (compressDataVec_hitReq_15_110 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_110 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_110 ? source2Pipe[143:136] : 8'h0)
    | (compressDataVec_hitReq_18_110 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_110 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_110 ? source2Pipe[167:160] : 8'h0)
    | (compressDataVec_hitReq_21_110 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_110 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_110 ? source2Pipe[191:184] : 8'h0)
    | (compressDataVec_hitReq_24_110 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_110 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_110 ? source2Pipe[215:208] : 8'h0)
    | (compressDataVec_hitReq_27_110 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_110 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_110 ? source2Pipe[239:232] : 8'h0)
    | (compressDataVec_hitReq_30_110 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_110 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_110 ? source2Pipe[263:256] : 8'h0)
    | (compressDataVec_hitReq_33_110 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_110 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_110 ? source2Pipe[287:280] : 8'h0)
    | (compressDataVec_hitReq_36_110 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_110 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_110 ? source2Pipe[311:304] : 8'h0)
    | (compressDataVec_hitReq_39_110 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_110 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_110 ? source2Pipe[335:328] : 8'h0)
    | (compressDataVec_hitReq_42_110 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_110 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_110 ? source2Pipe[359:352] : 8'h0)
    | (compressDataVec_hitReq_45_110 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_110 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_110 ? source2Pipe[383:376] : 8'h0)
    | (compressDataVec_hitReq_48_110 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_110 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_110 ? source2Pipe[407:400] : 8'h0)
    | (compressDataVec_hitReq_51_110 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_110 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_110 ? source2Pipe[431:424] : 8'h0)
    | (compressDataVec_hitReq_54_110 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_110 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_110 ? source2Pipe[455:448] : 8'h0)
    | (compressDataVec_hitReq_57_110 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_110 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_110 ? source2Pipe[479:472] : 8'h0)
    | (compressDataVec_hitReq_60_110 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_110 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_110 ? source2Pipe[503:496] : 8'h0)
    | (compressDataVec_hitReq_63_110 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_111 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h6F;
  wire          compressDataVec_hitReq_1_111 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h6F;
  wire          compressDataVec_hitReq_2_111 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h6F;
  wire          compressDataVec_hitReq_3_111 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h6F;
  wire          compressDataVec_hitReq_4_111 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h6F;
  wire          compressDataVec_hitReq_5_111 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h6F;
  wire          compressDataVec_hitReq_6_111 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h6F;
  wire          compressDataVec_hitReq_7_111 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h6F;
  wire          compressDataVec_hitReq_8_111 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h6F;
  wire          compressDataVec_hitReq_9_111 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h6F;
  wire          compressDataVec_hitReq_10_111 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h6F;
  wire          compressDataVec_hitReq_11_111 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h6F;
  wire          compressDataVec_hitReq_12_111 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h6F;
  wire          compressDataVec_hitReq_13_111 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h6F;
  wire          compressDataVec_hitReq_14_111 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h6F;
  wire          compressDataVec_hitReq_15_111 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h6F;
  wire          compressDataVec_hitReq_16_111 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h6F;
  wire          compressDataVec_hitReq_17_111 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h6F;
  wire          compressDataVec_hitReq_18_111 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h6F;
  wire          compressDataVec_hitReq_19_111 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h6F;
  wire          compressDataVec_hitReq_20_111 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h6F;
  wire          compressDataVec_hitReq_21_111 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h6F;
  wire          compressDataVec_hitReq_22_111 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h6F;
  wire          compressDataVec_hitReq_23_111 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h6F;
  wire          compressDataVec_hitReq_24_111 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h6F;
  wire          compressDataVec_hitReq_25_111 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h6F;
  wire          compressDataVec_hitReq_26_111 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h6F;
  wire          compressDataVec_hitReq_27_111 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h6F;
  wire          compressDataVec_hitReq_28_111 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h6F;
  wire          compressDataVec_hitReq_29_111 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h6F;
  wire          compressDataVec_hitReq_30_111 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h6F;
  wire          compressDataVec_hitReq_31_111 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h6F;
  wire          compressDataVec_hitReq_32_111 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h6F;
  wire          compressDataVec_hitReq_33_111 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h6F;
  wire          compressDataVec_hitReq_34_111 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h6F;
  wire          compressDataVec_hitReq_35_111 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h6F;
  wire          compressDataVec_hitReq_36_111 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h6F;
  wire          compressDataVec_hitReq_37_111 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h6F;
  wire          compressDataVec_hitReq_38_111 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h6F;
  wire          compressDataVec_hitReq_39_111 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h6F;
  wire          compressDataVec_hitReq_40_111 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h6F;
  wire          compressDataVec_hitReq_41_111 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h6F;
  wire          compressDataVec_hitReq_42_111 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h6F;
  wire          compressDataVec_hitReq_43_111 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h6F;
  wire          compressDataVec_hitReq_44_111 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h6F;
  wire          compressDataVec_hitReq_45_111 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h6F;
  wire          compressDataVec_hitReq_46_111 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h6F;
  wire          compressDataVec_hitReq_47_111 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h6F;
  wire          compressDataVec_hitReq_48_111 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h6F;
  wire          compressDataVec_hitReq_49_111 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h6F;
  wire          compressDataVec_hitReq_50_111 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h6F;
  wire          compressDataVec_hitReq_51_111 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h6F;
  wire          compressDataVec_hitReq_52_111 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h6F;
  wire          compressDataVec_hitReq_53_111 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h6F;
  wire          compressDataVec_hitReq_54_111 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h6F;
  wire          compressDataVec_hitReq_55_111 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h6F;
  wire          compressDataVec_hitReq_56_111 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h6F;
  wire          compressDataVec_hitReq_57_111 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h6F;
  wire          compressDataVec_hitReq_58_111 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h6F;
  wire          compressDataVec_hitReq_59_111 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h6F;
  wire          compressDataVec_hitReq_60_111 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h6F;
  wire          compressDataVec_hitReq_61_111 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h6F;
  wire          compressDataVec_hitReq_62_111 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h6F;
  wire          compressDataVec_hitReq_63_111 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h6F;
  wire [7:0]    compressDataVec_selectReqData_111 =
    (compressDataVec_hitReq_0_111 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_111 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_111 ? source2Pipe[23:16] : 8'h0)
    | (compressDataVec_hitReq_3_111 ? source2Pipe[31:24] : 8'h0) | (compressDataVec_hitReq_4_111 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_111 ? source2Pipe[47:40] : 8'h0)
    | (compressDataVec_hitReq_6_111 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_111 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_111 ? source2Pipe[71:64] : 8'h0)
    | (compressDataVec_hitReq_9_111 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_111 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_111 ? source2Pipe[95:88] : 8'h0)
    | (compressDataVec_hitReq_12_111 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_111 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_111 ? source2Pipe[119:112] : 8'h0)
    | (compressDataVec_hitReq_15_111 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_111 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_111 ? source2Pipe[143:136] : 8'h0)
    | (compressDataVec_hitReq_18_111 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_111 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_111 ? source2Pipe[167:160] : 8'h0)
    | (compressDataVec_hitReq_21_111 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_111 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_111 ? source2Pipe[191:184] : 8'h0)
    | (compressDataVec_hitReq_24_111 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_111 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_111 ? source2Pipe[215:208] : 8'h0)
    | (compressDataVec_hitReq_27_111 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_111 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_111 ? source2Pipe[239:232] : 8'h0)
    | (compressDataVec_hitReq_30_111 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_111 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_111 ? source2Pipe[263:256] : 8'h0)
    | (compressDataVec_hitReq_33_111 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_111 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_111 ? source2Pipe[287:280] : 8'h0)
    | (compressDataVec_hitReq_36_111 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_111 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_111 ? source2Pipe[311:304] : 8'h0)
    | (compressDataVec_hitReq_39_111 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_111 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_111 ? source2Pipe[335:328] : 8'h0)
    | (compressDataVec_hitReq_42_111 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_111 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_111 ? source2Pipe[359:352] : 8'h0)
    | (compressDataVec_hitReq_45_111 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_111 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_111 ? source2Pipe[383:376] : 8'h0)
    | (compressDataVec_hitReq_48_111 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_111 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_111 ? source2Pipe[407:400] : 8'h0)
    | (compressDataVec_hitReq_51_111 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_111 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_111 ? source2Pipe[431:424] : 8'h0)
    | (compressDataVec_hitReq_54_111 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_111 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_111 ? source2Pipe[455:448] : 8'h0)
    | (compressDataVec_hitReq_57_111 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_111 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_111 ? source2Pipe[479:472] : 8'h0)
    | (compressDataVec_hitReq_60_111 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_111 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_111 ? source2Pipe[503:496] : 8'h0)
    | (compressDataVec_hitReq_63_111 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_112 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h70;
  wire          compressDataVec_hitReq_1_112 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h70;
  wire          compressDataVec_hitReq_2_112 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h70;
  wire          compressDataVec_hitReq_3_112 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h70;
  wire          compressDataVec_hitReq_4_112 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h70;
  wire          compressDataVec_hitReq_5_112 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h70;
  wire          compressDataVec_hitReq_6_112 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h70;
  wire          compressDataVec_hitReq_7_112 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h70;
  wire          compressDataVec_hitReq_8_112 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h70;
  wire          compressDataVec_hitReq_9_112 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h70;
  wire          compressDataVec_hitReq_10_112 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h70;
  wire          compressDataVec_hitReq_11_112 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h70;
  wire          compressDataVec_hitReq_12_112 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h70;
  wire          compressDataVec_hitReq_13_112 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h70;
  wire          compressDataVec_hitReq_14_112 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h70;
  wire          compressDataVec_hitReq_15_112 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h70;
  wire          compressDataVec_hitReq_16_112 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h70;
  wire          compressDataVec_hitReq_17_112 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h70;
  wire          compressDataVec_hitReq_18_112 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h70;
  wire          compressDataVec_hitReq_19_112 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h70;
  wire          compressDataVec_hitReq_20_112 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h70;
  wire          compressDataVec_hitReq_21_112 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h70;
  wire          compressDataVec_hitReq_22_112 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h70;
  wire          compressDataVec_hitReq_23_112 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h70;
  wire          compressDataVec_hitReq_24_112 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h70;
  wire          compressDataVec_hitReq_25_112 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h70;
  wire          compressDataVec_hitReq_26_112 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h70;
  wire          compressDataVec_hitReq_27_112 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h70;
  wire          compressDataVec_hitReq_28_112 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h70;
  wire          compressDataVec_hitReq_29_112 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h70;
  wire          compressDataVec_hitReq_30_112 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h70;
  wire          compressDataVec_hitReq_31_112 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h70;
  wire          compressDataVec_hitReq_32_112 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h70;
  wire          compressDataVec_hitReq_33_112 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h70;
  wire          compressDataVec_hitReq_34_112 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h70;
  wire          compressDataVec_hitReq_35_112 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h70;
  wire          compressDataVec_hitReq_36_112 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h70;
  wire          compressDataVec_hitReq_37_112 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h70;
  wire          compressDataVec_hitReq_38_112 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h70;
  wire          compressDataVec_hitReq_39_112 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h70;
  wire          compressDataVec_hitReq_40_112 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h70;
  wire          compressDataVec_hitReq_41_112 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h70;
  wire          compressDataVec_hitReq_42_112 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h70;
  wire          compressDataVec_hitReq_43_112 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h70;
  wire          compressDataVec_hitReq_44_112 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h70;
  wire          compressDataVec_hitReq_45_112 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h70;
  wire          compressDataVec_hitReq_46_112 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h70;
  wire          compressDataVec_hitReq_47_112 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h70;
  wire          compressDataVec_hitReq_48_112 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h70;
  wire          compressDataVec_hitReq_49_112 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h70;
  wire          compressDataVec_hitReq_50_112 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h70;
  wire          compressDataVec_hitReq_51_112 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h70;
  wire          compressDataVec_hitReq_52_112 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h70;
  wire          compressDataVec_hitReq_53_112 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h70;
  wire          compressDataVec_hitReq_54_112 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h70;
  wire          compressDataVec_hitReq_55_112 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h70;
  wire          compressDataVec_hitReq_56_112 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h70;
  wire          compressDataVec_hitReq_57_112 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h70;
  wire          compressDataVec_hitReq_58_112 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h70;
  wire          compressDataVec_hitReq_59_112 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h70;
  wire          compressDataVec_hitReq_60_112 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h70;
  wire          compressDataVec_hitReq_61_112 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h70;
  wire          compressDataVec_hitReq_62_112 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h70;
  wire          compressDataVec_hitReq_63_112 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h70;
  wire [7:0]    compressDataVec_selectReqData_112 =
    (compressDataVec_hitReq_0_112 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_112 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_112 ? source2Pipe[23:16] : 8'h0)
    | (compressDataVec_hitReq_3_112 ? source2Pipe[31:24] : 8'h0) | (compressDataVec_hitReq_4_112 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_112 ? source2Pipe[47:40] : 8'h0)
    | (compressDataVec_hitReq_6_112 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_112 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_112 ? source2Pipe[71:64] : 8'h0)
    | (compressDataVec_hitReq_9_112 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_112 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_112 ? source2Pipe[95:88] : 8'h0)
    | (compressDataVec_hitReq_12_112 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_112 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_112 ? source2Pipe[119:112] : 8'h0)
    | (compressDataVec_hitReq_15_112 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_112 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_112 ? source2Pipe[143:136] : 8'h0)
    | (compressDataVec_hitReq_18_112 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_112 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_112 ? source2Pipe[167:160] : 8'h0)
    | (compressDataVec_hitReq_21_112 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_112 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_112 ? source2Pipe[191:184] : 8'h0)
    | (compressDataVec_hitReq_24_112 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_112 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_112 ? source2Pipe[215:208] : 8'h0)
    | (compressDataVec_hitReq_27_112 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_112 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_112 ? source2Pipe[239:232] : 8'h0)
    | (compressDataVec_hitReq_30_112 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_112 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_112 ? source2Pipe[263:256] : 8'h0)
    | (compressDataVec_hitReq_33_112 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_112 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_112 ? source2Pipe[287:280] : 8'h0)
    | (compressDataVec_hitReq_36_112 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_112 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_112 ? source2Pipe[311:304] : 8'h0)
    | (compressDataVec_hitReq_39_112 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_112 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_112 ? source2Pipe[335:328] : 8'h0)
    | (compressDataVec_hitReq_42_112 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_112 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_112 ? source2Pipe[359:352] : 8'h0)
    | (compressDataVec_hitReq_45_112 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_112 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_112 ? source2Pipe[383:376] : 8'h0)
    | (compressDataVec_hitReq_48_112 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_112 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_112 ? source2Pipe[407:400] : 8'h0)
    | (compressDataVec_hitReq_51_112 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_112 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_112 ? source2Pipe[431:424] : 8'h0)
    | (compressDataVec_hitReq_54_112 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_112 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_112 ? source2Pipe[455:448] : 8'h0)
    | (compressDataVec_hitReq_57_112 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_112 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_112 ? source2Pipe[479:472] : 8'h0)
    | (compressDataVec_hitReq_60_112 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_112 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_112 ? source2Pipe[503:496] : 8'h0)
    | (compressDataVec_hitReq_63_112 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_113 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h71;
  wire          compressDataVec_hitReq_1_113 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h71;
  wire          compressDataVec_hitReq_2_113 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h71;
  wire          compressDataVec_hitReq_3_113 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h71;
  wire          compressDataVec_hitReq_4_113 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h71;
  wire          compressDataVec_hitReq_5_113 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h71;
  wire          compressDataVec_hitReq_6_113 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h71;
  wire          compressDataVec_hitReq_7_113 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h71;
  wire          compressDataVec_hitReq_8_113 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h71;
  wire          compressDataVec_hitReq_9_113 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h71;
  wire          compressDataVec_hitReq_10_113 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h71;
  wire          compressDataVec_hitReq_11_113 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h71;
  wire          compressDataVec_hitReq_12_113 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h71;
  wire          compressDataVec_hitReq_13_113 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h71;
  wire          compressDataVec_hitReq_14_113 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h71;
  wire          compressDataVec_hitReq_15_113 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h71;
  wire          compressDataVec_hitReq_16_113 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h71;
  wire          compressDataVec_hitReq_17_113 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h71;
  wire          compressDataVec_hitReq_18_113 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h71;
  wire          compressDataVec_hitReq_19_113 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h71;
  wire          compressDataVec_hitReq_20_113 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h71;
  wire          compressDataVec_hitReq_21_113 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h71;
  wire          compressDataVec_hitReq_22_113 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h71;
  wire          compressDataVec_hitReq_23_113 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h71;
  wire          compressDataVec_hitReq_24_113 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h71;
  wire          compressDataVec_hitReq_25_113 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h71;
  wire          compressDataVec_hitReq_26_113 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h71;
  wire          compressDataVec_hitReq_27_113 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h71;
  wire          compressDataVec_hitReq_28_113 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h71;
  wire          compressDataVec_hitReq_29_113 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h71;
  wire          compressDataVec_hitReq_30_113 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h71;
  wire          compressDataVec_hitReq_31_113 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h71;
  wire          compressDataVec_hitReq_32_113 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h71;
  wire          compressDataVec_hitReq_33_113 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h71;
  wire          compressDataVec_hitReq_34_113 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h71;
  wire          compressDataVec_hitReq_35_113 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h71;
  wire          compressDataVec_hitReq_36_113 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h71;
  wire          compressDataVec_hitReq_37_113 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h71;
  wire          compressDataVec_hitReq_38_113 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h71;
  wire          compressDataVec_hitReq_39_113 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h71;
  wire          compressDataVec_hitReq_40_113 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h71;
  wire          compressDataVec_hitReq_41_113 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h71;
  wire          compressDataVec_hitReq_42_113 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h71;
  wire          compressDataVec_hitReq_43_113 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h71;
  wire          compressDataVec_hitReq_44_113 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h71;
  wire          compressDataVec_hitReq_45_113 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h71;
  wire          compressDataVec_hitReq_46_113 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h71;
  wire          compressDataVec_hitReq_47_113 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h71;
  wire          compressDataVec_hitReq_48_113 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h71;
  wire          compressDataVec_hitReq_49_113 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h71;
  wire          compressDataVec_hitReq_50_113 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h71;
  wire          compressDataVec_hitReq_51_113 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h71;
  wire          compressDataVec_hitReq_52_113 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h71;
  wire          compressDataVec_hitReq_53_113 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h71;
  wire          compressDataVec_hitReq_54_113 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h71;
  wire          compressDataVec_hitReq_55_113 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h71;
  wire          compressDataVec_hitReq_56_113 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h71;
  wire          compressDataVec_hitReq_57_113 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h71;
  wire          compressDataVec_hitReq_58_113 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h71;
  wire          compressDataVec_hitReq_59_113 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h71;
  wire          compressDataVec_hitReq_60_113 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h71;
  wire          compressDataVec_hitReq_61_113 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h71;
  wire          compressDataVec_hitReq_62_113 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h71;
  wire          compressDataVec_hitReq_63_113 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h71;
  wire [7:0]    compressDataVec_selectReqData_113 =
    (compressDataVec_hitReq_0_113 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_113 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_113 ? source2Pipe[23:16] : 8'h0)
    | (compressDataVec_hitReq_3_113 ? source2Pipe[31:24] : 8'h0) | (compressDataVec_hitReq_4_113 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_113 ? source2Pipe[47:40] : 8'h0)
    | (compressDataVec_hitReq_6_113 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_113 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_113 ? source2Pipe[71:64] : 8'h0)
    | (compressDataVec_hitReq_9_113 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_113 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_113 ? source2Pipe[95:88] : 8'h0)
    | (compressDataVec_hitReq_12_113 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_113 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_113 ? source2Pipe[119:112] : 8'h0)
    | (compressDataVec_hitReq_15_113 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_113 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_113 ? source2Pipe[143:136] : 8'h0)
    | (compressDataVec_hitReq_18_113 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_113 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_113 ? source2Pipe[167:160] : 8'h0)
    | (compressDataVec_hitReq_21_113 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_113 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_113 ? source2Pipe[191:184] : 8'h0)
    | (compressDataVec_hitReq_24_113 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_113 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_113 ? source2Pipe[215:208] : 8'h0)
    | (compressDataVec_hitReq_27_113 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_113 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_113 ? source2Pipe[239:232] : 8'h0)
    | (compressDataVec_hitReq_30_113 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_113 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_113 ? source2Pipe[263:256] : 8'h0)
    | (compressDataVec_hitReq_33_113 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_113 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_113 ? source2Pipe[287:280] : 8'h0)
    | (compressDataVec_hitReq_36_113 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_113 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_113 ? source2Pipe[311:304] : 8'h0)
    | (compressDataVec_hitReq_39_113 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_113 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_113 ? source2Pipe[335:328] : 8'h0)
    | (compressDataVec_hitReq_42_113 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_113 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_113 ? source2Pipe[359:352] : 8'h0)
    | (compressDataVec_hitReq_45_113 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_113 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_113 ? source2Pipe[383:376] : 8'h0)
    | (compressDataVec_hitReq_48_113 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_113 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_113 ? source2Pipe[407:400] : 8'h0)
    | (compressDataVec_hitReq_51_113 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_113 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_113 ? source2Pipe[431:424] : 8'h0)
    | (compressDataVec_hitReq_54_113 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_113 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_113 ? source2Pipe[455:448] : 8'h0)
    | (compressDataVec_hitReq_57_113 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_113 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_113 ? source2Pipe[479:472] : 8'h0)
    | (compressDataVec_hitReq_60_113 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_113 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_113 ? source2Pipe[503:496] : 8'h0)
    | (compressDataVec_hitReq_63_113 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_114 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h72;
  wire          compressDataVec_hitReq_1_114 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h72;
  wire          compressDataVec_hitReq_2_114 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h72;
  wire          compressDataVec_hitReq_3_114 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h72;
  wire          compressDataVec_hitReq_4_114 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h72;
  wire          compressDataVec_hitReq_5_114 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h72;
  wire          compressDataVec_hitReq_6_114 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h72;
  wire          compressDataVec_hitReq_7_114 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h72;
  wire          compressDataVec_hitReq_8_114 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h72;
  wire          compressDataVec_hitReq_9_114 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h72;
  wire          compressDataVec_hitReq_10_114 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h72;
  wire          compressDataVec_hitReq_11_114 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h72;
  wire          compressDataVec_hitReq_12_114 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h72;
  wire          compressDataVec_hitReq_13_114 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h72;
  wire          compressDataVec_hitReq_14_114 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h72;
  wire          compressDataVec_hitReq_15_114 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h72;
  wire          compressDataVec_hitReq_16_114 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h72;
  wire          compressDataVec_hitReq_17_114 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h72;
  wire          compressDataVec_hitReq_18_114 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h72;
  wire          compressDataVec_hitReq_19_114 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h72;
  wire          compressDataVec_hitReq_20_114 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h72;
  wire          compressDataVec_hitReq_21_114 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h72;
  wire          compressDataVec_hitReq_22_114 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h72;
  wire          compressDataVec_hitReq_23_114 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h72;
  wire          compressDataVec_hitReq_24_114 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h72;
  wire          compressDataVec_hitReq_25_114 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h72;
  wire          compressDataVec_hitReq_26_114 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h72;
  wire          compressDataVec_hitReq_27_114 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h72;
  wire          compressDataVec_hitReq_28_114 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h72;
  wire          compressDataVec_hitReq_29_114 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h72;
  wire          compressDataVec_hitReq_30_114 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h72;
  wire          compressDataVec_hitReq_31_114 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h72;
  wire          compressDataVec_hitReq_32_114 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h72;
  wire          compressDataVec_hitReq_33_114 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h72;
  wire          compressDataVec_hitReq_34_114 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h72;
  wire          compressDataVec_hitReq_35_114 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h72;
  wire          compressDataVec_hitReq_36_114 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h72;
  wire          compressDataVec_hitReq_37_114 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h72;
  wire          compressDataVec_hitReq_38_114 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h72;
  wire          compressDataVec_hitReq_39_114 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h72;
  wire          compressDataVec_hitReq_40_114 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h72;
  wire          compressDataVec_hitReq_41_114 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h72;
  wire          compressDataVec_hitReq_42_114 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h72;
  wire          compressDataVec_hitReq_43_114 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h72;
  wire          compressDataVec_hitReq_44_114 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h72;
  wire          compressDataVec_hitReq_45_114 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h72;
  wire          compressDataVec_hitReq_46_114 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h72;
  wire          compressDataVec_hitReq_47_114 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h72;
  wire          compressDataVec_hitReq_48_114 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h72;
  wire          compressDataVec_hitReq_49_114 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h72;
  wire          compressDataVec_hitReq_50_114 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h72;
  wire          compressDataVec_hitReq_51_114 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h72;
  wire          compressDataVec_hitReq_52_114 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h72;
  wire          compressDataVec_hitReq_53_114 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h72;
  wire          compressDataVec_hitReq_54_114 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h72;
  wire          compressDataVec_hitReq_55_114 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h72;
  wire          compressDataVec_hitReq_56_114 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h72;
  wire          compressDataVec_hitReq_57_114 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h72;
  wire          compressDataVec_hitReq_58_114 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h72;
  wire          compressDataVec_hitReq_59_114 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h72;
  wire          compressDataVec_hitReq_60_114 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h72;
  wire          compressDataVec_hitReq_61_114 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h72;
  wire          compressDataVec_hitReq_62_114 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h72;
  wire          compressDataVec_hitReq_63_114 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h72;
  wire [7:0]    compressDataVec_selectReqData_114 =
    (compressDataVec_hitReq_0_114 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_114 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_114 ? source2Pipe[23:16] : 8'h0)
    | (compressDataVec_hitReq_3_114 ? source2Pipe[31:24] : 8'h0) | (compressDataVec_hitReq_4_114 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_114 ? source2Pipe[47:40] : 8'h0)
    | (compressDataVec_hitReq_6_114 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_114 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_114 ? source2Pipe[71:64] : 8'h0)
    | (compressDataVec_hitReq_9_114 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_114 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_114 ? source2Pipe[95:88] : 8'h0)
    | (compressDataVec_hitReq_12_114 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_114 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_114 ? source2Pipe[119:112] : 8'h0)
    | (compressDataVec_hitReq_15_114 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_114 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_114 ? source2Pipe[143:136] : 8'h0)
    | (compressDataVec_hitReq_18_114 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_114 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_114 ? source2Pipe[167:160] : 8'h0)
    | (compressDataVec_hitReq_21_114 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_114 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_114 ? source2Pipe[191:184] : 8'h0)
    | (compressDataVec_hitReq_24_114 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_114 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_114 ? source2Pipe[215:208] : 8'h0)
    | (compressDataVec_hitReq_27_114 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_114 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_114 ? source2Pipe[239:232] : 8'h0)
    | (compressDataVec_hitReq_30_114 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_114 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_114 ? source2Pipe[263:256] : 8'h0)
    | (compressDataVec_hitReq_33_114 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_114 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_114 ? source2Pipe[287:280] : 8'h0)
    | (compressDataVec_hitReq_36_114 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_114 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_114 ? source2Pipe[311:304] : 8'h0)
    | (compressDataVec_hitReq_39_114 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_114 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_114 ? source2Pipe[335:328] : 8'h0)
    | (compressDataVec_hitReq_42_114 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_114 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_114 ? source2Pipe[359:352] : 8'h0)
    | (compressDataVec_hitReq_45_114 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_114 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_114 ? source2Pipe[383:376] : 8'h0)
    | (compressDataVec_hitReq_48_114 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_114 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_114 ? source2Pipe[407:400] : 8'h0)
    | (compressDataVec_hitReq_51_114 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_114 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_114 ? source2Pipe[431:424] : 8'h0)
    | (compressDataVec_hitReq_54_114 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_114 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_114 ? source2Pipe[455:448] : 8'h0)
    | (compressDataVec_hitReq_57_114 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_114 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_114 ? source2Pipe[479:472] : 8'h0)
    | (compressDataVec_hitReq_60_114 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_114 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_114 ? source2Pipe[503:496] : 8'h0)
    | (compressDataVec_hitReq_63_114 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_115 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h73;
  wire          compressDataVec_hitReq_1_115 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h73;
  wire          compressDataVec_hitReq_2_115 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h73;
  wire          compressDataVec_hitReq_3_115 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h73;
  wire          compressDataVec_hitReq_4_115 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h73;
  wire          compressDataVec_hitReq_5_115 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h73;
  wire          compressDataVec_hitReq_6_115 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h73;
  wire          compressDataVec_hitReq_7_115 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h73;
  wire          compressDataVec_hitReq_8_115 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h73;
  wire          compressDataVec_hitReq_9_115 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h73;
  wire          compressDataVec_hitReq_10_115 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h73;
  wire          compressDataVec_hitReq_11_115 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h73;
  wire          compressDataVec_hitReq_12_115 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h73;
  wire          compressDataVec_hitReq_13_115 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h73;
  wire          compressDataVec_hitReq_14_115 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h73;
  wire          compressDataVec_hitReq_15_115 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h73;
  wire          compressDataVec_hitReq_16_115 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h73;
  wire          compressDataVec_hitReq_17_115 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h73;
  wire          compressDataVec_hitReq_18_115 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h73;
  wire          compressDataVec_hitReq_19_115 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h73;
  wire          compressDataVec_hitReq_20_115 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h73;
  wire          compressDataVec_hitReq_21_115 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h73;
  wire          compressDataVec_hitReq_22_115 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h73;
  wire          compressDataVec_hitReq_23_115 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h73;
  wire          compressDataVec_hitReq_24_115 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h73;
  wire          compressDataVec_hitReq_25_115 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h73;
  wire          compressDataVec_hitReq_26_115 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h73;
  wire          compressDataVec_hitReq_27_115 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h73;
  wire          compressDataVec_hitReq_28_115 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h73;
  wire          compressDataVec_hitReq_29_115 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h73;
  wire          compressDataVec_hitReq_30_115 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h73;
  wire          compressDataVec_hitReq_31_115 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h73;
  wire          compressDataVec_hitReq_32_115 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h73;
  wire          compressDataVec_hitReq_33_115 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h73;
  wire          compressDataVec_hitReq_34_115 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h73;
  wire          compressDataVec_hitReq_35_115 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h73;
  wire          compressDataVec_hitReq_36_115 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h73;
  wire          compressDataVec_hitReq_37_115 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h73;
  wire          compressDataVec_hitReq_38_115 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h73;
  wire          compressDataVec_hitReq_39_115 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h73;
  wire          compressDataVec_hitReq_40_115 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h73;
  wire          compressDataVec_hitReq_41_115 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h73;
  wire          compressDataVec_hitReq_42_115 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h73;
  wire          compressDataVec_hitReq_43_115 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h73;
  wire          compressDataVec_hitReq_44_115 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h73;
  wire          compressDataVec_hitReq_45_115 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h73;
  wire          compressDataVec_hitReq_46_115 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h73;
  wire          compressDataVec_hitReq_47_115 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h73;
  wire          compressDataVec_hitReq_48_115 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h73;
  wire          compressDataVec_hitReq_49_115 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h73;
  wire          compressDataVec_hitReq_50_115 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h73;
  wire          compressDataVec_hitReq_51_115 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h73;
  wire          compressDataVec_hitReq_52_115 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h73;
  wire          compressDataVec_hitReq_53_115 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h73;
  wire          compressDataVec_hitReq_54_115 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h73;
  wire          compressDataVec_hitReq_55_115 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h73;
  wire          compressDataVec_hitReq_56_115 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h73;
  wire          compressDataVec_hitReq_57_115 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h73;
  wire          compressDataVec_hitReq_58_115 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h73;
  wire          compressDataVec_hitReq_59_115 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h73;
  wire          compressDataVec_hitReq_60_115 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h73;
  wire          compressDataVec_hitReq_61_115 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h73;
  wire          compressDataVec_hitReq_62_115 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h73;
  wire          compressDataVec_hitReq_63_115 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h73;
  wire [7:0]    compressDataVec_selectReqData_115 =
    (compressDataVec_hitReq_0_115 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_115 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_115 ? source2Pipe[23:16] : 8'h0)
    | (compressDataVec_hitReq_3_115 ? source2Pipe[31:24] : 8'h0) | (compressDataVec_hitReq_4_115 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_115 ? source2Pipe[47:40] : 8'h0)
    | (compressDataVec_hitReq_6_115 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_115 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_115 ? source2Pipe[71:64] : 8'h0)
    | (compressDataVec_hitReq_9_115 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_115 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_115 ? source2Pipe[95:88] : 8'h0)
    | (compressDataVec_hitReq_12_115 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_115 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_115 ? source2Pipe[119:112] : 8'h0)
    | (compressDataVec_hitReq_15_115 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_115 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_115 ? source2Pipe[143:136] : 8'h0)
    | (compressDataVec_hitReq_18_115 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_115 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_115 ? source2Pipe[167:160] : 8'h0)
    | (compressDataVec_hitReq_21_115 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_115 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_115 ? source2Pipe[191:184] : 8'h0)
    | (compressDataVec_hitReq_24_115 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_115 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_115 ? source2Pipe[215:208] : 8'h0)
    | (compressDataVec_hitReq_27_115 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_115 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_115 ? source2Pipe[239:232] : 8'h0)
    | (compressDataVec_hitReq_30_115 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_115 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_115 ? source2Pipe[263:256] : 8'h0)
    | (compressDataVec_hitReq_33_115 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_115 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_115 ? source2Pipe[287:280] : 8'h0)
    | (compressDataVec_hitReq_36_115 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_115 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_115 ? source2Pipe[311:304] : 8'h0)
    | (compressDataVec_hitReq_39_115 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_115 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_115 ? source2Pipe[335:328] : 8'h0)
    | (compressDataVec_hitReq_42_115 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_115 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_115 ? source2Pipe[359:352] : 8'h0)
    | (compressDataVec_hitReq_45_115 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_115 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_115 ? source2Pipe[383:376] : 8'h0)
    | (compressDataVec_hitReq_48_115 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_115 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_115 ? source2Pipe[407:400] : 8'h0)
    | (compressDataVec_hitReq_51_115 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_115 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_115 ? source2Pipe[431:424] : 8'h0)
    | (compressDataVec_hitReq_54_115 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_115 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_115 ? source2Pipe[455:448] : 8'h0)
    | (compressDataVec_hitReq_57_115 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_115 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_115 ? source2Pipe[479:472] : 8'h0)
    | (compressDataVec_hitReq_60_115 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_115 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_115 ? source2Pipe[503:496] : 8'h0)
    | (compressDataVec_hitReq_63_115 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_116 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h74;
  wire          compressDataVec_hitReq_1_116 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h74;
  wire          compressDataVec_hitReq_2_116 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h74;
  wire          compressDataVec_hitReq_3_116 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h74;
  wire          compressDataVec_hitReq_4_116 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h74;
  wire          compressDataVec_hitReq_5_116 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h74;
  wire          compressDataVec_hitReq_6_116 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h74;
  wire          compressDataVec_hitReq_7_116 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h74;
  wire          compressDataVec_hitReq_8_116 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h74;
  wire          compressDataVec_hitReq_9_116 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h74;
  wire          compressDataVec_hitReq_10_116 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h74;
  wire          compressDataVec_hitReq_11_116 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h74;
  wire          compressDataVec_hitReq_12_116 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h74;
  wire          compressDataVec_hitReq_13_116 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h74;
  wire          compressDataVec_hitReq_14_116 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h74;
  wire          compressDataVec_hitReq_15_116 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h74;
  wire          compressDataVec_hitReq_16_116 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h74;
  wire          compressDataVec_hitReq_17_116 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h74;
  wire          compressDataVec_hitReq_18_116 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h74;
  wire          compressDataVec_hitReq_19_116 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h74;
  wire          compressDataVec_hitReq_20_116 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h74;
  wire          compressDataVec_hitReq_21_116 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h74;
  wire          compressDataVec_hitReq_22_116 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h74;
  wire          compressDataVec_hitReq_23_116 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h74;
  wire          compressDataVec_hitReq_24_116 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h74;
  wire          compressDataVec_hitReq_25_116 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h74;
  wire          compressDataVec_hitReq_26_116 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h74;
  wire          compressDataVec_hitReq_27_116 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h74;
  wire          compressDataVec_hitReq_28_116 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h74;
  wire          compressDataVec_hitReq_29_116 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h74;
  wire          compressDataVec_hitReq_30_116 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h74;
  wire          compressDataVec_hitReq_31_116 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h74;
  wire          compressDataVec_hitReq_32_116 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h74;
  wire          compressDataVec_hitReq_33_116 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h74;
  wire          compressDataVec_hitReq_34_116 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h74;
  wire          compressDataVec_hitReq_35_116 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h74;
  wire          compressDataVec_hitReq_36_116 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h74;
  wire          compressDataVec_hitReq_37_116 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h74;
  wire          compressDataVec_hitReq_38_116 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h74;
  wire          compressDataVec_hitReq_39_116 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h74;
  wire          compressDataVec_hitReq_40_116 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h74;
  wire          compressDataVec_hitReq_41_116 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h74;
  wire          compressDataVec_hitReq_42_116 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h74;
  wire          compressDataVec_hitReq_43_116 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h74;
  wire          compressDataVec_hitReq_44_116 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h74;
  wire          compressDataVec_hitReq_45_116 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h74;
  wire          compressDataVec_hitReq_46_116 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h74;
  wire          compressDataVec_hitReq_47_116 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h74;
  wire          compressDataVec_hitReq_48_116 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h74;
  wire          compressDataVec_hitReq_49_116 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h74;
  wire          compressDataVec_hitReq_50_116 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h74;
  wire          compressDataVec_hitReq_51_116 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h74;
  wire          compressDataVec_hitReq_52_116 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h74;
  wire          compressDataVec_hitReq_53_116 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h74;
  wire          compressDataVec_hitReq_54_116 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h74;
  wire          compressDataVec_hitReq_55_116 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h74;
  wire          compressDataVec_hitReq_56_116 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h74;
  wire          compressDataVec_hitReq_57_116 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h74;
  wire          compressDataVec_hitReq_58_116 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h74;
  wire          compressDataVec_hitReq_59_116 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h74;
  wire          compressDataVec_hitReq_60_116 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h74;
  wire          compressDataVec_hitReq_61_116 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h74;
  wire          compressDataVec_hitReq_62_116 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h74;
  wire          compressDataVec_hitReq_63_116 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h74;
  wire [7:0]    compressDataVec_selectReqData_116 =
    (compressDataVec_hitReq_0_116 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_116 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_116 ? source2Pipe[23:16] : 8'h0)
    | (compressDataVec_hitReq_3_116 ? source2Pipe[31:24] : 8'h0) | (compressDataVec_hitReq_4_116 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_116 ? source2Pipe[47:40] : 8'h0)
    | (compressDataVec_hitReq_6_116 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_116 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_116 ? source2Pipe[71:64] : 8'h0)
    | (compressDataVec_hitReq_9_116 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_116 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_116 ? source2Pipe[95:88] : 8'h0)
    | (compressDataVec_hitReq_12_116 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_116 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_116 ? source2Pipe[119:112] : 8'h0)
    | (compressDataVec_hitReq_15_116 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_116 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_116 ? source2Pipe[143:136] : 8'h0)
    | (compressDataVec_hitReq_18_116 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_116 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_116 ? source2Pipe[167:160] : 8'h0)
    | (compressDataVec_hitReq_21_116 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_116 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_116 ? source2Pipe[191:184] : 8'h0)
    | (compressDataVec_hitReq_24_116 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_116 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_116 ? source2Pipe[215:208] : 8'h0)
    | (compressDataVec_hitReq_27_116 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_116 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_116 ? source2Pipe[239:232] : 8'h0)
    | (compressDataVec_hitReq_30_116 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_116 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_116 ? source2Pipe[263:256] : 8'h0)
    | (compressDataVec_hitReq_33_116 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_116 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_116 ? source2Pipe[287:280] : 8'h0)
    | (compressDataVec_hitReq_36_116 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_116 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_116 ? source2Pipe[311:304] : 8'h0)
    | (compressDataVec_hitReq_39_116 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_116 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_116 ? source2Pipe[335:328] : 8'h0)
    | (compressDataVec_hitReq_42_116 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_116 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_116 ? source2Pipe[359:352] : 8'h0)
    | (compressDataVec_hitReq_45_116 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_116 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_116 ? source2Pipe[383:376] : 8'h0)
    | (compressDataVec_hitReq_48_116 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_116 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_116 ? source2Pipe[407:400] : 8'h0)
    | (compressDataVec_hitReq_51_116 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_116 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_116 ? source2Pipe[431:424] : 8'h0)
    | (compressDataVec_hitReq_54_116 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_116 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_116 ? source2Pipe[455:448] : 8'h0)
    | (compressDataVec_hitReq_57_116 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_116 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_116 ? source2Pipe[479:472] : 8'h0)
    | (compressDataVec_hitReq_60_116 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_116 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_116 ? source2Pipe[503:496] : 8'h0)
    | (compressDataVec_hitReq_63_116 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_117 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h75;
  wire          compressDataVec_hitReq_1_117 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h75;
  wire          compressDataVec_hitReq_2_117 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h75;
  wire          compressDataVec_hitReq_3_117 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h75;
  wire          compressDataVec_hitReq_4_117 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h75;
  wire          compressDataVec_hitReq_5_117 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h75;
  wire          compressDataVec_hitReq_6_117 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h75;
  wire          compressDataVec_hitReq_7_117 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h75;
  wire          compressDataVec_hitReq_8_117 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h75;
  wire          compressDataVec_hitReq_9_117 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h75;
  wire          compressDataVec_hitReq_10_117 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h75;
  wire          compressDataVec_hitReq_11_117 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h75;
  wire          compressDataVec_hitReq_12_117 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h75;
  wire          compressDataVec_hitReq_13_117 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h75;
  wire          compressDataVec_hitReq_14_117 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h75;
  wire          compressDataVec_hitReq_15_117 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h75;
  wire          compressDataVec_hitReq_16_117 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h75;
  wire          compressDataVec_hitReq_17_117 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h75;
  wire          compressDataVec_hitReq_18_117 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h75;
  wire          compressDataVec_hitReq_19_117 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h75;
  wire          compressDataVec_hitReq_20_117 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h75;
  wire          compressDataVec_hitReq_21_117 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h75;
  wire          compressDataVec_hitReq_22_117 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h75;
  wire          compressDataVec_hitReq_23_117 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h75;
  wire          compressDataVec_hitReq_24_117 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h75;
  wire          compressDataVec_hitReq_25_117 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h75;
  wire          compressDataVec_hitReq_26_117 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h75;
  wire          compressDataVec_hitReq_27_117 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h75;
  wire          compressDataVec_hitReq_28_117 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h75;
  wire          compressDataVec_hitReq_29_117 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h75;
  wire          compressDataVec_hitReq_30_117 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h75;
  wire          compressDataVec_hitReq_31_117 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h75;
  wire          compressDataVec_hitReq_32_117 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h75;
  wire          compressDataVec_hitReq_33_117 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h75;
  wire          compressDataVec_hitReq_34_117 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h75;
  wire          compressDataVec_hitReq_35_117 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h75;
  wire          compressDataVec_hitReq_36_117 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h75;
  wire          compressDataVec_hitReq_37_117 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h75;
  wire          compressDataVec_hitReq_38_117 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h75;
  wire          compressDataVec_hitReq_39_117 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h75;
  wire          compressDataVec_hitReq_40_117 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h75;
  wire          compressDataVec_hitReq_41_117 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h75;
  wire          compressDataVec_hitReq_42_117 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h75;
  wire          compressDataVec_hitReq_43_117 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h75;
  wire          compressDataVec_hitReq_44_117 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h75;
  wire          compressDataVec_hitReq_45_117 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h75;
  wire          compressDataVec_hitReq_46_117 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h75;
  wire          compressDataVec_hitReq_47_117 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h75;
  wire          compressDataVec_hitReq_48_117 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h75;
  wire          compressDataVec_hitReq_49_117 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h75;
  wire          compressDataVec_hitReq_50_117 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h75;
  wire          compressDataVec_hitReq_51_117 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h75;
  wire          compressDataVec_hitReq_52_117 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h75;
  wire          compressDataVec_hitReq_53_117 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h75;
  wire          compressDataVec_hitReq_54_117 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h75;
  wire          compressDataVec_hitReq_55_117 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h75;
  wire          compressDataVec_hitReq_56_117 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h75;
  wire          compressDataVec_hitReq_57_117 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h75;
  wire          compressDataVec_hitReq_58_117 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h75;
  wire          compressDataVec_hitReq_59_117 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h75;
  wire          compressDataVec_hitReq_60_117 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h75;
  wire          compressDataVec_hitReq_61_117 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h75;
  wire          compressDataVec_hitReq_62_117 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h75;
  wire          compressDataVec_hitReq_63_117 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h75;
  wire [7:0]    compressDataVec_selectReqData_117 =
    (compressDataVec_hitReq_0_117 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_117 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_117 ? source2Pipe[23:16] : 8'h0)
    | (compressDataVec_hitReq_3_117 ? source2Pipe[31:24] : 8'h0) | (compressDataVec_hitReq_4_117 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_117 ? source2Pipe[47:40] : 8'h0)
    | (compressDataVec_hitReq_6_117 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_117 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_117 ? source2Pipe[71:64] : 8'h0)
    | (compressDataVec_hitReq_9_117 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_117 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_117 ? source2Pipe[95:88] : 8'h0)
    | (compressDataVec_hitReq_12_117 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_117 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_117 ? source2Pipe[119:112] : 8'h0)
    | (compressDataVec_hitReq_15_117 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_117 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_117 ? source2Pipe[143:136] : 8'h0)
    | (compressDataVec_hitReq_18_117 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_117 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_117 ? source2Pipe[167:160] : 8'h0)
    | (compressDataVec_hitReq_21_117 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_117 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_117 ? source2Pipe[191:184] : 8'h0)
    | (compressDataVec_hitReq_24_117 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_117 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_117 ? source2Pipe[215:208] : 8'h0)
    | (compressDataVec_hitReq_27_117 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_117 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_117 ? source2Pipe[239:232] : 8'h0)
    | (compressDataVec_hitReq_30_117 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_117 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_117 ? source2Pipe[263:256] : 8'h0)
    | (compressDataVec_hitReq_33_117 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_117 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_117 ? source2Pipe[287:280] : 8'h0)
    | (compressDataVec_hitReq_36_117 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_117 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_117 ? source2Pipe[311:304] : 8'h0)
    | (compressDataVec_hitReq_39_117 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_117 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_117 ? source2Pipe[335:328] : 8'h0)
    | (compressDataVec_hitReq_42_117 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_117 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_117 ? source2Pipe[359:352] : 8'h0)
    | (compressDataVec_hitReq_45_117 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_117 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_117 ? source2Pipe[383:376] : 8'h0)
    | (compressDataVec_hitReq_48_117 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_117 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_117 ? source2Pipe[407:400] : 8'h0)
    | (compressDataVec_hitReq_51_117 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_117 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_117 ? source2Pipe[431:424] : 8'h0)
    | (compressDataVec_hitReq_54_117 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_117 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_117 ? source2Pipe[455:448] : 8'h0)
    | (compressDataVec_hitReq_57_117 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_117 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_117 ? source2Pipe[479:472] : 8'h0)
    | (compressDataVec_hitReq_60_117 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_117 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_117 ? source2Pipe[503:496] : 8'h0)
    | (compressDataVec_hitReq_63_117 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_118 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h76;
  wire          compressDataVec_hitReq_1_118 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h76;
  wire          compressDataVec_hitReq_2_118 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h76;
  wire          compressDataVec_hitReq_3_118 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h76;
  wire          compressDataVec_hitReq_4_118 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h76;
  wire          compressDataVec_hitReq_5_118 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h76;
  wire          compressDataVec_hitReq_6_118 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h76;
  wire          compressDataVec_hitReq_7_118 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h76;
  wire          compressDataVec_hitReq_8_118 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h76;
  wire          compressDataVec_hitReq_9_118 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h76;
  wire          compressDataVec_hitReq_10_118 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h76;
  wire          compressDataVec_hitReq_11_118 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h76;
  wire          compressDataVec_hitReq_12_118 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h76;
  wire          compressDataVec_hitReq_13_118 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h76;
  wire          compressDataVec_hitReq_14_118 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h76;
  wire          compressDataVec_hitReq_15_118 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h76;
  wire          compressDataVec_hitReq_16_118 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h76;
  wire          compressDataVec_hitReq_17_118 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h76;
  wire          compressDataVec_hitReq_18_118 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h76;
  wire          compressDataVec_hitReq_19_118 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h76;
  wire          compressDataVec_hitReq_20_118 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h76;
  wire          compressDataVec_hitReq_21_118 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h76;
  wire          compressDataVec_hitReq_22_118 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h76;
  wire          compressDataVec_hitReq_23_118 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h76;
  wire          compressDataVec_hitReq_24_118 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h76;
  wire          compressDataVec_hitReq_25_118 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h76;
  wire          compressDataVec_hitReq_26_118 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h76;
  wire          compressDataVec_hitReq_27_118 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h76;
  wire          compressDataVec_hitReq_28_118 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h76;
  wire          compressDataVec_hitReq_29_118 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h76;
  wire          compressDataVec_hitReq_30_118 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h76;
  wire          compressDataVec_hitReq_31_118 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h76;
  wire          compressDataVec_hitReq_32_118 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h76;
  wire          compressDataVec_hitReq_33_118 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h76;
  wire          compressDataVec_hitReq_34_118 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h76;
  wire          compressDataVec_hitReq_35_118 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h76;
  wire          compressDataVec_hitReq_36_118 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h76;
  wire          compressDataVec_hitReq_37_118 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h76;
  wire          compressDataVec_hitReq_38_118 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h76;
  wire          compressDataVec_hitReq_39_118 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h76;
  wire          compressDataVec_hitReq_40_118 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h76;
  wire          compressDataVec_hitReq_41_118 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h76;
  wire          compressDataVec_hitReq_42_118 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h76;
  wire          compressDataVec_hitReq_43_118 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h76;
  wire          compressDataVec_hitReq_44_118 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h76;
  wire          compressDataVec_hitReq_45_118 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h76;
  wire          compressDataVec_hitReq_46_118 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h76;
  wire          compressDataVec_hitReq_47_118 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h76;
  wire          compressDataVec_hitReq_48_118 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h76;
  wire          compressDataVec_hitReq_49_118 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h76;
  wire          compressDataVec_hitReq_50_118 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h76;
  wire          compressDataVec_hitReq_51_118 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h76;
  wire          compressDataVec_hitReq_52_118 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h76;
  wire          compressDataVec_hitReq_53_118 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h76;
  wire          compressDataVec_hitReq_54_118 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h76;
  wire          compressDataVec_hitReq_55_118 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h76;
  wire          compressDataVec_hitReq_56_118 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h76;
  wire          compressDataVec_hitReq_57_118 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h76;
  wire          compressDataVec_hitReq_58_118 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h76;
  wire          compressDataVec_hitReq_59_118 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h76;
  wire          compressDataVec_hitReq_60_118 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h76;
  wire          compressDataVec_hitReq_61_118 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h76;
  wire          compressDataVec_hitReq_62_118 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h76;
  wire          compressDataVec_hitReq_63_118 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h76;
  wire [7:0]    compressDataVec_selectReqData_118 =
    (compressDataVec_hitReq_0_118 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_118 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_118 ? source2Pipe[23:16] : 8'h0)
    | (compressDataVec_hitReq_3_118 ? source2Pipe[31:24] : 8'h0) | (compressDataVec_hitReq_4_118 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_118 ? source2Pipe[47:40] : 8'h0)
    | (compressDataVec_hitReq_6_118 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_118 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_118 ? source2Pipe[71:64] : 8'h0)
    | (compressDataVec_hitReq_9_118 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_118 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_118 ? source2Pipe[95:88] : 8'h0)
    | (compressDataVec_hitReq_12_118 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_118 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_118 ? source2Pipe[119:112] : 8'h0)
    | (compressDataVec_hitReq_15_118 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_118 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_118 ? source2Pipe[143:136] : 8'h0)
    | (compressDataVec_hitReq_18_118 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_118 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_118 ? source2Pipe[167:160] : 8'h0)
    | (compressDataVec_hitReq_21_118 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_118 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_118 ? source2Pipe[191:184] : 8'h0)
    | (compressDataVec_hitReq_24_118 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_118 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_118 ? source2Pipe[215:208] : 8'h0)
    | (compressDataVec_hitReq_27_118 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_118 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_118 ? source2Pipe[239:232] : 8'h0)
    | (compressDataVec_hitReq_30_118 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_118 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_118 ? source2Pipe[263:256] : 8'h0)
    | (compressDataVec_hitReq_33_118 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_118 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_118 ? source2Pipe[287:280] : 8'h0)
    | (compressDataVec_hitReq_36_118 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_118 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_118 ? source2Pipe[311:304] : 8'h0)
    | (compressDataVec_hitReq_39_118 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_118 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_118 ? source2Pipe[335:328] : 8'h0)
    | (compressDataVec_hitReq_42_118 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_118 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_118 ? source2Pipe[359:352] : 8'h0)
    | (compressDataVec_hitReq_45_118 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_118 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_118 ? source2Pipe[383:376] : 8'h0)
    | (compressDataVec_hitReq_48_118 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_118 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_118 ? source2Pipe[407:400] : 8'h0)
    | (compressDataVec_hitReq_51_118 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_118 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_118 ? source2Pipe[431:424] : 8'h0)
    | (compressDataVec_hitReq_54_118 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_118 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_118 ? source2Pipe[455:448] : 8'h0)
    | (compressDataVec_hitReq_57_118 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_118 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_118 ? source2Pipe[479:472] : 8'h0)
    | (compressDataVec_hitReq_60_118 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_118 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_118 ? source2Pipe[503:496] : 8'h0)
    | (compressDataVec_hitReq_63_118 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_119 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h77;
  wire          compressDataVec_hitReq_1_119 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h77;
  wire          compressDataVec_hitReq_2_119 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h77;
  wire          compressDataVec_hitReq_3_119 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h77;
  wire          compressDataVec_hitReq_4_119 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h77;
  wire          compressDataVec_hitReq_5_119 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h77;
  wire          compressDataVec_hitReq_6_119 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h77;
  wire          compressDataVec_hitReq_7_119 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h77;
  wire          compressDataVec_hitReq_8_119 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h77;
  wire          compressDataVec_hitReq_9_119 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h77;
  wire          compressDataVec_hitReq_10_119 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h77;
  wire          compressDataVec_hitReq_11_119 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h77;
  wire          compressDataVec_hitReq_12_119 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h77;
  wire          compressDataVec_hitReq_13_119 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h77;
  wire          compressDataVec_hitReq_14_119 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h77;
  wire          compressDataVec_hitReq_15_119 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h77;
  wire          compressDataVec_hitReq_16_119 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h77;
  wire          compressDataVec_hitReq_17_119 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h77;
  wire          compressDataVec_hitReq_18_119 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h77;
  wire          compressDataVec_hitReq_19_119 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h77;
  wire          compressDataVec_hitReq_20_119 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h77;
  wire          compressDataVec_hitReq_21_119 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h77;
  wire          compressDataVec_hitReq_22_119 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h77;
  wire          compressDataVec_hitReq_23_119 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h77;
  wire          compressDataVec_hitReq_24_119 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h77;
  wire          compressDataVec_hitReq_25_119 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h77;
  wire          compressDataVec_hitReq_26_119 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h77;
  wire          compressDataVec_hitReq_27_119 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h77;
  wire          compressDataVec_hitReq_28_119 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h77;
  wire          compressDataVec_hitReq_29_119 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h77;
  wire          compressDataVec_hitReq_30_119 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h77;
  wire          compressDataVec_hitReq_31_119 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h77;
  wire          compressDataVec_hitReq_32_119 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h77;
  wire          compressDataVec_hitReq_33_119 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h77;
  wire          compressDataVec_hitReq_34_119 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h77;
  wire          compressDataVec_hitReq_35_119 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h77;
  wire          compressDataVec_hitReq_36_119 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h77;
  wire          compressDataVec_hitReq_37_119 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h77;
  wire          compressDataVec_hitReq_38_119 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h77;
  wire          compressDataVec_hitReq_39_119 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h77;
  wire          compressDataVec_hitReq_40_119 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h77;
  wire          compressDataVec_hitReq_41_119 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h77;
  wire          compressDataVec_hitReq_42_119 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h77;
  wire          compressDataVec_hitReq_43_119 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h77;
  wire          compressDataVec_hitReq_44_119 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h77;
  wire          compressDataVec_hitReq_45_119 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h77;
  wire          compressDataVec_hitReq_46_119 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h77;
  wire          compressDataVec_hitReq_47_119 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h77;
  wire          compressDataVec_hitReq_48_119 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h77;
  wire          compressDataVec_hitReq_49_119 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h77;
  wire          compressDataVec_hitReq_50_119 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h77;
  wire          compressDataVec_hitReq_51_119 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h77;
  wire          compressDataVec_hitReq_52_119 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h77;
  wire          compressDataVec_hitReq_53_119 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h77;
  wire          compressDataVec_hitReq_54_119 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h77;
  wire          compressDataVec_hitReq_55_119 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h77;
  wire          compressDataVec_hitReq_56_119 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h77;
  wire          compressDataVec_hitReq_57_119 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h77;
  wire          compressDataVec_hitReq_58_119 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h77;
  wire          compressDataVec_hitReq_59_119 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h77;
  wire          compressDataVec_hitReq_60_119 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h77;
  wire          compressDataVec_hitReq_61_119 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h77;
  wire          compressDataVec_hitReq_62_119 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h77;
  wire          compressDataVec_hitReq_63_119 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h77;
  wire [7:0]    compressDataVec_selectReqData_119 =
    (compressDataVec_hitReq_0_119 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_119 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_119 ? source2Pipe[23:16] : 8'h0)
    | (compressDataVec_hitReq_3_119 ? source2Pipe[31:24] : 8'h0) | (compressDataVec_hitReq_4_119 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_119 ? source2Pipe[47:40] : 8'h0)
    | (compressDataVec_hitReq_6_119 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_119 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_119 ? source2Pipe[71:64] : 8'h0)
    | (compressDataVec_hitReq_9_119 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_119 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_119 ? source2Pipe[95:88] : 8'h0)
    | (compressDataVec_hitReq_12_119 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_119 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_119 ? source2Pipe[119:112] : 8'h0)
    | (compressDataVec_hitReq_15_119 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_119 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_119 ? source2Pipe[143:136] : 8'h0)
    | (compressDataVec_hitReq_18_119 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_119 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_119 ? source2Pipe[167:160] : 8'h0)
    | (compressDataVec_hitReq_21_119 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_119 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_119 ? source2Pipe[191:184] : 8'h0)
    | (compressDataVec_hitReq_24_119 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_119 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_119 ? source2Pipe[215:208] : 8'h0)
    | (compressDataVec_hitReq_27_119 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_119 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_119 ? source2Pipe[239:232] : 8'h0)
    | (compressDataVec_hitReq_30_119 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_119 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_119 ? source2Pipe[263:256] : 8'h0)
    | (compressDataVec_hitReq_33_119 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_119 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_119 ? source2Pipe[287:280] : 8'h0)
    | (compressDataVec_hitReq_36_119 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_119 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_119 ? source2Pipe[311:304] : 8'h0)
    | (compressDataVec_hitReq_39_119 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_119 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_119 ? source2Pipe[335:328] : 8'h0)
    | (compressDataVec_hitReq_42_119 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_119 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_119 ? source2Pipe[359:352] : 8'h0)
    | (compressDataVec_hitReq_45_119 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_119 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_119 ? source2Pipe[383:376] : 8'h0)
    | (compressDataVec_hitReq_48_119 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_119 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_119 ? source2Pipe[407:400] : 8'h0)
    | (compressDataVec_hitReq_51_119 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_119 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_119 ? source2Pipe[431:424] : 8'h0)
    | (compressDataVec_hitReq_54_119 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_119 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_119 ? source2Pipe[455:448] : 8'h0)
    | (compressDataVec_hitReq_57_119 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_119 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_119 ? source2Pipe[479:472] : 8'h0)
    | (compressDataVec_hitReq_60_119 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_119 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_119 ? source2Pipe[503:496] : 8'h0)
    | (compressDataVec_hitReq_63_119 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_120 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h78;
  wire          compressDataVec_hitReq_1_120 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h78;
  wire          compressDataVec_hitReq_2_120 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h78;
  wire          compressDataVec_hitReq_3_120 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h78;
  wire          compressDataVec_hitReq_4_120 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h78;
  wire          compressDataVec_hitReq_5_120 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h78;
  wire          compressDataVec_hitReq_6_120 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h78;
  wire          compressDataVec_hitReq_7_120 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h78;
  wire          compressDataVec_hitReq_8_120 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h78;
  wire          compressDataVec_hitReq_9_120 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h78;
  wire          compressDataVec_hitReq_10_120 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h78;
  wire          compressDataVec_hitReq_11_120 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h78;
  wire          compressDataVec_hitReq_12_120 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h78;
  wire          compressDataVec_hitReq_13_120 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h78;
  wire          compressDataVec_hitReq_14_120 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h78;
  wire          compressDataVec_hitReq_15_120 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h78;
  wire          compressDataVec_hitReq_16_120 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h78;
  wire          compressDataVec_hitReq_17_120 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h78;
  wire          compressDataVec_hitReq_18_120 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h78;
  wire          compressDataVec_hitReq_19_120 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h78;
  wire          compressDataVec_hitReq_20_120 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h78;
  wire          compressDataVec_hitReq_21_120 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h78;
  wire          compressDataVec_hitReq_22_120 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h78;
  wire          compressDataVec_hitReq_23_120 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h78;
  wire          compressDataVec_hitReq_24_120 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h78;
  wire          compressDataVec_hitReq_25_120 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h78;
  wire          compressDataVec_hitReq_26_120 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h78;
  wire          compressDataVec_hitReq_27_120 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h78;
  wire          compressDataVec_hitReq_28_120 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h78;
  wire          compressDataVec_hitReq_29_120 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h78;
  wire          compressDataVec_hitReq_30_120 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h78;
  wire          compressDataVec_hitReq_31_120 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h78;
  wire          compressDataVec_hitReq_32_120 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h78;
  wire          compressDataVec_hitReq_33_120 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h78;
  wire          compressDataVec_hitReq_34_120 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h78;
  wire          compressDataVec_hitReq_35_120 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h78;
  wire          compressDataVec_hitReq_36_120 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h78;
  wire          compressDataVec_hitReq_37_120 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h78;
  wire          compressDataVec_hitReq_38_120 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h78;
  wire          compressDataVec_hitReq_39_120 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h78;
  wire          compressDataVec_hitReq_40_120 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h78;
  wire          compressDataVec_hitReq_41_120 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h78;
  wire          compressDataVec_hitReq_42_120 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h78;
  wire          compressDataVec_hitReq_43_120 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h78;
  wire          compressDataVec_hitReq_44_120 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h78;
  wire          compressDataVec_hitReq_45_120 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h78;
  wire          compressDataVec_hitReq_46_120 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h78;
  wire          compressDataVec_hitReq_47_120 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h78;
  wire          compressDataVec_hitReq_48_120 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h78;
  wire          compressDataVec_hitReq_49_120 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h78;
  wire          compressDataVec_hitReq_50_120 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h78;
  wire          compressDataVec_hitReq_51_120 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h78;
  wire          compressDataVec_hitReq_52_120 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h78;
  wire          compressDataVec_hitReq_53_120 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h78;
  wire          compressDataVec_hitReq_54_120 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h78;
  wire          compressDataVec_hitReq_55_120 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h78;
  wire          compressDataVec_hitReq_56_120 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h78;
  wire          compressDataVec_hitReq_57_120 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h78;
  wire          compressDataVec_hitReq_58_120 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h78;
  wire          compressDataVec_hitReq_59_120 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h78;
  wire          compressDataVec_hitReq_60_120 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h78;
  wire          compressDataVec_hitReq_61_120 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h78;
  wire          compressDataVec_hitReq_62_120 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h78;
  wire          compressDataVec_hitReq_63_120 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h78;
  wire [7:0]    compressDataVec_selectReqData_120 =
    (compressDataVec_hitReq_0_120 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_120 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_120 ? source2Pipe[23:16] : 8'h0)
    | (compressDataVec_hitReq_3_120 ? source2Pipe[31:24] : 8'h0) | (compressDataVec_hitReq_4_120 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_120 ? source2Pipe[47:40] : 8'h0)
    | (compressDataVec_hitReq_6_120 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_120 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_120 ? source2Pipe[71:64] : 8'h0)
    | (compressDataVec_hitReq_9_120 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_120 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_120 ? source2Pipe[95:88] : 8'h0)
    | (compressDataVec_hitReq_12_120 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_120 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_120 ? source2Pipe[119:112] : 8'h0)
    | (compressDataVec_hitReq_15_120 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_120 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_120 ? source2Pipe[143:136] : 8'h0)
    | (compressDataVec_hitReq_18_120 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_120 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_120 ? source2Pipe[167:160] : 8'h0)
    | (compressDataVec_hitReq_21_120 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_120 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_120 ? source2Pipe[191:184] : 8'h0)
    | (compressDataVec_hitReq_24_120 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_120 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_120 ? source2Pipe[215:208] : 8'h0)
    | (compressDataVec_hitReq_27_120 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_120 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_120 ? source2Pipe[239:232] : 8'h0)
    | (compressDataVec_hitReq_30_120 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_120 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_120 ? source2Pipe[263:256] : 8'h0)
    | (compressDataVec_hitReq_33_120 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_120 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_120 ? source2Pipe[287:280] : 8'h0)
    | (compressDataVec_hitReq_36_120 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_120 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_120 ? source2Pipe[311:304] : 8'h0)
    | (compressDataVec_hitReq_39_120 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_120 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_120 ? source2Pipe[335:328] : 8'h0)
    | (compressDataVec_hitReq_42_120 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_120 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_120 ? source2Pipe[359:352] : 8'h0)
    | (compressDataVec_hitReq_45_120 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_120 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_120 ? source2Pipe[383:376] : 8'h0)
    | (compressDataVec_hitReq_48_120 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_120 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_120 ? source2Pipe[407:400] : 8'h0)
    | (compressDataVec_hitReq_51_120 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_120 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_120 ? source2Pipe[431:424] : 8'h0)
    | (compressDataVec_hitReq_54_120 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_120 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_120 ? source2Pipe[455:448] : 8'h0)
    | (compressDataVec_hitReq_57_120 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_120 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_120 ? source2Pipe[479:472] : 8'h0)
    | (compressDataVec_hitReq_60_120 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_120 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_120 ? source2Pipe[503:496] : 8'h0)
    | (compressDataVec_hitReq_63_120 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_121 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h79;
  wire          compressDataVec_hitReq_1_121 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h79;
  wire          compressDataVec_hitReq_2_121 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h79;
  wire          compressDataVec_hitReq_3_121 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h79;
  wire          compressDataVec_hitReq_4_121 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h79;
  wire          compressDataVec_hitReq_5_121 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h79;
  wire          compressDataVec_hitReq_6_121 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h79;
  wire          compressDataVec_hitReq_7_121 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h79;
  wire          compressDataVec_hitReq_8_121 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h79;
  wire          compressDataVec_hitReq_9_121 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h79;
  wire          compressDataVec_hitReq_10_121 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h79;
  wire          compressDataVec_hitReq_11_121 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h79;
  wire          compressDataVec_hitReq_12_121 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h79;
  wire          compressDataVec_hitReq_13_121 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h79;
  wire          compressDataVec_hitReq_14_121 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h79;
  wire          compressDataVec_hitReq_15_121 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h79;
  wire          compressDataVec_hitReq_16_121 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h79;
  wire          compressDataVec_hitReq_17_121 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h79;
  wire          compressDataVec_hitReq_18_121 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h79;
  wire          compressDataVec_hitReq_19_121 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h79;
  wire          compressDataVec_hitReq_20_121 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h79;
  wire          compressDataVec_hitReq_21_121 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h79;
  wire          compressDataVec_hitReq_22_121 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h79;
  wire          compressDataVec_hitReq_23_121 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h79;
  wire          compressDataVec_hitReq_24_121 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h79;
  wire          compressDataVec_hitReq_25_121 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h79;
  wire          compressDataVec_hitReq_26_121 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h79;
  wire          compressDataVec_hitReq_27_121 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h79;
  wire          compressDataVec_hitReq_28_121 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h79;
  wire          compressDataVec_hitReq_29_121 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h79;
  wire          compressDataVec_hitReq_30_121 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h79;
  wire          compressDataVec_hitReq_31_121 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h79;
  wire          compressDataVec_hitReq_32_121 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h79;
  wire          compressDataVec_hitReq_33_121 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h79;
  wire          compressDataVec_hitReq_34_121 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h79;
  wire          compressDataVec_hitReq_35_121 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h79;
  wire          compressDataVec_hitReq_36_121 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h79;
  wire          compressDataVec_hitReq_37_121 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h79;
  wire          compressDataVec_hitReq_38_121 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h79;
  wire          compressDataVec_hitReq_39_121 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h79;
  wire          compressDataVec_hitReq_40_121 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h79;
  wire          compressDataVec_hitReq_41_121 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h79;
  wire          compressDataVec_hitReq_42_121 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h79;
  wire          compressDataVec_hitReq_43_121 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h79;
  wire          compressDataVec_hitReq_44_121 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h79;
  wire          compressDataVec_hitReq_45_121 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h79;
  wire          compressDataVec_hitReq_46_121 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h79;
  wire          compressDataVec_hitReq_47_121 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h79;
  wire          compressDataVec_hitReq_48_121 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h79;
  wire          compressDataVec_hitReq_49_121 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h79;
  wire          compressDataVec_hitReq_50_121 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h79;
  wire          compressDataVec_hitReq_51_121 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h79;
  wire          compressDataVec_hitReq_52_121 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h79;
  wire          compressDataVec_hitReq_53_121 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h79;
  wire          compressDataVec_hitReq_54_121 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h79;
  wire          compressDataVec_hitReq_55_121 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h79;
  wire          compressDataVec_hitReq_56_121 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h79;
  wire          compressDataVec_hitReq_57_121 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h79;
  wire          compressDataVec_hitReq_58_121 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h79;
  wire          compressDataVec_hitReq_59_121 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h79;
  wire          compressDataVec_hitReq_60_121 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h79;
  wire          compressDataVec_hitReq_61_121 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h79;
  wire          compressDataVec_hitReq_62_121 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h79;
  wire          compressDataVec_hitReq_63_121 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h79;
  wire [7:0]    compressDataVec_selectReqData_121 =
    (compressDataVec_hitReq_0_121 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_121 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_121 ? source2Pipe[23:16] : 8'h0)
    | (compressDataVec_hitReq_3_121 ? source2Pipe[31:24] : 8'h0) | (compressDataVec_hitReq_4_121 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_121 ? source2Pipe[47:40] : 8'h0)
    | (compressDataVec_hitReq_6_121 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_121 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_121 ? source2Pipe[71:64] : 8'h0)
    | (compressDataVec_hitReq_9_121 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_121 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_121 ? source2Pipe[95:88] : 8'h0)
    | (compressDataVec_hitReq_12_121 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_121 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_121 ? source2Pipe[119:112] : 8'h0)
    | (compressDataVec_hitReq_15_121 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_121 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_121 ? source2Pipe[143:136] : 8'h0)
    | (compressDataVec_hitReq_18_121 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_121 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_121 ? source2Pipe[167:160] : 8'h0)
    | (compressDataVec_hitReq_21_121 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_121 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_121 ? source2Pipe[191:184] : 8'h0)
    | (compressDataVec_hitReq_24_121 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_121 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_121 ? source2Pipe[215:208] : 8'h0)
    | (compressDataVec_hitReq_27_121 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_121 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_121 ? source2Pipe[239:232] : 8'h0)
    | (compressDataVec_hitReq_30_121 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_121 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_121 ? source2Pipe[263:256] : 8'h0)
    | (compressDataVec_hitReq_33_121 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_121 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_121 ? source2Pipe[287:280] : 8'h0)
    | (compressDataVec_hitReq_36_121 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_121 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_121 ? source2Pipe[311:304] : 8'h0)
    | (compressDataVec_hitReq_39_121 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_121 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_121 ? source2Pipe[335:328] : 8'h0)
    | (compressDataVec_hitReq_42_121 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_121 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_121 ? source2Pipe[359:352] : 8'h0)
    | (compressDataVec_hitReq_45_121 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_121 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_121 ? source2Pipe[383:376] : 8'h0)
    | (compressDataVec_hitReq_48_121 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_121 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_121 ? source2Pipe[407:400] : 8'h0)
    | (compressDataVec_hitReq_51_121 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_121 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_121 ? source2Pipe[431:424] : 8'h0)
    | (compressDataVec_hitReq_54_121 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_121 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_121 ? source2Pipe[455:448] : 8'h0)
    | (compressDataVec_hitReq_57_121 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_121 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_121 ? source2Pipe[479:472] : 8'h0)
    | (compressDataVec_hitReq_60_121 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_121 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_121 ? source2Pipe[503:496] : 8'h0)
    | (compressDataVec_hitReq_63_121 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_122 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h7A;
  wire          compressDataVec_hitReq_1_122 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h7A;
  wire          compressDataVec_hitReq_2_122 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h7A;
  wire          compressDataVec_hitReq_3_122 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h7A;
  wire          compressDataVec_hitReq_4_122 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h7A;
  wire          compressDataVec_hitReq_5_122 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h7A;
  wire          compressDataVec_hitReq_6_122 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h7A;
  wire          compressDataVec_hitReq_7_122 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h7A;
  wire          compressDataVec_hitReq_8_122 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h7A;
  wire          compressDataVec_hitReq_9_122 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h7A;
  wire          compressDataVec_hitReq_10_122 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h7A;
  wire          compressDataVec_hitReq_11_122 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h7A;
  wire          compressDataVec_hitReq_12_122 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h7A;
  wire          compressDataVec_hitReq_13_122 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h7A;
  wire          compressDataVec_hitReq_14_122 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h7A;
  wire          compressDataVec_hitReq_15_122 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h7A;
  wire          compressDataVec_hitReq_16_122 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h7A;
  wire          compressDataVec_hitReq_17_122 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h7A;
  wire          compressDataVec_hitReq_18_122 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h7A;
  wire          compressDataVec_hitReq_19_122 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h7A;
  wire          compressDataVec_hitReq_20_122 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h7A;
  wire          compressDataVec_hitReq_21_122 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h7A;
  wire          compressDataVec_hitReq_22_122 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h7A;
  wire          compressDataVec_hitReq_23_122 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h7A;
  wire          compressDataVec_hitReq_24_122 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h7A;
  wire          compressDataVec_hitReq_25_122 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h7A;
  wire          compressDataVec_hitReq_26_122 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h7A;
  wire          compressDataVec_hitReq_27_122 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h7A;
  wire          compressDataVec_hitReq_28_122 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h7A;
  wire          compressDataVec_hitReq_29_122 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h7A;
  wire          compressDataVec_hitReq_30_122 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h7A;
  wire          compressDataVec_hitReq_31_122 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h7A;
  wire          compressDataVec_hitReq_32_122 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h7A;
  wire          compressDataVec_hitReq_33_122 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h7A;
  wire          compressDataVec_hitReq_34_122 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h7A;
  wire          compressDataVec_hitReq_35_122 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h7A;
  wire          compressDataVec_hitReq_36_122 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h7A;
  wire          compressDataVec_hitReq_37_122 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h7A;
  wire          compressDataVec_hitReq_38_122 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h7A;
  wire          compressDataVec_hitReq_39_122 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h7A;
  wire          compressDataVec_hitReq_40_122 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h7A;
  wire          compressDataVec_hitReq_41_122 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h7A;
  wire          compressDataVec_hitReq_42_122 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h7A;
  wire          compressDataVec_hitReq_43_122 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h7A;
  wire          compressDataVec_hitReq_44_122 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h7A;
  wire          compressDataVec_hitReq_45_122 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h7A;
  wire          compressDataVec_hitReq_46_122 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h7A;
  wire          compressDataVec_hitReq_47_122 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h7A;
  wire          compressDataVec_hitReq_48_122 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h7A;
  wire          compressDataVec_hitReq_49_122 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h7A;
  wire          compressDataVec_hitReq_50_122 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h7A;
  wire          compressDataVec_hitReq_51_122 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h7A;
  wire          compressDataVec_hitReq_52_122 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h7A;
  wire          compressDataVec_hitReq_53_122 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h7A;
  wire          compressDataVec_hitReq_54_122 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h7A;
  wire          compressDataVec_hitReq_55_122 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h7A;
  wire          compressDataVec_hitReq_56_122 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h7A;
  wire          compressDataVec_hitReq_57_122 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h7A;
  wire          compressDataVec_hitReq_58_122 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h7A;
  wire          compressDataVec_hitReq_59_122 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h7A;
  wire          compressDataVec_hitReq_60_122 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h7A;
  wire          compressDataVec_hitReq_61_122 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h7A;
  wire          compressDataVec_hitReq_62_122 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h7A;
  wire          compressDataVec_hitReq_63_122 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h7A;
  wire [7:0]    compressDataVec_selectReqData_122 =
    (compressDataVec_hitReq_0_122 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_122 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_122 ? source2Pipe[23:16] : 8'h0)
    | (compressDataVec_hitReq_3_122 ? source2Pipe[31:24] : 8'h0) | (compressDataVec_hitReq_4_122 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_122 ? source2Pipe[47:40] : 8'h0)
    | (compressDataVec_hitReq_6_122 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_122 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_122 ? source2Pipe[71:64] : 8'h0)
    | (compressDataVec_hitReq_9_122 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_122 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_122 ? source2Pipe[95:88] : 8'h0)
    | (compressDataVec_hitReq_12_122 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_122 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_122 ? source2Pipe[119:112] : 8'h0)
    | (compressDataVec_hitReq_15_122 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_122 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_122 ? source2Pipe[143:136] : 8'h0)
    | (compressDataVec_hitReq_18_122 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_122 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_122 ? source2Pipe[167:160] : 8'h0)
    | (compressDataVec_hitReq_21_122 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_122 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_122 ? source2Pipe[191:184] : 8'h0)
    | (compressDataVec_hitReq_24_122 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_122 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_122 ? source2Pipe[215:208] : 8'h0)
    | (compressDataVec_hitReq_27_122 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_122 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_122 ? source2Pipe[239:232] : 8'h0)
    | (compressDataVec_hitReq_30_122 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_122 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_122 ? source2Pipe[263:256] : 8'h0)
    | (compressDataVec_hitReq_33_122 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_122 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_122 ? source2Pipe[287:280] : 8'h0)
    | (compressDataVec_hitReq_36_122 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_122 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_122 ? source2Pipe[311:304] : 8'h0)
    | (compressDataVec_hitReq_39_122 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_122 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_122 ? source2Pipe[335:328] : 8'h0)
    | (compressDataVec_hitReq_42_122 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_122 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_122 ? source2Pipe[359:352] : 8'h0)
    | (compressDataVec_hitReq_45_122 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_122 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_122 ? source2Pipe[383:376] : 8'h0)
    | (compressDataVec_hitReq_48_122 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_122 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_122 ? source2Pipe[407:400] : 8'h0)
    | (compressDataVec_hitReq_51_122 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_122 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_122 ? source2Pipe[431:424] : 8'h0)
    | (compressDataVec_hitReq_54_122 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_122 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_122 ? source2Pipe[455:448] : 8'h0)
    | (compressDataVec_hitReq_57_122 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_122 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_122 ? source2Pipe[479:472] : 8'h0)
    | (compressDataVec_hitReq_60_122 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_122 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_122 ? source2Pipe[503:496] : 8'h0)
    | (compressDataVec_hitReq_63_122 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_123 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h7B;
  wire          compressDataVec_hitReq_1_123 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h7B;
  wire          compressDataVec_hitReq_2_123 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h7B;
  wire          compressDataVec_hitReq_3_123 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h7B;
  wire          compressDataVec_hitReq_4_123 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h7B;
  wire          compressDataVec_hitReq_5_123 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h7B;
  wire          compressDataVec_hitReq_6_123 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h7B;
  wire          compressDataVec_hitReq_7_123 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h7B;
  wire          compressDataVec_hitReq_8_123 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h7B;
  wire          compressDataVec_hitReq_9_123 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h7B;
  wire          compressDataVec_hitReq_10_123 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h7B;
  wire          compressDataVec_hitReq_11_123 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h7B;
  wire          compressDataVec_hitReq_12_123 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h7B;
  wire          compressDataVec_hitReq_13_123 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h7B;
  wire          compressDataVec_hitReq_14_123 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h7B;
  wire          compressDataVec_hitReq_15_123 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h7B;
  wire          compressDataVec_hitReq_16_123 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h7B;
  wire          compressDataVec_hitReq_17_123 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h7B;
  wire          compressDataVec_hitReq_18_123 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h7B;
  wire          compressDataVec_hitReq_19_123 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h7B;
  wire          compressDataVec_hitReq_20_123 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h7B;
  wire          compressDataVec_hitReq_21_123 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h7B;
  wire          compressDataVec_hitReq_22_123 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h7B;
  wire          compressDataVec_hitReq_23_123 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h7B;
  wire          compressDataVec_hitReq_24_123 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h7B;
  wire          compressDataVec_hitReq_25_123 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h7B;
  wire          compressDataVec_hitReq_26_123 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h7B;
  wire          compressDataVec_hitReq_27_123 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h7B;
  wire          compressDataVec_hitReq_28_123 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h7B;
  wire          compressDataVec_hitReq_29_123 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h7B;
  wire          compressDataVec_hitReq_30_123 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h7B;
  wire          compressDataVec_hitReq_31_123 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h7B;
  wire          compressDataVec_hitReq_32_123 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h7B;
  wire          compressDataVec_hitReq_33_123 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h7B;
  wire          compressDataVec_hitReq_34_123 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h7B;
  wire          compressDataVec_hitReq_35_123 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h7B;
  wire          compressDataVec_hitReq_36_123 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h7B;
  wire          compressDataVec_hitReq_37_123 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h7B;
  wire          compressDataVec_hitReq_38_123 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h7B;
  wire          compressDataVec_hitReq_39_123 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h7B;
  wire          compressDataVec_hitReq_40_123 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h7B;
  wire          compressDataVec_hitReq_41_123 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h7B;
  wire          compressDataVec_hitReq_42_123 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h7B;
  wire          compressDataVec_hitReq_43_123 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h7B;
  wire          compressDataVec_hitReq_44_123 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h7B;
  wire          compressDataVec_hitReq_45_123 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h7B;
  wire          compressDataVec_hitReq_46_123 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h7B;
  wire          compressDataVec_hitReq_47_123 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h7B;
  wire          compressDataVec_hitReq_48_123 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h7B;
  wire          compressDataVec_hitReq_49_123 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h7B;
  wire          compressDataVec_hitReq_50_123 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h7B;
  wire          compressDataVec_hitReq_51_123 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h7B;
  wire          compressDataVec_hitReq_52_123 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h7B;
  wire          compressDataVec_hitReq_53_123 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h7B;
  wire          compressDataVec_hitReq_54_123 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h7B;
  wire          compressDataVec_hitReq_55_123 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h7B;
  wire          compressDataVec_hitReq_56_123 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h7B;
  wire          compressDataVec_hitReq_57_123 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h7B;
  wire          compressDataVec_hitReq_58_123 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h7B;
  wire          compressDataVec_hitReq_59_123 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h7B;
  wire          compressDataVec_hitReq_60_123 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h7B;
  wire          compressDataVec_hitReq_61_123 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h7B;
  wire          compressDataVec_hitReq_62_123 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h7B;
  wire          compressDataVec_hitReq_63_123 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h7B;
  wire [7:0]    compressDataVec_selectReqData_123 =
    (compressDataVec_hitReq_0_123 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_123 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_123 ? source2Pipe[23:16] : 8'h0)
    | (compressDataVec_hitReq_3_123 ? source2Pipe[31:24] : 8'h0) | (compressDataVec_hitReq_4_123 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_123 ? source2Pipe[47:40] : 8'h0)
    | (compressDataVec_hitReq_6_123 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_123 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_123 ? source2Pipe[71:64] : 8'h0)
    | (compressDataVec_hitReq_9_123 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_123 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_123 ? source2Pipe[95:88] : 8'h0)
    | (compressDataVec_hitReq_12_123 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_123 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_123 ? source2Pipe[119:112] : 8'h0)
    | (compressDataVec_hitReq_15_123 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_123 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_123 ? source2Pipe[143:136] : 8'h0)
    | (compressDataVec_hitReq_18_123 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_123 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_123 ? source2Pipe[167:160] : 8'h0)
    | (compressDataVec_hitReq_21_123 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_123 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_123 ? source2Pipe[191:184] : 8'h0)
    | (compressDataVec_hitReq_24_123 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_123 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_123 ? source2Pipe[215:208] : 8'h0)
    | (compressDataVec_hitReq_27_123 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_123 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_123 ? source2Pipe[239:232] : 8'h0)
    | (compressDataVec_hitReq_30_123 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_123 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_123 ? source2Pipe[263:256] : 8'h0)
    | (compressDataVec_hitReq_33_123 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_123 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_123 ? source2Pipe[287:280] : 8'h0)
    | (compressDataVec_hitReq_36_123 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_123 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_123 ? source2Pipe[311:304] : 8'h0)
    | (compressDataVec_hitReq_39_123 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_123 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_123 ? source2Pipe[335:328] : 8'h0)
    | (compressDataVec_hitReq_42_123 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_123 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_123 ? source2Pipe[359:352] : 8'h0)
    | (compressDataVec_hitReq_45_123 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_123 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_123 ? source2Pipe[383:376] : 8'h0)
    | (compressDataVec_hitReq_48_123 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_123 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_123 ? source2Pipe[407:400] : 8'h0)
    | (compressDataVec_hitReq_51_123 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_123 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_123 ? source2Pipe[431:424] : 8'h0)
    | (compressDataVec_hitReq_54_123 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_123 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_123 ? source2Pipe[455:448] : 8'h0)
    | (compressDataVec_hitReq_57_123 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_123 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_123 ? source2Pipe[479:472] : 8'h0)
    | (compressDataVec_hitReq_60_123 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_123 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_123 ? source2Pipe[503:496] : 8'h0)
    | (compressDataVec_hitReq_63_123 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_124 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h7C;
  wire          compressDataVec_hitReq_1_124 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h7C;
  wire          compressDataVec_hitReq_2_124 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h7C;
  wire          compressDataVec_hitReq_3_124 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h7C;
  wire          compressDataVec_hitReq_4_124 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h7C;
  wire          compressDataVec_hitReq_5_124 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h7C;
  wire          compressDataVec_hitReq_6_124 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h7C;
  wire          compressDataVec_hitReq_7_124 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h7C;
  wire          compressDataVec_hitReq_8_124 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h7C;
  wire          compressDataVec_hitReq_9_124 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h7C;
  wire          compressDataVec_hitReq_10_124 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h7C;
  wire          compressDataVec_hitReq_11_124 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h7C;
  wire          compressDataVec_hitReq_12_124 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h7C;
  wire          compressDataVec_hitReq_13_124 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h7C;
  wire          compressDataVec_hitReq_14_124 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h7C;
  wire          compressDataVec_hitReq_15_124 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h7C;
  wire          compressDataVec_hitReq_16_124 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h7C;
  wire          compressDataVec_hitReq_17_124 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h7C;
  wire          compressDataVec_hitReq_18_124 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h7C;
  wire          compressDataVec_hitReq_19_124 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h7C;
  wire          compressDataVec_hitReq_20_124 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h7C;
  wire          compressDataVec_hitReq_21_124 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h7C;
  wire          compressDataVec_hitReq_22_124 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h7C;
  wire          compressDataVec_hitReq_23_124 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h7C;
  wire          compressDataVec_hitReq_24_124 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h7C;
  wire          compressDataVec_hitReq_25_124 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h7C;
  wire          compressDataVec_hitReq_26_124 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h7C;
  wire          compressDataVec_hitReq_27_124 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h7C;
  wire          compressDataVec_hitReq_28_124 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h7C;
  wire          compressDataVec_hitReq_29_124 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h7C;
  wire          compressDataVec_hitReq_30_124 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h7C;
  wire          compressDataVec_hitReq_31_124 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h7C;
  wire          compressDataVec_hitReq_32_124 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h7C;
  wire          compressDataVec_hitReq_33_124 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h7C;
  wire          compressDataVec_hitReq_34_124 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h7C;
  wire          compressDataVec_hitReq_35_124 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h7C;
  wire          compressDataVec_hitReq_36_124 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h7C;
  wire          compressDataVec_hitReq_37_124 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h7C;
  wire          compressDataVec_hitReq_38_124 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h7C;
  wire          compressDataVec_hitReq_39_124 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h7C;
  wire          compressDataVec_hitReq_40_124 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h7C;
  wire          compressDataVec_hitReq_41_124 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h7C;
  wire          compressDataVec_hitReq_42_124 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h7C;
  wire          compressDataVec_hitReq_43_124 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h7C;
  wire          compressDataVec_hitReq_44_124 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h7C;
  wire          compressDataVec_hitReq_45_124 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h7C;
  wire          compressDataVec_hitReq_46_124 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h7C;
  wire          compressDataVec_hitReq_47_124 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h7C;
  wire          compressDataVec_hitReq_48_124 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h7C;
  wire          compressDataVec_hitReq_49_124 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h7C;
  wire          compressDataVec_hitReq_50_124 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h7C;
  wire          compressDataVec_hitReq_51_124 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h7C;
  wire          compressDataVec_hitReq_52_124 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h7C;
  wire          compressDataVec_hitReq_53_124 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h7C;
  wire          compressDataVec_hitReq_54_124 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h7C;
  wire          compressDataVec_hitReq_55_124 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h7C;
  wire          compressDataVec_hitReq_56_124 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h7C;
  wire          compressDataVec_hitReq_57_124 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h7C;
  wire          compressDataVec_hitReq_58_124 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h7C;
  wire          compressDataVec_hitReq_59_124 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h7C;
  wire          compressDataVec_hitReq_60_124 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h7C;
  wire          compressDataVec_hitReq_61_124 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h7C;
  wire          compressDataVec_hitReq_62_124 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h7C;
  wire          compressDataVec_hitReq_63_124 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h7C;
  wire [7:0]    compressDataVec_selectReqData_124 =
    (compressDataVec_hitReq_0_124 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_124 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_124 ? source2Pipe[23:16] : 8'h0)
    | (compressDataVec_hitReq_3_124 ? source2Pipe[31:24] : 8'h0) | (compressDataVec_hitReq_4_124 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_124 ? source2Pipe[47:40] : 8'h0)
    | (compressDataVec_hitReq_6_124 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_124 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_124 ? source2Pipe[71:64] : 8'h0)
    | (compressDataVec_hitReq_9_124 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_124 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_124 ? source2Pipe[95:88] : 8'h0)
    | (compressDataVec_hitReq_12_124 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_124 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_124 ? source2Pipe[119:112] : 8'h0)
    | (compressDataVec_hitReq_15_124 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_124 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_124 ? source2Pipe[143:136] : 8'h0)
    | (compressDataVec_hitReq_18_124 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_124 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_124 ? source2Pipe[167:160] : 8'h0)
    | (compressDataVec_hitReq_21_124 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_124 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_124 ? source2Pipe[191:184] : 8'h0)
    | (compressDataVec_hitReq_24_124 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_124 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_124 ? source2Pipe[215:208] : 8'h0)
    | (compressDataVec_hitReq_27_124 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_124 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_124 ? source2Pipe[239:232] : 8'h0)
    | (compressDataVec_hitReq_30_124 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_124 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_124 ? source2Pipe[263:256] : 8'h0)
    | (compressDataVec_hitReq_33_124 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_124 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_124 ? source2Pipe[287:280] : 8'h0)
    | (compressDataVec_hitReq_36_124 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_124 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_124 ? source2Pipe[311:304] : 8'h0)
    | (compressDataVec_hitReq_39_124 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_124 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_124 ? source2Pipe[335:328] : 8'h0)
    | (compressDataVec_hitReq_42_124 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_124 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_124 ? source2Pipe[359:352] : 8'h0)
    | (compressDataVec_hitReq_45_124 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_124 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_124 ? source2Pipe[383:376] : 8'h0)
    | (compressDataVec_hitReq_48_124 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_124 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_124 ? source2Pipe[407:400] : 8'h0)
    | (compressDataVec_hitReq_51_124 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_124 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_124 ? source2Pipe[431:424] : 8'h0)
    | (compressDataVec_hitReq_54_124 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_124 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_124 ? source2Pipe[455:448] : 8'h0)
    | (compressDataVec_hitReq_57_124 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_124 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_124 ? source2Pipe[479:472] : 8'h0)
    | (compressDataVec_hitReq_60_124 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_124 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_124 ? source2Pipe[503:496] : 8'h0)
    | (compressDataVec_hitReq_63_124 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_125 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h7D;
  wire          compressDataVec_hitReq_1_125 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h7D;
  wire          compressDataVec_hitReq_2_125 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h7D;
  wire          compressDataVec_hitReq_3_125 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h7D;
  wire          compressDataVec_hitReq_4_125 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h7D;
  wire          compressDataVec_hitReq_5_125 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h7D;
  wire          compressDataVec_hitReq_6_125 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h7D;
  wire          compressDataVec_hitReq_7_125 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h7D;
  wire          compressDataVec_hitReq_8_125 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h7D;
  wire          compressDataVec_hitReq_9_125 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h7D;
  wire          compressDataVec_hitReq_10_125 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h7D;
  wire          compressDataVec_hitReq_11_125 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h7D;
  wire          compressDataVec_hitReq_12_125 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h7D;
  wire          compressDataVec_hitReq_13_125 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h7D;
  wire          compressDataVec_hitReq_14_125 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h7D;
  wire          compressDataVec_hitReq_15_125 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h7D;
  wire          compressDataVec_hitReq_16_125 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h7D;
  wire          compressDataVec_hitReq_17_125 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h7D;
  wire          compressDataVec_hitReq_18_125 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h7D;
  wire          compressDataVec_hitReq_19_125 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h7D;
  wire          compressDataVec_hitReq_20_125 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h7D;
  wire          compressDataVec_hitReq_21_125 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h7D;
  wire          compressDataVec_hitReq_22_125 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h7D;
  wire          compressDataVec_hitReq_23_125 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h7D;
  wire          compressDataVec_hitReq_24_125 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h7D;
  wire          compressDataVec_hitReq_25_125 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h7D;
  wire          compressDataVec_hitReq_26_125 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h7D;
  wire          compressDataVec_hitReq_27_125 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h7D;
  wire          compressDataVec_hitReq_28_125 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h7D;
  wire          compressDataVec_hitReq_29_125 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h7D;
  wire          compressDataVec_hitReq_30_125 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h7D;
  wire          compressDataVec_hitReq_31_125 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h7D;
  wire          compressDataVec_hitReq_32_125 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h7D;
  wire          compressDataVec_hitReq_33_125 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h7D;
  wire          compressDataVec_hitReq_34_125 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h7D;
  wire          compressDataVec_hitReq_35_125 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h7D;
  wire          compressDataVec_hitReq_36_125 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h7D;
  wire          compressDataVec_hitReq_37_125 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h7D;
  wire          compressDataVec_hitReq_38_125 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h7D;
  wire          compressDataVec_hitReq_39_125 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h7D;
  wire          compressDataVec_hitReq_40_125 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h7D;
  wire          compressDataVec_hitReq_41_125 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h7D;
  wire          compressDataVec_hitReq_42_125 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h7D;
  wire          compressDataVec_hitReq_43_125 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h7D;
  wire          compressDataVec_hitReq_44_125 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h7D;
  wire          compressDataVec_hitReq_45_125 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h7D;
  wire          compressDataVec_hitReq_46_125 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h7D;
  wire          compressDataVec_hitReq_47_125 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h7D;
  wire          compressDataVec_hitReq_48_125 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h7D;
  wire          compressDataVec_hitReq_49_125 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h7D;
  wire          compressDataVec_hitReq_50_125 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h7D;
  wire          compressDataVec_hitReq_51_125 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h7D;
  wire          compressDataVec_hitReq_52_125 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h7D;
  wire          compressDataVec_hitReq_53_125 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h7D;
  wire          compressDataVec_hitReq_54_125 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h7D;
  wire          compressDataVec_hitReq_55_125 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h7D;
  wire          compressDataVec_hitReq_56_125 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h7D;
  wire          compressDataVec_hitReq_57_125 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h7D;
  wire          compressDataVec_hitReq_58_125 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h7D;
  wire          compressDataVec_hitReq_59_125 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h7D;
  wire          compressDataVec_hitReq_60_125 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h7D;
  wire          compressDataVec_hitReq_61_125 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h7D;
  wire          compressDataVec_hitReq_62_125 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h7D;
  wire          compressDataVec_hitReq_63_125 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h7D;
  wire [7:0]    compressDataVec_selectReqData_125 =
    (compressDataVec_hitReq_0_125 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_125 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_125 ? source2Pipe[23:16] : 8'h0)
    | (compressDataVec_hitReq_3_125 ? source2Pipe[31:24] : 8'h0) | (compressDataVec_hitReq_4_125 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_125 ? source2Pipe[47:40] : 8'h0)
    | (compressDataVec_hitReq_6_125 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_125 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_125 ? source2Pipe[71:64] : 8'h0)
    | (compressDataVec_hitReq_9_125 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_125 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_125 ? source2Pipe[95:88] : 8'h0)
    | (compressDataVec_hitReq_12_125 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_125 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_125 ? source2Pipe[119:112] : 8'h0)
    | (compressDataVec_hitReq_15_125 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_125 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_125 ? source2Pipe[143:136] : 8'h0)
    | (compressDataVec_hitReq_18_125 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_125 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_125 ? source2Pipe[167:160] : 8'h0)
    | (compressDataVec_hitReq_21_125 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_125 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_125 ? source2Pipe[191:184] : 8'h0)
    | (compressDataVec_hitReq_24_125 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_125 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_125 ? source2Pipe[215:208] : 8'h0)
    | (compressDataVec_hitReq_27_125 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_125 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_125 ? source2Pipe[239:232] : 8'h0)
    | (compressDataVec_hitReq_30_125 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_125 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_125 ? source2Pipe[263:256] : 8'h0)
    | (compressDataVec_hitReq_33_125 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_125 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_125 ? source2Pipe[287:280] : 8'h0)
    | (compressDataVec_hitReq_36_125 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_125 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_125 ? source2Pipe[311:304] : 8'h0)
    | (compressDataVec_hitReq_39_125 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_125 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_125 ? source2Pipe[335:328] : 8'h0)
    | (compressDataVec_hitReq_42_125 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_125 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_125 ? source2Pipe[359:352] : 8'h0)
    | (compressDataVec_hitReq_45_125 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_125 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_125 ? source2Pipe[383:376] : 8'h0)
    | (compressDataVec_hitReq_48_125 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_125 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_125 ? source2Pipe[407:400] : 8'h0)
    | (compressDataVec_hitReq_51_125 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_125 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_125 ? source2Pipe[431:424] : 8'h0)
    | (compressDataVec_hitReq_54_125 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_125 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_125 ? source2Pipe[455:448] : 8'h0)
    | (compressDataVec_hitReq_57_125 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_125 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_125 ? source2Pipe[479:472] : 8'h0)
    | (compressDataVec_hitReq_60_125 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_125 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_125 ? source2Pipe[503:496] : 8'h0)
    | (compressDataVec_hitReq_63_125 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_126 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h7E;
  wire          compressDataVec_hitReq_1_126 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h7E;
  wire          compressDataVec_hitReq_2_126 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h7E;
  wire          compressDataVec_hitReq_3_126 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h7E;
  wire          compressDataVec_hitReq_4_126 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h7E;
  wire          compressDataVec_hitReq_5_126 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h7E;
  wire          compressDataVec_hitReq_6_126 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h7E;
  wire          compressDataVec_hitReq_7_126 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h7E;
  wire          compressDataVec_hitReq_8_126 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h7E;
  wire          compressDataVec_hitReq_9_126 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h7E;
  wire          compressDataVec_hitReq_10_126 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h7E;
  wire          compressDataVec_hitReq_11_126 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h7E;
  wire          compressDataVec_hitReq_12_126 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h7E;
  wire          compressDataVec_hitReq_13_126 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h7E;
  wire          compressDataVec_hitReq_14_126 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h7E;
  wire          compressDataVec_hitReq_15_126 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h7E;
  wire          compressDataVec_hitReq_16_126 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h7E;
  wire          compressDataVec_hitReq_17_126 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h7E;
  wire          compressDataVec_hitReq_18_126 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h7E;
  wire          compressDataVec_hitReq_19_126 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h7E;
  wire          compressDataVec_hitReq_20_126 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h7E;
  wire          compressDataVec_hitReq_21_126 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h7E;
  wire          compressDataVec_hitReq_22_126 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h7E;
  wire          compressDataVec_hitReq_23_126 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h7E;
  wire          compressDataVec_hitReq_24_126 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h7E;
  wire          compressDataVec_hitReq_25_126 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h7E;
  wire          compressDataVec_hitReq_26_126 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h7E;
  wire          compressDataVec_hitReq_27_126 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h7E;
  wire          compressDataVec_hitReq_28_126 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h7E;
  wire          compressDataVec_hitReq_29_126 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h7E;
  wire          compressDataVec_hitReq_30_126 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h7E;
  wire          compressDataVec_hitReq_31_126 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h7E;
  wire          compressDataVec_hitReq_32_126 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h7E;
  wire          compressDataVec_hitReq_33_126 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h7E;
  wire          compressDataVec_hitReq_34_126 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h7E;
  wire          compressDataVec_hitReq_35_126 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h7E;
  wire          compressDataVec_hitReq_36_126 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h7E;
  wire          compressDataVec_hitReq_37_126 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h7E;
  wire          compressDataVec_hitReq_38_126 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h7E;
  wire          compressDataVec_hitReq_39_126 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h7E;
  wire          compressDataVec_hitReq_40_126 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h7E;
  wire          compressDataVec_hitReq_41_126 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h7E;
  wire          compressDataVec_hitReq_42_126 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h7E;
  wire          compressDataVec_hitReq_43_126 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h7E;
  wire          compressDataVec_hitReq_44_126 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h7E;
  wire          compressDataVec_hitReq_45_126 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h7E;
  wire          compressDataVec_hitReq_46_126 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h7E;
  wire          compressDataVec_hitReq_47_126 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h7E;
  wire          compressDataVec_hitReq_48_126 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h7E;
  wire          compressDataVec_hitReq_49_126 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h7E;
  wire          compressDataVec_hitReq_50_126 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h7E;
  wire          compressDataVec_hitReq_51_126 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h7E;
  wire          compressDataVec_hitReq_52_126 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h7E;
  wire          compressDataVec_hitReq_53_126 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h7E;
  wire          compressDataVec_hitReq_54_126 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h7E;
  wire          compressDataVec_hitReq_55_126 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h7E;
  wire          compressDataVec_hitReq_56_126 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h7E;
  wire          compressDataVec_hitReq_57_126 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h7E;
  wire          compressDataVec_hitReq_58_126 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h7E;
  wire          compressDataVec_hitReq_59_126 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h7E;
  wire          compressDataVec_hitReq_60_126 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h7E;
  wire          compressDataVec_hitReq_61_126 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h7E;
  wire          compressDataVec_hitReq_62_126 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h7E;
  wire          compressDataVec_hitReq_63_126 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h7E;
  wire [7:0]    compressDataVec_selectReqData_126 =
    (compressDataVec_hitReq_0_126 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_126 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_126 ? source2Pipe[23:16] : 8'h0)
    | (compressDataVec_hitReq_3_126 ? source2Pipe[31:24] : 8'h0) | (compressDataVec_hitReq_4_126 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_126 ? source2Pipe[47:40] : 8'h0)
    | (compressDataVec_hitReq_6_126 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_126 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_126 ? source2Pipe[71:64] : 8'h0)
    | (compressDataVec_hitReq_9_126 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_126 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_126 ? source2Pipe[95:88] : 8'h0)
    | (compressDataVec_hitReq_12_126 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_126 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_126 ? source2Pipe[119:112] : 8'h0)
    | (compressDataVec_hitReq_15_126 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_126 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_126 ? source2Pipe[143:136] : 8'h0)
    | (compressDataVec_hitReq_18_126 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_126 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_126 ? source2Pipe[167:160] : 8'h0)
    | (compressDataVec_hitReq_21_126 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_126 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_126 ? source2Pipe[191:184] : 8'h0)
    | (compressDataVec_hitReq_24_126 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_126 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_126 ? source2Pipe[215:208] : 8'h0)
    | (compressDataVec_hitReq_27_126 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_126 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_126 ? source2Pipe[239:232] : 8'h0)
    | (compressDataVec_hitReq_30_126 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_126 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_126 ? source2Pipe[263:256] : 8'h0)
    | (compressDataVec_hitReq_33_126 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_126 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_126 ? source2Pipe[287:280] : 8'h0)
    | (compressDataVec_hitReq_36_126 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_126 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_126 ? source2Pipe[311:304] : 8'h0)
    | (compressDataVec_hitReq_39_126 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_126 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_126 ? source2Pipe[335:328] : 8'h0)
    | (compressDataVec_hitReq_42_126 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_126 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_126 ? source2Pipe[359:352] : 8'h0)
    | (compressDataVec_hitReq_45_126 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_126 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_126 ? source2Pipe[383:376] : 8'h0)
    | (compressDataVec_hitReq_48_126 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_126 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_126 ? source2Pipe[407:400] : 8'h0)
    | (compressDataVec_hitReq_51_126 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_126 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_126 ? source2Pipe[431:424] : 8'h0)
    | (compressDataVec_hitReq_54_126 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_126 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_126 ? source2Pipe[455:448] : 8'h0)
    | (compressDataVec_hitReq_57_126 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_126 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_126 ? source2Pipe[479:472] : 8'h0)
    | (compressDataVec_hitReq_60_126 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_126 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_126 ? source2Pipe[503:496] : 8'h0)
    | (compressDataVec_hitReq_63_126 ? source2Pipe[511:504] : 8'h0);
  wire          compressDataVec_hitReq_0_127 = compressMaskVecPipe_0 & compressVecPipe_0 == 11'h7F;
  wire          compressDataVec_hitReq_1_127 = compressMaskVecPipe_1 & compressVecPipe_1 == 11'h7F;
  wire          compressDataVec_hitReq_2_127 = compressMaskVecPipe_2 & compressVecPipe_2 == 11'h7F;
  wire          compressDataVec_hitReq_3_127 = compressMaskVecPipe_3 & compressVecPipe_3 == 11'h7F;
  wire          compressDataVec_hitReq_4_127 = compressMaskVecPipe_4 & compressVecPipe_4 == 11'h7F;
  wire          compressDataVec_hitReq_5_127 = compressMaskVecPipe_5 & compressVecPipe_5 == 11'h7F;
  wire          compressDataVec_hitReq_6_127 = compressMaskVecPipe_6 & compressVecPipe_6 == 11'h7F;
  wire          compressDataVec_hitReq_7_127 = compressMaskVecPipe_7 & compressVecPipe_7 == 11'h7F;
  wire          compressDataVec_hitReq_8_127 = compressMaskVecPipe_8 & compressVecPipe_8 == 11'h7F;
  wire          compressDataVec_hitReq_9_127 = compressMaskVecPipe_9 & compressVecPipe_9 == 11'h7F;
  wire          compressDataVec_hitReq_10_127 = compressMaskVecPipe_10 & compressVecPipe_10 == 11'h7F;
  wire          compressDataVec_hitReq_11_127 = compressMaskVecPipe_11 & compressVecPipe_11 == 11'h7F;
  wire          compressDataVec_hitReq_12_127 = compressMaskVecPipe_12 & compressVecPipe_12 == 11'h7F;
  wire          compressDataVec_hitReq_13_127 = compressMaskVecPipe_13 & compressVecPipe_13 == 11'h7F;
  wire          compressDataVec_hitReq_14_127 = compressMaskVecPipe_14 & compressVecPipe_14 == 11'h7F;
  wire          compressDataVec_hitReq_15_127 = compressMaskVecPipe_15 & compressVecPipe_15 == 11'h7F;
  wire          compressDataVec_hitReq_16_127 = compressMaskVecPipe_16 & compressVecPipe_16 == 11'h7F;
  wire          compressDataVec_hitReq_17_127 = compressMaskVecPipe_17 & compressVecPipe_17 == 11'h7F;
  wire          compressDataVec_hitReq_18_127 = compressMaskVecPipe_18 & compressVecPipe_18 == 11'h7F;
  wire          compressDataVec_hitReq_19_127 = compressMaskVecPipe_19 & compressVecPipe_19 == 11'h7F;
  wire          compressDataVec_hitReq_20_127 = compressMaskVecPipe_20 & compressVecPipe_20 == 11'h7F;
  wire          compressDataVec_hitReq_21_127 = compressMaskVecPipe_21 & compressVecPipe_21 == 11'h7F;
  wire          compressDataVec_hitReq_22_127 = compressMaskVecPipe_22 & compressVecPipe_22 == 11'h7F;
  wire          compressDataVec_hitReq_23_127 = compressMaskVecPipe_23 & compressVecPipe_23 == 11'h7F;
  wire          compressDataVec_hitReq_24_127 = compressMaskVecPipe_24 & compressVecPipe_24 == 11'h7F;
  wire          compressDataVec_hitReq_25_127 = compressMaskVecPipe_25 & compressVecPipe_25 == 11'h7F;
  wire          compressDataVec_hitReq_26_127 = compressMaskVecPipe_26 & compressVecPipe_26 == 11'h7F;
  wire          compressDataVec_hitReq_27_127 = compressMaskVecPipe_27 & compressVecPipe_27 == 11'h7F;
  wire          compressDataVec_hitReq_28_127 = compressMaskVecPipe_28 & compressVecPipe_28 == 11'h7F;
  wire          compressDataVec_hitReq_29_127 = compressMaskVecPipe_29 & compressVecPipe_29 == 11'h7F;
  wire          compressDataVec_hitReq_30_127 = compressMaskVecPipe_30 & compressVecPipe_30 == 11'h7F;
  wire          compressDataVec_hitReq_31_127 = compressMaskVecPipe_31 & compressVecPipe_31 == 11'h7F;
  wire          compressDataVec_hitReq_32_127 = compressMaskVecPipe_32 & compressVecPipe_32 == 11'h7F;
  wire          compressDataVec_hitReq_33_127 = compressMaskVecPipe_33 & compressVecPipe_33 == 11'h7F;
  wire          compressDataVec_hitReq_34_127 = compressMaskVecPipe_34 & compressVecPipe_34 == 11'h7F;
  wire          compressDataVec_hitReq_35_127 = compressMaskVecPipe_35 & compressVecPipe_35 == 11'h7F;
  wire          compressDataVec_hitReq_36_127 = compressMaskVecPipe_36 & compressVecPipe_36 == 11'h7F;
  wire          compressDataVec_hitReq_37_127 = compressMaskVecPipe_37 & compressVecPipe_37 == 11'h7F;
  wire          compressDataVec_hitReq_38_127 = compressMaskVecPipe_38 & compressVecPipe_38 == 11'h7F;
  wire          compressDataVec_hitReq_39_127 = compressMaskVecPipe_39 & compressVecPipe_39 == 11'h7F;
  wire          compressDataVec_hitReq_40_127 = compressMaskVecPipe_40 & compressVecPipe_40 == 11'h7F;
  wire          compressDataVec_hitReq_41_127 = compressMaskVecPipe_41 & compressVecPipe_41 == 11'h7F;
  wire          compressDataVec_hitReq_42_127 = compressMaskVecPipe_42 & compressVecPipe_42 == 11'h7F;
  wire          compressDataVec_hitReq_43_127 = compressMaskVecPipe_43 & compressVecPipe_43 == 11'h7F;
  wire          compressDataVec_hitReq_44_127 = compressMaskVecPipe_44 & compressVecPipe_44 == 11'h7F;
  wire          compressDataVec_hitReq_45_127 = compressMaskVecPipe_45 & compressVecPipe_45 == 11'h7F;
  wire          compressDataVec_hitReq_46_127 = compressMaskVecPipe_46 & compressVecPipe_46 == 11'h7F;
  wire          compressDataVec_hitReq_47_127 = compressMaskVecPipe_47 & compressVecPipe_47 == 11'h7F;
  wire          compressDataVec_hitReq_48_127 = compressMaskVecPipe_48 & compressVecPipe_48 == 11'h7F;
  wire          compressDataVec_hitReq_49_127 = compressMaskVecPipe_49 & compressVecPipe_49 == 11'h7F;
  wire          compressDataVec_hitReq_50_127 = compressMaskVecPipe_50 & compressVecPipe_50 == 11'h7F;
  wire          compressDataVec_hitReq_51_127 = compressMaskVecPipe_51 & compressVecPipe_51 == 11'h7F;
  wire          compressDataVec_hitReq_52_127 = compressMaskVecPipe_52 & compressVecPipe_52 == 11'h7F;
  wire          compressDataVec_hitReq_53_127 = compressMaskVecPipe_53 & compressVecPipe_53 == 11'h7F;
  wire          compressDataVec_hitReq_54_127 = compressMaskVecPipe_54 & compressVecPipe_54 == 11'h7F;
  wire          compressDataVec_hitReq_55_127 = compressMaskVecPipe_55 & compressVecPipe_55 == 11'h7F;
  wire          compressDataVec_hitReq_56_127 = compressMaskVecPipe_56 & compressVecPipe_56 == 11'h7F;
  wire          compressDataVec_hitReq_57_127 = compressMaskVecPipe_57 & compressVecPipe_57 == 11'h7F;
  wire          compressDataVec_hitReq_58_127 = compressMaskVecPipe_58 & compressVecPipe_58 == 11'h7F;
  wire          compressDataVec_hitReq_59_127 = compressMaskVecPipe_59 & compressVecPipe_59 == 11'h7F;
  wire          compressDataVec_hitReq_60_127 = compressMaskVecPipe_60 & compressVecPipe_60 == 11'h7F;
  wire          compressDataVec_hitReq_61_127 = compressMaskVecPipe_61 & compressVecPipe_61 == 11'h7F;
  wire          compressDataVec_hitReq_62_127 = compressMaskVecPipe_62 & compressVecPipe_62 == 11'h7F;
  wire          compressDataVec_hitReq_63_127 = compressMaskVecPipe_63 & compressVecPipe_63 == 11'h7F;
  wire [7:0]    compressDataVec_selectReqData_127 =
    (compressDataVec_hitReq_0_127 ? source2Pipe[7:0] : 8'h0) | (compressDataVec_hitReq_1_127 ? source2Pipe[15:8] : 8'h0) | (compressDataVec_hitReq_2_127 ? source2Pipe[23:16] : 8'h0)
    | (compressDataVec_hitReq_3_127 ? source2Pipe[31:24] : 8'h0) | (compressDataVec_hitReq_4_127 ? source2Pipe[39:32] : 8'h0) | (compressDataVec_hitReq_5_127 ? source2Pipe[47:40] : 8'h0)
    | (compressDataVec_hitReq_6_127 ? source2Pipe[55:48] : 8'h0) | (compressDataVec_hitReq_7_127 ? source2Pipe[63:56] : 8'h0) | (compressDataVec_hitReq_8_127 ? source2Pipe[71:64] : 8'h0)
    | (compressDataVec_hitReq_9_127 ? source2Pipe[79:72] : 8'h0) | (compressDataVec_hitReq_10_127 ? source2Pipe[87:80] : 8'h0) | (compressDataVec_hitReq_11_127 ? source2Pipe[95:88] : 8'h0)
    | (compressDataVec_hitReq_12_127 ? source2Pipe[103:96] : 8'h0) | (compressDataVec_hitReq_13_127 ? source2Pipe[111:104] : 8'h0) | (compressDataVec_hitReq_14_127 ? source2Pipe[119:112] : 8'h0)
    | (compressDataVec_hitReq_15_127 ? source2Pipe[127:120] : 8'h0) | (compressDataVec_hitReq_16_127 ? source2Pipe[135:128] : 8'h0) | (compressDataVec_hitReq_17_127 ? source2Pipe[143:136] : 8'h0)
    | (compressDataVec_hitReq_18_127 ? source2Pipe[151:144] : 8'h0) | (compressDataVec_hitReq_19_127 ? source2Pipe[159:152] : 8'h0) | (compressDataVec_hitReq_20_127 ? source2Pipe[167:160] : 8'h0)
    | (compressDataVec_hitReq_21_127 ? source2Pipe[175:168] : 8'h0) | (compressDataVec_hitReq_22_127 ? source2Pipe[183:176] : 8'h0) | (compressDataVec_hitReq_23_127 ? source2Pipe[191:184] : 8'h0)
    | (compressDataVec_hitReq_24_127 ? source2Pipe[199:192] : 8'h0) | (compressDataVec_hitReq_25_127 ? source2Pipe[207:200] : 8'h0) | (compressDataVec_hitReq_26_127 ? source2Pipe[215:208] : 8'h0)
    | (compressDataVec_hitReq_27_127 ? source2Pipe[223:216] : 8'h0) | (compressDataVec_hitReq_28_127 ? source2Pipe[231:224] : 8'h0) | (compressDataVec_hitReq_29_127 ? source2Pipe[239:232] : 8'h0)
    | (compressDataVec_hitReq_30_127 ? source2Pipe[247:240] : 8'h0) | (compressDataVec_hitReq_31_127 ? source2Pipe[255:248] : 8'h0) | (compressDataVec_hitReq_32_127 ? source2Pipe[263:256] : 8'h0)
    | (compressDataVec_hitReq_33_127 ? source2Pipe[271:264] : 8'h0) | (compressDataVec_hitReq_34_127 ? source2Pipe[279:272] : 8'h0) | (compressDataVec_hitReq_35_127 ? source2Pipe[287:280] : 8'h0)
    | (compressDataVec_hitReq_36_127 ? source2Pipe[295:288] : 8'h0) | (compressDataVec_hitReq_37_127 ? source2Pipe[303:296] : 8'h0) | (compressDataVec_hitReq_38_127 ? source2Pipe[311:304] : 8'h0)
    | (compressDataVec_hitReq_39_127 ? source2Pipe[319:312] : 8'h0) | (compressDataVec_hitReq_40_127 ? source2Pipe[327:320] : 8'h0) | (compressDataVec_hitReq_41_127 ? source2Pipe[335:328] : 8'h0)
    | (compressDataVec_hitReq_42_127 ? source2Pipe[343:336] : 8'h0) | (compressDataVec_hitReq_43_127 ? source2Pipe[351:344] : 8'h0) | (compressDataVec_hitReq_44_127 ? source2Pipe[359:352] : 8'h0)
    | (compressDataVec_hitReq_45_127 ? source2Pipe[367:360] : 8'h0) | (compressDataVec_hitReq_46_127 ? source2Pipe[375:368] : 8'h0) | (compressDataVec_hitReq_47_127 ? source2Pipe[383:376] : 8'h0)
    | (compressDataVec_hitReq_48_127 ? source2Pipe[391:384] : 8'h0) | (compressDataVec_hitReq_49_127 ? source2Pipe[399:392] : 8'h0) | (compressDataVec_hitReq_50_127 ? source2Pipe[407:400] : 8'h0)
    | (compressDataVec_hitReq_51_127 ? source2Pipe[415:408] : 8'h0) | (compressDataVec_hitReq_52_127 ? source2Pipe[423:416] : 8'h0) | (compressDataVec_hitReq_53_127 ? source2Pipe[431:424] : 8'h0)
    | (compressDataVec_hitReq_54_127 ? source2Pipe[439:432] : 8'h0) | (compressDataVec_hitReq_55_127 ? source2Pipe[447:440] : 8'h0) | (compressDataVec_hitReq_56_127 ? source2Pipe[455:448] : 8'h0)
    | (compressDataVec_hitReq_57_127 ? source2Pipe[463:456] : 8'h0) | (compressDataVec_hitReq_58_127 ? source2Pipe[471:464] : 8'h0) | (compressDataVec_hitReq_59_127 ? source2Pipe[479:472] : 8'h0)
    | (compressDataVec_hitReq_60_127 ? source2Pipe[487:480] : 8'h0) | (compressDataVec_hitReq_61_127 ? source2Pipe[495:488] : 8'h0) | (compressDataVec_hitReq_62_127 ? source2Pipe[503:496] : 8'h0)
    | (compressDataVec_hitReq_63_127 ? source2Pipe[511:504] : 8'h0);
  wire [15:0]   compressDataVec_lo_lo_lo_lo_lo_lo = {compressDataVec_useTail_1 ? compressDataReg[15:8] : compressDataVec_selectReqData_1, compressDataVec_useTail ? compressDataReg[7:0] : compressDataVec_selectReqData};
  wire [15:0]   compressDataVec_lo_lo_lo_lo_lo_hi = {compressDataVec_useTail_3 ? compressDataReg[31:24] : compressDataVec_selectReqData_3, compressDataVec_useTail_2 ? compressDataReg[23:16] : compressDataVec_selectReqData_2};
  wire [31:0]   compressDataVec_lo_lo_lo_lo_lo = {compressDataVec_lo_lo_lo_lo_lo_hi, compressDataVec_lo_lo_lo_lo_lo_lo};
  wire [15:0]   compressDataVec_lo_lo_lo_lo_hi_lo = {compressDataVec_useTail_5 ? compressDataReg[47:40] : compressDataVec_selectReqData_5, compressDataVec_useTail_4 ? compressDataReg[39:32] : compressDataVec_selectReqData_4};
  wire [15:0]   compressDataVec_lo_lo_lo_lo_hi_hi = {compressDataVec_useTail_7 ? compressDataReg[63:56] : compressDataVec_selectReqData_7, compressDataVec_useTail_6 ? compressDataReg[55:48] : compressDataVec_selectReqData_6};
  wire [31:0]   compressDataVec_lo_lo_lo_lo_hi = {compressDataVec_lo_lo_lo_lo_hi_hi, compressDataVec_lo_lo_lo_lo_hi_lo};
  wire [63:0]   compressDataVec_lo_lo_lo_lo = {compressDataVec_lo_lo_lo_lo_hi, compressDataVec_lo_lo_lo_lo_lo};
  wire [15:0]   compressDataVec_lo_lo_lo_hi_lo_lo = {compressDataVec_useTail_9 ? compressDataReg[79:72] : compressDataVec_selectReqData_9, compressDataVec_useTail_8 ? compressDataReg[71:64] : compressDataVec_selectReqData_8};
  wire [15:0]   compressDataVec_lo_lo_lo_hi_lo_hi = {compressDataVec_useTail_11 ? compressDataReg[95:88] : compressDataVec_selectReqData_11, compressDataVec_useTail_10 ? compressDataReg[87:80] : compressDataVec_selectReqData_10};
  wire [31:0]   compressDataVec_lo_lo_lo_hi_lo = {compressDataVec_lo_lo_lo_hi_lo_hi, compressDataVec_lo_lo_lo_hi_lo_lo};
  wire [15:0]   compressDataVec_lo_lo_lo_hi_hi_lo = {compressDataVec_useTail_13 ? compressDataReg[111:104] : compressDataVec_selectReqData_13, compressDataVec_useTail_12 ? compressDataReg[103:96] : compressDataVec_selectReqData_12};
  wire [15:0]   compressDataVec_lo_lo_lo_hi_hi_hi = {compressDataVec_useTail_15 ? compressDataReg[127:120] : compressDataVec_selectReqData_15, compressDataVec_useTail_14 ? compressDataReg[119:112] : compressDataVec_selectReqData_14};
  wire [31:0]   compressDataVec_lo_lo_lo_hi_hi = {compressDataVec_lo_lo_lo_hi_hi_hi, compressDataVec_lo_lo_lo_hi_hi_lo};
  wire [63:0]   compressDataVec_lo_lo_lo_hi = {compressDataVec_lo_lo_lo_hi_hi, compressDataVec_lo_lo_lo_hi_lo};
  wire [127:0]  compressDataVec_lo_lo_lo = {compressDataVec_lo_lo_lo_hi, compressDataVec_lo_lo_lo_lo};
  wire [15:0]   compressDataVec_lo_lo_hi_lo_lo_lo = {compressDataVec_useTail_17 ? compressDataReg[143:136] : compressDataVec_selectReqData_17, compressDataVec_useTail_16 ? compressDataReg[135:128] : compressDataVec_selectReqData_16};
  wire [15:0]   compressDataVec_lo_lo_hi_lo_lo_hi = {compressDataVec_useTail_19 ? compressDataReg[159:152] : compressDataVec_selectReqData_19, compressDataVec_useTail_18 ? compressDataReg[151:144] : compressDataVec_selectReqData_18};
  wire [31:0]   compressDataVec_lo_lo_hi_lo_lo = {compressDataVec_lo_lo_hi_lo_lo_hi, compressDataVec_lo_lo_hi_lo_lo_lo};
  wire [15:0]   compressDataVec_lo_lo_hi_lo_hi_lo = {compressDataVec_useTail_21 ? compressDataReg[175:168] : compressDataVec_selectReqData_21, compressDataVec_useTail_20 ? compressDataReg[167:160] : compressDataVec_selectReqData_20};
  wire [15:0]   compressDataVec_lo_lo_hi_lo_hi_hi = {compressDataVec_useTail_23 ? compressDataReg[191:184] : compressDataVec_selectReqData_23, compressDataVec_useTail_22 ? compressDataReg[183:176] : compressDataVec_selectReqData_22};
  wire [31:0]   compressDataVec_lo_lo_hi_lo_hi = {compressDataVec_lo_lo_hi_lo_hi_hi, compressDataVec_lo_lo_hi_lo_hi_lo};
  wire [63:0]   compressDataVec_lo_lo_hi_lo = {compressDataVec_lo_lo_hi_lo_hi, compressDataVec_lo_lo_hi_lo_lo};
  wire [15:0]   compressDataVec_lo_lo_hi_hi_lo_lo = {compressDataVec_useTail_25 ? compressDataReg[207:200] : compressDataVec_selectReqData_25, compressDataVec_useTail_24 ? compressDataReg[199:192] : compressDataVec_selectReqData_24};
  wire [15:0]   compressDataVec_lo_lo_hi_hi_lo_hi = {compressDataVec_useTail_27 ? compressDataReg[223:216] : compressDataVec_selectReqData_27, compressDataVec_useTail_26 ? compressDataReg[215:208] : compressDataVec_selectReqData_26};
  wire [31:0]   compressDataVec_lo_lo_hi_hi_lo = {compressDataVec_lo_lo_hi_hi_lo_hi, compressDataVec_lo_lo_hi_hi_lo_lo};
  wire [15:0]   compressDataVec_lo_lo_hi_hi_hi_lo = {compressDataVec_useTail_29 ? compressDataReg[239:232] : compressDataVec_selectReqData_29, compressDataVec_useTail_28 ? compressDataReg[231:224] : compressDataVec_selectReqData_28};
  wire [15:0]   compressDataVec_lo_lo_hi_hi_hi_hi = {compressDataVec_useTail_31 ? compressDataReg[255:248] : compressDataVec_selectReqData_31, compressDataVec_useTail_30 ? compressDataReg[247:240] : compressDataVec_selectReqData_30};
  wire [31:0]   compressDataVec_lo_lo_hi_hi_hi = {compressDataVec_lo_lo_hi_hi_hi_hi, compressDataVec_lo_lo_hi_hi_hi_lo};
  wire [63:0]   compressDataVec_lo_lo_hi_hi = {compressDataVec_lo_lo_hi_hi_hi, compressDataVec_lo_lo_hi_hi_lo};
  wire [127:0]  compressDataVec_lo_lo_hi = {compressDataVec_lo_lo_hi_hi, compressDataVec_lo_lo_hi_lo};
  wire [255:0]  compressDataVec_lo_lo = {compressDataVec_lo_lo_hi, compressDataVec_lo_lo_lo};
  wire [15:0]   compressDataVec_lo_hi_lo_lo_lo_lo = {compressDataVec_useTail_33 ? compressDataReg[271:264] : compressDataVec_selectReqData_33, compressDataVec_useTail_32 ? compressDataReg[263:256] : compressDataVec_selectReqData_32};
  wire [15:0]   compressDataVec_lo_hi_lo_lo_lo_hi = {compressDataVec_useTail_35 ? compressDataReg[287:280] : compressDataVec_selectReqData_35, compressDataVec_useTail_34 ? compressDataReg[279:272] : compressDataVec_selectReqData_34};
  wire [31:0]   compressDataVec_lo_hi_lo_lo_lo = {compressDataVec_lo_hi_lo_lo_lo_hi, compressDataVec_lo_hi_lo_lo_lo_lo};
  wire [15:0]   compressDataVec_lo_hi_lo_lo_hi_lo = {compressDataVec_useTail_37 ? compressDataReg[303:296] : compressDataVec_selectReqData_37, compressDataVec_useTail_36 ? compressDataReg[295:288] : compressDataVec_selectReqData_36};
  wire [15:0]   compressDataVec_lo_hi_lo_lo_hi_hi = {compressDataVec_useTail_39 ? compressDataReg[319:312] : compressDataVec_selectReqData_39, compressDataVec_useTail_38 ? compressDataReg[311:304] : compressDataVec_selectReqData_38};
  wire [31:0]   compressDataVec_lo_hi_lo_lo_hi = {compressDataVec_lo_hi_lo_lo_hi_hi, compressDataVec_lo_hi_lo_lo_hi_lo};
  wire [63:0]   compressDataVec_lo_hi_lo_lo = {compressDataVec_lo_hi_lo_lo_hi, compressDataVec_lo_hi_lo_lo_lo};
  wire [15:0]   compressDataVec_lo_hi_lo_hi_lo_lo = {compressDataVec_useTail_41 ? compressDataReg[335:328] : compressDataVec_selectReqData_41, compressDataVec_useTail_40 ? compressDataReg[327:320] : compressDataVec_selectReqData_40};
  wire [15:0]   compressDataVec_lo_hi_lo_hi_lo_hi = {compressDataVec_useTail_43 ? compressDataReg[351:344] : compressDataVec_selectReqData_43, compressDataVec_useTail_42 ? compressDataReg[343:336] : compressDataVec_selectReqData_42};
  wire [31:0]   compressDataVec_lo_hi_lo_hi_lo = {compressDataVec_lo_hi_lo_hi_lo_hi, compressDataVec_lo_hi_lo_hi_lo_lo};
  wire [15:0]   compressDataVec_lo_hi_lo_hi_hi_lo = {compressDataVec_useTail_45 ? compressDataReg[367:360] : compressDataVec_selectReqData_45, compressDataVec_useTail_44 ? compressDataReg[359:352] : compressDataVec_selectReqData_44};
  wire [15:0]   compressDataVec_lo_hi_lo_hi_hi_hi = {compressDataVec_useTail_47 ? compressDataReg[383:376] : compressDataVec_selectReqData_47, compressDataVec_useTail_46 ? compressDataReg[375:368] : compressDataVec_selectReqData_46};
  wire [31:0]   compressDataVec_lo_hi_lo_hi_hi = {compressDataVec_lo_hi_lo_hi_hi_hi, compressDataVec_lo_hi_lo_hi_hi_lo};
  wire [63:0]   compressDataVec_lo_hi_lo_hi = {compressDataVec_lo_hi_lo_hi_hi, compressDataVec_lo_hi_lo_hi_lo};
  wire [127:0]  compressDataVec_lo_hi_lo = {compressDataVec_lo_hi_lo_hi, compressDataVec_lo_hi_lo_lo};
  wire [15:0]   compressDataVec_lo_hi_hi_lo_lo_lo = {compressDataVec_useTail_49 ? compressDataReg[399:392] : compressDataVec_selectReqData_49, compressDataVec_useTail_48 ? compressDataReg[391:384] : compressDataVec_selectReqData_48};
  wire [15:0]   compressDataVec_lo_hi_hi_lo_lo_hi = {compressDataVec_useTail_51 ? compressDataReg[415:408] : compressDataVec_selectReqData_51, compressDataVec_useTail_50 ? compressDataReg[407:400] : compressDataVec_selectReqData_50};
  wire [31:0]   compressDataVec_lo_hi_hi_lo_lo = {compressDataVec_lo_hi_hi_lo_lo_hi, compressDataVec_lo_hi_hi_lo_lo_lo};
  wire [15:0]   compressDataVec_lo_hi_hi_lo_hi_lo = {compressDataVec_useTail_53 ? compressDataReg[431:424] : compressDataVec_selectReqData_53, compressDataVec_useTail_52 ? compressDataReg[423:416] : compressDataVec_selectReqData_52};
  wire [15:0]   compressDataVec_lo_hi_hi_lo_hi_hi = {compressDataVec_useTail_55 ? compressDataReg[447:440] : compressDataVec_selectReqData_55, compressDataVec_useTail_54 ? compressDataReg[439:432] : compressDataVec_selectReqData_54};
  wire [31:0]   compressDataVec_lo_hi_hi_lo_hi = {compressDataVec_lo_hi_hi_lo_hi_hi, compressDataVec_lo_hi_hi_lo_hi_lo};
  wire [63:0]   compressDataVec_lo_hi_hi_lo = {compressDataVec_lo_hi_hi_lo_hi, compressDataVec_lo_hi_hi_lo_lo};
  wire [15:0]   compressDataVec_lo_hi_hi_hi_lo_lo = {compressDataVec_useTail_57 ? compressDataReg[463:456] : compressDataVec_selectReqData_57, compressDataVec_useTail_56 ? compressDataReg[455:448] : compressDataVec_selectReqData_56};
  wire [15:0]   compressDataVec_lo_hi_hi_hi_lo_hi = {compressDataVec_useTail_59 ? compressDataReg[479:472] : compressDataVec_selectReqData_59, compressDataVec_useTail_58 ? compressDataReg[471:464] : compressDataVec_selectReqData_58};
  wire [31:0]   compressDataVec_lo_hi_hi_hi_lo = {compressDataVec_lo_hi_hi_hi_lo_hi, compressDataVec_lo_hi_hi_hi_lo_lo};
  wire [15:0]   compressDataVec_lo_hi_hi_hi_hi_lo = {compressDataVec_useTail_61 ? compressDataReg[495:488] : compressDataVec_selectReqData_61, compressDataVec_useTail_60 ? compressDataReg[487:480] : compressDataVec_selectReqData_60};
  wire [15:0]   compressDataVec_lo_hi_hi_hi_hi_hi = {compressDataVec_selectReqData_63, compressDataVec_useTail_62 ? compressDataReg[503:496] : compressDataVec_selectReqData_62};
  wire [31:0]   compressDataVec_lo_hi_hi_hi_hi = {compressDataVec_lo_hi_hi_hi_hi_hi, compressDataVec_lo_hi_hi_hi_hi_lo};
  wire [63:0]   compressDataVec_lo_hi_hi_hi = {compressDataVec_lo_hi_hi_hi_hi, compressDataVec_lo_hi_hi_hi_lo};
  wire [127:0]  compressDataVec_lo_hi_hi = {compressDataVec_lo_hi_hi_hi, compressDataVec_lo_hi_hi_lo};
  wire [255:0]  compressDataVec_lo_hi = {compressDataVec_lo_hi_hi, compressDataVec_lo_hi_lo};
  wire [511:0]  compressDataVec_lo = {compressDataVec_lo_hi, compressDataVec_lo_lo};
  wire [15:0]   compressDataVec_hi_lo_lo_lo_lo_lo = {compressDataVec_selectReqData_65, compressDataVec_selectReqData_64};
  wire [15:0]   compressDataVec_hi_lo_lo_lo_lo_hi = {compressDataVec_selectReqData_67, compressDataVec_selectReqData_66};
  wire [31:0]   compressDataVec_hi_lo_lo_lo_lo = {compressDataVec_hi_lo_lo_lo_lo_hi, compressDataVec_hi_lo_lo_lo_lo_lo};
  wire [15:0]   compressDataVec_hi_lo_lo_lo_hi_lo = {compressDataVec_selectReqData_69, compressDataVec_selectReqData_68};
  wire [15:0]   compressDataVec_hi_lo_lo_lo_hi_hi = {compressDataVec_selectReqData_71, compressDataVec_selectReqData_70};
  wire [31:0]   compressDataVec_hi_lo_lo_lo_hi = {compressDataVec_hi_lo_lo_lo_hi_hi, compressDataVec_hi_lo_lo_lo_hi_lo};
  wire [63:0]   compressDataVec_hi_lo_lo_lo = {compressDataVec_hi_lo_lo_lo_hi, compressDataVec_hi_lo_lo_lo_lo};
  wire [15:0]   compressDataVec_hi_lo_lo_hi_lo_lo = {compressDataVec_selectReqData_73, compressDataVec_selectReqData_72};
  wire [15:0]   compressDataVec_hi_lo_lo_hi_lo_hi = {compressDataVec_selectReqData_75, compressDataVec_selectReqData_74};
  wire [31:0]   compressDataVec_hi_lo_lo_hi_lo = {compressDataVec_hi_lo_lo_hi_lo_hi, compressDataVec_hi_lo_lo_hi_lo_lo};
  wire [15:0]   compressDataVec_hi_lo_lo_hi_hi_lo = {compressDataVec_selectReqData_77, compressDataVec_selectReqData_76};
  wire [15:0]   compressDataVec_hi_lo_lo_hi_hi_hi = {compressDataVec_selectReqData_79, compressDataVec_selectReqData_78};
  wire [31:0]   compressDataVec_hi_lo_lo_hi_hi = {compressDataVec_hi_lo_lo_hi_hi_hi, compressDataVec_hi_lo_lo_hi_hi_lo};
  wire [63:0]   compressDataVec_hi_lo_lo_hi = {compressDataVec_hi_lo_lo_hi_hi, compressDataVec_hi_lo_lo_hi_lo};
  wire [127:0]  compressDataVec_hi_lo_lo = {compressDataVec_hi_lo_lo_hi, compressDataVec_hi_lo_lo_lo};
  wire [15:0]   compressDataVec_hi_lo_hi_lo_lo_lo = {compressDataVec_selectReqData_81, compressDataVec_selectReqData_80};
  wire [15:0]   compressDataVec_hi_lo_hi_lo_lo_hi = {compressDataVec_selectReqData_83, compressDataVec_selectReqData_82};
  wire [31:0]   compressDataVec_hi_lo_hi_lo_lo = {compressDataVec_hi_lo_hi_lo_lo_hi, compressDataVec_hi_lo_hi_lo_lo_lo};
  wire [15:0]   compressDataVec_hi_lo_hi_lo_hi_lo = {compressDataVec_selectReqData_85, compressDataVec_selectReqData_84};
  wire [15:0]   compressDataVec_hi_lo_hi_lo_hi_hi = {compressDataVec_selectReqData_87, compressDataVec_selectReqData_86};
  wire [31:0]   compressDataVec_hi_lo_hi_lo_hi = {compressDataVec_hi_lo_hi_lo_hi_hi, compressDataVec_hi_lo_hi_lo_hi_lo};
  wire [63:0]   compressDataVec_hi_lo_hi_lo = {compressDataVec_hi_lo_hi_lo_hi, compressDataVec_hi_lo_hi_lo_lo};
  wire [15:0]   compressDataVec_hi_lo_hi_hi_lo_lo = {compressDataVec_selectReqData_89, compressDataVec_selectReqData_88};
  wire [15:0]   compressDataVec_hi_lo_hi_hi_lo_hi = {compressDataVec_selectReqData_91, compressDataVec_selectReqData_90};
  wire [31:0]   compressDataVec_hi_lo_hi_hi_lo = {compressDataVec_hi_lo_hi_hi_lo_hi, compressDataVec_hi_lo_hi_hi_lo_lo};
  wire [15:0]   compressDataVec_hi_lo_hi_hi_hi_lo = {compressDataVec_selectReqData_93, compressDataVec_selectReqData_92};
  wire [15:0]   compressDataVec_hi_lo_hi_hi_hi_hi = {compressDataVec_selectReqData_95, compressDataVec_selectReqData_94};
  wire [31:0]   compressDataVec_hi_lo_hi_hi_hi = {compressDataVec_hi_lo_hi_hi_hi_hi, compressDataVec_hi_lo_hi_hi_hi_lo};
  wire [63:0]   compressDataVec_hi_lo_hi_hi = {compressDataVec_hi_lo_hi_hi_hi, compressDataVec_hi_lo_hi_hi_lo};
  wire [127:0]  compressDataVec_hi_lo_hi = {compressDataVec_hi_lo_hi_hi, compressDataVec_hi_lo_hi_lo};
  wire [255:0]  compressDataVec_hi_lo = {compressDataVec_hi_lo_hi, compressDataVec_hi_lo_lo};
  wire [15:0]   compressDataVec_hi_hi_lo_lo_lo_lo = {compressDataVec_selectReqData_97, compressDataVec_selectReqData_96};
  wire [15:0]   compressDataVec_hi_hi_lo_lo_lo_hi = {compressDataVec_selectReqData_99, compressDataVec_selectReqData_98};
  wire [31:0]   compressDataVec_hi_hi_lo_lo_lo = {compressDataVec_hi_hi_lo_lo_lo_hi, compressDataVec_hi_hi_lo_lo_lo_lo};
  wire [15:0]   compressDataVec_hi_hi_lo_lo_hi_lo = {compressDataVec_selectReqData_101, compressDataVec_selectReqData_100};
  wire [15:0]   compressDataVec_hi_hi_lo_lo_hi_hi = {compressDataVec_selectReqData_103, compressDataVec_selectReqData_102};
  wire [31:0]   compressDataVec_hi_hi_lo_lo_hi = {compressDataVec_hi_hi_lo_lo_hi_hi, compressDataVec_hi_hi_lo_lo_hi_lo};
  wire [63:0]   compressDataVec_hi_hi_lo_lo = {compressDataVec_hi_hi_lo_lo_hi, compressDataVec_hi_hi_lo_lo_lo};
  wire [15:0]   compressDataVec_hi_hi_lo_hi_lo_lo = {compressDataVec_selectReqData_105, compressDataVec_selectReqData_104};
  wire [15:0]   compressDataVec_hi_hi_lo_hi_lo_hi = {compressDataVec_selectReqData_107, compressDataVec_selectReqData_106};
  wire [31:0]   compressDataVec_hi_hi_lo_hi_lo = {compressDataVec_hi_hi_lo_hi_lo_hi, compressDataVec_hi_hi_lo_hi_lo_lo};
  wire [15:0]   compressDataVec_hi_hi_lo_hi_hi_lo = {compressDataVec_selectReqData_109, compressDataVec_selectReqData_108};
  wire [15:0]   compressDataVec_hi_hi_lo_hi_hi_hi = {compressDataVec_selectReqData_111, compressDataVec_selectReqData_110};
  wire [31:0]   compressDataVec_hi_hi_lo_hi_hi = {compressDataVec_hi_hi_lo_hi_hi_hi, compressDataVec_hi_hi_lo_hi_hi_lo};
  wire [63:0]   compressDataVec_hi_hi_lo_hi = {compressDataVec_hi_hi_lo_hi_hi, compressDataVec_hi_hi_lo_hi_lo};
  wire [127:0]  compressDataVec_hi_hi_lo = {compressDataVec_hi_hi_lo_hi, compressDataVec_hi_hi_lo_lo};
  wire [15:0]   compressDataVec_hi_hi_hi_lo_lo_lo = {compressDataVec_selectReqData_113, compressDataVec_selectReqData_112};
  wire [15:0]   compressDataVec_hi_hi_hi_lo_lo_hi = {compressDataVec_selectReqData_115, compressDataVec_selectReqData_114};
  wire [31:0]   compressDataVec_hi_hi_hi_lo_lo = {compressDataVec_hi_hi_hi_lo_lo_hi, compressDataVec_hi_hi_hi_lo_lo_lo};
  wire [15:0]   compressDataVec_hi_hi_hi_lo_hi_lo = {compressDataVec_selectReqData_117, compressDataVec_selectReqData_116};
  wire [15:0]   compressDataVec_hi_hi_hi_lo_hi_hi = {compressDataVec_selectReqData_119, compressDataVec_selectReqData_118};
  wire [31:0]   compressDataVec_hi_hi_hi_lo_hi = {compressDataVec_hi_hi_hi_lo_hi_hi, compressDataVec_hi_hi_hi_lo_hi_lo};
  wire [63:0]   compressDataVec_hi_hi_hi_lo = {compressDataVec_hi_hi_hi_lo_hi, compressDataVec_hi_hi_hi_lo_lo};
  wire [15:0]   compressDataVec_hi_hi_hi_hi_lo_lo = {compressDataVec_selectReqData_121, compressDataVec_selectReqData_120};
  wire [15:0]   compressDataVec_hi_hi_hi_hi_lo_hi = {compressDataVec_selectReqData_123, compressDataVec_selectReqData_122};
  wire [31:0]   compressDataVec_hi_hi_hi_hi_lo = {compressDataVec_hi_hi_hi_hi_lo_hi, compressDataVec_hi_hi_hi_hi_lo_lo};
  wire [15:0]   compressDataVec_hi_hi_hi_hi_hi_lo = {compressDataVec_selectReqData_125, compressDataVec_selectReqData_124};
  wire [15:0]   compressDataVec_hi_hi_hi_hi_hi_hi = {compressDataVec_selectReqData_127, compressDataVec_selectReqData_126};
  wire [31:0]   compressDataVec_hi_hi_hi_hi_hi = {compressDataVec_hi_hi_hi_hi_hi_hi, compressDataVec_hi_hi_hi_hi_hi_lo};
  wire [63:0]   compressDataVec_hi_hi_hi_hi = {compressDataVec_hi_hi_hi_hi_hi, compressDataVec_hi_hi_hi_hi_lo};
  wire [127:0]  compressDataVec_hi_hi_hi = {compressDataVec_hi_hi_hi_hi, compressDataVec_hi_hi_hi_lo};
  wire [255:0]  compressDataVec_hi_hi = {compressDataVec_hi_hi_hi, compressDataVec_hi_hi_lo};
  wire [511:0]  compressDataVec_hi = {compressDataVec_hi_hi, compressDataVec_hi_lo};
  wire [1023:0] compressDataVec_0 = {compressDataVec_hi, compressDataVec_lo};
  wire [15:0]   compressDataVec_selectReqData_128 =
    (compressDataVec_hitReq_0_128 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_128 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_128 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_128 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_128 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_128 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_128 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_128 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_128 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_128 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_128 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_128 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_128 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_128 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_128 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_128 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_128 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_128 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_128 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_128 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_128 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_128 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_128 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_128 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_128 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_128 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_128 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_128 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_128 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_128 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_128 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_128 ? source2Pipe[511:496] : 16'h0);
  wire          compressDataVec_useTail_64;
  assign compressDataVec_useTail_64 = |tailCount;
  wire [15:0]   compressDataVec_selectReqData_129 =
    (compressDataVec_hitReq_0_129 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_129 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_129 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_129 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_129 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_129 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_129 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_129 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_129 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_129 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_129 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_129 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_129 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_129 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_129 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_129 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_129 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_129 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_129 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_129 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_129 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_129 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_129 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_129 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_129 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_129 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_129 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_129 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_129 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_129 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_129 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_129 ? source2Pipe[511:496] : 16'h0);
  wire          compressDataVec_useTail_65;
  assign compressDataVec_useTail_65 = |(tailCount[5:1]);
  wire [15:0]   compressDataVec_selectReqData_130 =
    (compressDataVec_hitReq_0_130 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_130 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_130 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_130 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_130 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_130 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_130 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_130 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_130 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_130 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_130 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_130 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_130 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_130 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_130 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_130 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_130 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_130 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_130 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_130 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_130 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_130 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_130 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_130 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_130 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_130 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_130 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_130 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_130 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_130 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_130 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_130 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_131 =
    (compressDataVec_hitReq_0_131 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_131 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_131 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_131 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_131 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_131 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_131 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_131 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_131 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_131 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_131 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_131 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_131 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_131 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_131 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_131 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_131 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_131 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_131 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_131 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_131 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_131 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_131 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_131 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_131 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_131 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_131 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_131 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_131 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_131 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_131 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_131 ? source2Pipe[511:496] : 16'h0);
  wire          compressDataVec_useTail_67;
  assign compressDataVec_useTail_67 = |(tailCount[5:2]);
  wire [15:0]   compressDataVec_selectReqData_132 =
    (compressDataVec_hitReq_0_132 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_132 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_132 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_132 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_132 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_132 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_132 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_132 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_132 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_132 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_132 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_132 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_132 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_132 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_132 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_132 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_132 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_132 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_132 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_132 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_132 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_132 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_132 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_132 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_132 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_132 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_132 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_132 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_132 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_132 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_132 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_132 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_133 =
    (compressDataVec_hitReq_0_133 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_133 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_133 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_133 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_133 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_133 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_133 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_133 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_133 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_133 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_133 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_133 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_133 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_133 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_133 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_133 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_133 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_133 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_133 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_133 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_133 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_133 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_133 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_133 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_133 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_133 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_133 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_133 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_133 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_133 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_133 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_133 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_134 =
    (compressDataVec_hitReq_0_134 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_134 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_134 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_134 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_134 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_134 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_134 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_134 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_134 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_134 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_134 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_134 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_134 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_134 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_134 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_134 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_134 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_134 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_134 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_134 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_134 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_134 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_134 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_134 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_134 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_134 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_134 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_134 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_134 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_134 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_134 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_134 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_135 =
    (compressDataVec_hitReq_0_135 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_135 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_135 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_135 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_135 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_135 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_135 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_135 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_135 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_135 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_135 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_135 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_135 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_135 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_135 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_135 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_135 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_135 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_135 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_135 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_135 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_135 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_135 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_135 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_135 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_135 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_135 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_135 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_135 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_135 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_135 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_135 ? source2Pipe[511:496] : 16'h0);
  wire          compressDataVec_useTail_71;
  assign compressDataVec_useTail_71 = |(tailCount[5:3]);
  wire [15:0]   compressDataVec_selectReqData_136 =
    (compressDataVec_hitReq_0_136 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_136 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_136 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_136 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_136 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_136 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_136 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_136 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_136 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_136 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_136 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_136 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_136 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_136 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_136 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_136 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_136 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_136 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_136 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_136 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_136 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_136 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_136 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_136 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_136 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_136 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_136 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_136 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_136 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_136 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_136 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_136 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_137 =
    (compressDataVec_hitReq_0_137 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_137 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_137 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_137 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_137 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_137 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_137 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_137 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_137 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_137 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_137 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_137 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_137 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_137 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_137 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_137 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_137 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_137 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_137 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_137 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_137 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_137 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_137 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_137 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_137 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_137 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_137 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_137 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_137 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_137 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_137 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_137 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_138 =
    (compressDataVec_hitReq_0_138 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_138 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_138 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_138 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_138 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_138 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_138 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_138 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_138 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_138 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_138 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_138 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_138 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_138 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_138 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_138 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_138 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_138 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_138 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_138 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_138 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_138 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_138 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_138 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_138 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_138 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_138 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_138 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_138 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_138 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_138 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_138 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_139 =
    (compressDataVec_hitReq_0_139 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_139 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_139 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_139 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_139 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_139 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_139 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_139 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_139 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_139 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_139 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_139 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_139 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_139 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_139 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_139 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_139 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_139 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_139 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_139 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_139 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_139 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_139 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_139 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_139 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_139 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_139 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_139 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_139 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_139 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_139 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_139 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_140 =
    (compressDataVec_hitReq_0_140 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_140 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_140 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_140 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_140 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_140 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_140 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_140 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_140 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_140 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_140 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_140 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_140 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_140 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_140 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_140 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_140 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_140 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_140 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_140 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_140 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_140 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_140 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_140 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_140 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_140 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_140 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_140 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_140 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_140 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_140 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_140 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_141 =
    (compressDataVec_hitReq_0_141 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_141 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_141 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_141 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_141 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_141 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_141 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_141 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_141 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_141 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_141 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_141 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_141 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_141 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_141 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_141 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_141 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_141 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_141 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_141 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_141 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_141 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_141 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_141 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_141 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_141 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_141 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_141 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_141 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_141 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_141 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_141 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_142 =
    (compressDataVec_hitReq_0_142 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_142 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_142 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_142 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_142 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_142 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_142 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_142 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_142 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_142 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_142 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_142 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_142 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_142 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_142 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_142 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_142 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_142 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_142 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_142 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_142 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_142 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_142 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_142 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_142 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_142 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_142 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_142 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_142 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_142 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_142 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_142 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_143 =
    (compressDataVec_hitReq_0_143 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_143 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_143 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_143 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_143 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_143 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_143 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_143 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_143 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_143 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_143 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_143 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_143 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_143 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_143 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_143 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_143 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_143 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_143 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_143 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_143 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_143 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_143 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_143 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_143 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_143 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_143 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_143 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_143 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_143 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_143 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_143 ? source2Pipe[511:496] : 16'h0);
  wire          compressDataVec_useTail_79;
  assign compressDataVec_useTail_79 = |(tailCount[5:4]);
  wire [15:0]   compressDataVec_selectReqData_144 =
    (compressDataVec_hitReq_0_144 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_144 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_144 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_144 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_144 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_144 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_144 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_144 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_144 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_144 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_144 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_144 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_144 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_144 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_144 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_144 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_144 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_144 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_144 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_144 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_144 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_144 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_144 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_144 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_144 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_144 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_144 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_144 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_144 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_144 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_144 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_144 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_145 =
    (compressDataVec_hitReq_0_145 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_145 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_145 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_145 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_145 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_145 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_145 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_145 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_145 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_145 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_145 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_145 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_145 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_145 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_145 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_145 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_145 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_145 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_145 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_145 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_145 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_145 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_145 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_145 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_145 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_145 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_145 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_145 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_145 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_145 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_145 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_145 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_146 =
    (compressDataVec_hitReq_0_146 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_146 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_146 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_146 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_146 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_146 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_146 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_146 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_146 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_146 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_146 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_146 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_146 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_146 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_146 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_146 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_146 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_146 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_146 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_146 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_146 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_146 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_146 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_146 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_146 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_146 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_146 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_146 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_146 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_146 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_146 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_146 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_147 =
    (compressDataVec_hitReq_0_147 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_147 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_147 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_147 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_147 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_147 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_147 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_147 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_147 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_147 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_147 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_147 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_147 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_147 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_147 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_147 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_147 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_147 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_147 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_147 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_147 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_147 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_147 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_147 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_147 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_147 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_147 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_147 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_147 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_147 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_147 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_147 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_148 =
    (compressDataVec_hitReq_0_148 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_148 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_148 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_148 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_148 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_148 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_148 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_148 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_148 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_148 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_148 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_148 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_148 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_148 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_148 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_148 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_148 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_148 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_148 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_148 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_148 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_148 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_148 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_148 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_148 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_148 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_148 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_148 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_148 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_148 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_148 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_148 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_149 =
    (compressDataVec_hitReq_0_149 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_149 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_149 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_149 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_149 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_149 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_149 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_149 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_149 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_149 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_149 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_149 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_149 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_149 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_149 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_149 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_149 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_149 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_149 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_149 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_149 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_149 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_149 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_149 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_149 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_149 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_149 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_149 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_149 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_149 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_149 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_149 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_150 =
    (compressDataVec_hitReq_0_150 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_150 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_150 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_150 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_150 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_150 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_150 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_150 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_150 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_150 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_150 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_150 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_150 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_150 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_150 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_150 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_150 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_150 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_150 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_150 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_150 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_150 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_150 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_150 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_150 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_150 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_150 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_150 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_150 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_150 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_150 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_150 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_151 =
    (compressDataVec_hitReq_0_151 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_151 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_151 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_151 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_151 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_151 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_151 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_151 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_151 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_151 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_151 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_151 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_151 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_151 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_151 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_151 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_151 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_151 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_151 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_151 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_151 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_151 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_151 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_151 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_151 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_151 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_151 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_151 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_151 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_151 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_151 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_151 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_152 =
    (compressDataVec_hitReq_0_152 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_152 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_152 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_152 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_152 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_152 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_152 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_152 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_152 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_152 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_152 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_152 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_152 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_152 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_152 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_152 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_152 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_152 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_152 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_152 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_152 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_152 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_152 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_152 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_152 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_152 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_152 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_152 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_152 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_152 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_152 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_152 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_153 =
    (compressDataVec_hitReq_0_153 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_153 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_153 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_153 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_153 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_153 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_153 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_153 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_153 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_153 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_153 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_153 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_153 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_153 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_153 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_153 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_153 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_153 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_153 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_153 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_153 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_153 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_153 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_153 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_153 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_153 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_153 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_153 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_153 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_153 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_153 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_153 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_154 =
    (compressDataVec_hitReq_0_154 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_154 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_154 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_154 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_154 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_154 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_154 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_154 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_154 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_154 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_154 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_154 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_154 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_154 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_154 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_154 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_154 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_154 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_154 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_154 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_154 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_154 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_154 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_154 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_154 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_154 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_154 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_154 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_154 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_154 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_154 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_154 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_155 =
    (compressDataVec_hitReq_0_155 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_155 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_155 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_155 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_155 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_155 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_155 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_155 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_155 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_155 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_155 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_155 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_155 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_155 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_155 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_155 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_155 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_155 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_155 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_155 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_155 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_155 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_155 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_155 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_155 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_155 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_155 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_155 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_155 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_155 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_155 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_155 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_156 =
    (compressDataVec_hitReq_0_156 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_156 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_156 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_156 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_156 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_156 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_156 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_156 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_156 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_156 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_156 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_156 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_156 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_156 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_156 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_156 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_156 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_156 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_156 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_156 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_156 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_156 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_156 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_156 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_156 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_156 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_156 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_156 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_156 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_156 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_156 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_156 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_157 =
    (compressDataVec_hitReq_0_157 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_157 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_157 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_157 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_157 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_157 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_157 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_157 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_157 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_157 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_157 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_157 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_157 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_157 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_157 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_157 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_157 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_157 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_157 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_157 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_157 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_157 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_157 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_157 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_157 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_157 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_157 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_157 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_157 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_157 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_157 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_157 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_158 =
    (compressDataVec_hitReq_0_158 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_158 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_158 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_158 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_158 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_158 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_158 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_158 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_158 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_158 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_158 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_158 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_158 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_158 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_158 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_158 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_158 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_158 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_158 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_158 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_158 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_158 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_158 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_158 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_158 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_158 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_158 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_158 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_158 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_158 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_158 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_158 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_159 =
    (compressDataVec_hitReq_0_159 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_159 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_159 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_159 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_159 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_159 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_159 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_159 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_159 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_159 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_159 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_159 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_159 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_159 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_159 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_159 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_159 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_159 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_159 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_159 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_159 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_159 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_159 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_159 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_159 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_159 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_159 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_159 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_159 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_159 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_159 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_159 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_160 =
    (compressDataVec_hitReq_0_160 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_160 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_160 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_160 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_160 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_160 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_160 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_160 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_160 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_160 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_160 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_160 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_160 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_160 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_160 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_160 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_160 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_160 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_160 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_160 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_160 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_160 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_160 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_160 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_160 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_160 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_160 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_160 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_160 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_160 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_160 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_160 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_161 =
    (compressDataVec_hitReq_0_161 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_161 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_161 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_161 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_161 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_161 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_161 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_161 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_161 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_161 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_161 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_161 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_161 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_161 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_161 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_161 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_161 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_161 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_161 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_161 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_161 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_161 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_161 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_161 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_161 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_161 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_161 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_161 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_161 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_161 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_161 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_161 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_162 =
    (compressDataVec_hitReq_0_162 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_162 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_162 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_162 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_162 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_162 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_162 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_162 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_162 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_162 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_162 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_162 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_162 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_162 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_162 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_162 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_162 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_162 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_162 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_162 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_162 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_162 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_162 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_162 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_162 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_162 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_162 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_162 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_162 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_162 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_162 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_162 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_163 =
    (compressDataVec_hitReq_0_163 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_163 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_163 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_163 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_163 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_163 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_163 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_163 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_163 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_163 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_163 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_163 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_163 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_163 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_163 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_163 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_163 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_163 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_163 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_163 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_163 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_163 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_163 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_163 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_163 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_163 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_163 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_163 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_163 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_163 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_163 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_163 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_164 =
    (compressDataVec_hitReq_0_164 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_164 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_164 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_164 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_164 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_164 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_164 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_164 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_164 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_164 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_164 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_164 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_164 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_164 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_164 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_164 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_164 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_164 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_164 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_164 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_164 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_164 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_164 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_164 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_164 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_164 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_164 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_164 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_164 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_164 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_164 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_164 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_165 =
    (compressDataVec_hitReq_0_165 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_165 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_165 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_165 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_165 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_165 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_165 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_165 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_165 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_165 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_165 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_165 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_165 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_165 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_165 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_165 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_165 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_165 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_165 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_165 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_165 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_165 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_165 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_165 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_165 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_165 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_165 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_165 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_165 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_165 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_165 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_165 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_166 =
    (compressDataVec_hitReq_0_166 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_166 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_166 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_166 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_166 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_166 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_166 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_166 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_166 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_166 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_166 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_166 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_166 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_166 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_166 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_166 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_166 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_166 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_166 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_166 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_166 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_166 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_166 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_166 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_166 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_166 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_166 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_166 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_166 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_166 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_166 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_166 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_167 =
    (compressDataVec_hitReq_0_167 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_167 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_167 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_167 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_167 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_167 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_167 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_167 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_167 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_167 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_167 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_167 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_167 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_167 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_167 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_167 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_167 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_167 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_167 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_167 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_167 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_167 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_167 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_167 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_167 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_167 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_167 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_167 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_167 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_167 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_167 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_167 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_168 =
    (compressDataVec_hitReq_0_168 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_168 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_168 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_168 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_168 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_168 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_168 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_168 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_168 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_168 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_168 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_168 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_168 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_168 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_168 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_168 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_168 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_168 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_168 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_168 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_168 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_168 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_168 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_168 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_168 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_168 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_168 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_168 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_168 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_168 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_168 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_168 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_169 =
    (compressDataVec_hitReq_0_169 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_169 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_169 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_169 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_169 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_169 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_169 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_169 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_169 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_169 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_169 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_169 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_169 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_169 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_169 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_169 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_169 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_169 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_169 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_169 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_169 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_169 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_169 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_169 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_169 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_169 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_169 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_169 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_169 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_169 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_169 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_169 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_170 =
    (compressDataVec_hitReq_0_170 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_170 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_170 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_170 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_170 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_170 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_170 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_170 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_170 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_170 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_170 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_170 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_170 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_170 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_170 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_170 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_170 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_170 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_170 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_170 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_170 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_170 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_170 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_170 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_170 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_170 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_170 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_170 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_170 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_170 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_170 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_170 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_171 =
    (compressDataVec_hitReq_0_171 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_171 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_171 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_171 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_171 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_171 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_171 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_171 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_171 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_171 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_171 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_171 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_171 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_171 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_171 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_171 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_171 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_171 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_171 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_171 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_171 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_171 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_171 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_171 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_171 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_171 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_171 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_171 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_171 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_171 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_171 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_171 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_172 =
    (compressDataVec_hitReq_0_172 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_172 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_172 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_172 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_172 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_172 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_172 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_172 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_172 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_172 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_172 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_172 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_172 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_172 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_172 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_172 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_172 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_172 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_172 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_172 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_172 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_172 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_172 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_172 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_172 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_172 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_172 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_172 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_172 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_172 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_172 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_172 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_173 =
    (compressDataVec_hitReq_0_173 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_173 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_173 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_173 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_173 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_173 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_173 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_173 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_173 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_173 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_173 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_173 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_173 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_173 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_173 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_173 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_173 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_173 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_173 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_173 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_173 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_173 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_173 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_173 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_173 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_173 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_173 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_173 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_173 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_173 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_173 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_173 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_174 =
    (compressDataVec_hitReq_0_174 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_174 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_174 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_174 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_174 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_174 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_174 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_174 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_174 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_174 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_174 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_174 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_174 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_174 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_174 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_174 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_174 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_174 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_174 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_174 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_174 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_174 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_174 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_174 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_174 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_174 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_174 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_174 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_174 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_174 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_174 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_174 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_175 =
    (compressDataVec_hitReq_0_175 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_175 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_175 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_175 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_175 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_175 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_175 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_175 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_175 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_175 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_175 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_175 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_175 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_175 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_175 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_175 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_175 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_175 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_175 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_175 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_175 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_175 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_175 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_175 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_175 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_175 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_175 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_175 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_175 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_175 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_175 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_175 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_176 =
    (compressDataVec_hitReq_0_176 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_176 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_176 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_176 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_176 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_176 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_176 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_176 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_176 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_176 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_176 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_176 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_176 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_176 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_176 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_176 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_176 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_176 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_176 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_176 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_176 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_176 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_176 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_176 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_176 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_176 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_176 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_176 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_176 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_176 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_176 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_176 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_177 =
    (compressDataVec_hitReq_0_177 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_177 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_177 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_177 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_177 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_177 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_177 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_177 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_177 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_177 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_177 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_177 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_177 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_177 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_177 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_177 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_177 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_177 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_177 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_177 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_177 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_177 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_177 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_177 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_177 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_177 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_177 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_177 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_177 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_177 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_177 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_177 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_178 =
    (compressDataVec_hitReq_0_178 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_178 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_178 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_178 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_178 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_178 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_178 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_178 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_178 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_178 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_178 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_178 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_178 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_178 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_178 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_178 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_178 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_178 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_178 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_178 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_178 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_178 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_178 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_178 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_178 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_178 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_178 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_178 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_178 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_178 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_178 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_178 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_179 =
    (compressDataVec_hitReq_0_179 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_179 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_179 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_179 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_179 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_179 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_179 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_179 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_179 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_179 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_179 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_179 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_179 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_179 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_179 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_179 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_179 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_179 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_179 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_179 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_179 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_179 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_179 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_179 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_179 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_179 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_179 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_179 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_179 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_179 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_179 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_179 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_180 =
    (compressDataVec_hitReq_0_180 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_180 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_180 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_180 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_180 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_180 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_180 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_180 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_180 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_180 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_180 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_180 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_180 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_180 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_180 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_180 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_180 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_180 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_180 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_180 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_180 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_180 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_180 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_180 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_180 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_180 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_180 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_180 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_180 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_180 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_180 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_180 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_181 =
    (compressDataVec_hitReq_0_181 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_181 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_181 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_181 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_181 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_181 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_181 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_181 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_181 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_181 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_181 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_181 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_181 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_181 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_181 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_181 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_181 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_181 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_181 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_181 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_181 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_181 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_181 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_181 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_181 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_181 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_181 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_181 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_181 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_181 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_181 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_181 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_182 =
    (compressDataVec_hitReq_0_182 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_182 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_182 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_182 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_182 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_182 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_182 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_182 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_182 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_182 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_182 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_182 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_182 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_182 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_182 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_182 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_182 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_182 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_182 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_182 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_182 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_182 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_182 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_182 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_182 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_182 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_182 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_182 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_182 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_182 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_182 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_182 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_183 =
    (compressDataVec_hitReq_0_183 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_183 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_183 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_183 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_183 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_183 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_183 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_183 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_183 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_183 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_183 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_183 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_183 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_183 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_183 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_183 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_183 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_183 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_183 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_183 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_183 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_183 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_183 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_183 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_183 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_183 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_183 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_183 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_183 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_183 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_183 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_183 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_184 =
    (compressDataVec_hitReq_0_184 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_184 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_184 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_184 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_184 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_184 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_184 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_184 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_184 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_184 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_184 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_184 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_184 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_184 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_184 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_184 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_184 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_184 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_184 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_184 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_184 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_184 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_184 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_184 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_184 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_184 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_184 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_184 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_184 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_184 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_184 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_184 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_185 =
    (compressDataVec_hitReq_0_185 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_185 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_185 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_185 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_185 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_185 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_185 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_185 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_185 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_185 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_185 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_185 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_185 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_185 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_185 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_185 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_185 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_185 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_185 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_185 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_185 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_185 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_185 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_185 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_185 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_185 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_185 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_185 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_185 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_185 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_185 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_185 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_186 =
    (compressDataVec_hitReq_0_186 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_186 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_186 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_186 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_186 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_186 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_186 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_186 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_186 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_186 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_186 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_186 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_186 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_186 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_186 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_186 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_186 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_186 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_186 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_186 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_186 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_186 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_186 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_186 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_186 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_186 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_186 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_186 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_186 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_186 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_186 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_186 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_187 =
    (compressDataVec_hitReq_0_187 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_187 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_187 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_187 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_187 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_187 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_187 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_187 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_187 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_187 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_187 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_187 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_187 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_187 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_187 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_187 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_187 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_187 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_187 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_187 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_187 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_187 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_187 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_187 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_187 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_187 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_187 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_187 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_187 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_187 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_187 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_187 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_188 =
    (compressDataVec_hitReq_0_188 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_188 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_188 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_188 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_188 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_188 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_188 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_188 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_188 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_188 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_188 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_188 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_188 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_188 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_188 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_188 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_188 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_188 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_188 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_188 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_188 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_188 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_188 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_188 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_188 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_188 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_188 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_188 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_188 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_188 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_188 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_188 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_189 =
    (compressDataVec_hitReq_0_189 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_189 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_189 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_189 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_189 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_189 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_189 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_189 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_189 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_189 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_189 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_189 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_189 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_189 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_189 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_189 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_189 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_189 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_189 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_189 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_189 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_189 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_189 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_189 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_189 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_189 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_189 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_189 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_189 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_189 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_189 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_189 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_190 =
    (compressDataVec_hitReq_0_190 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_190 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_190 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_190 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_190 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_190 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_190 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_190 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_190 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_190 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_190 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_190 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_190 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_190 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_190 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_190 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_190 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_190 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_190 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_190 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_190 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_190 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_190 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_190 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_190 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_190 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_190 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_190 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_190 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_190 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_190 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_190 ? source2Pipe[511:496] : 16'h0);
  wire [15:0]   compressDataVec_selectReqData_191 =
    (compressDataVec_hitReq_0_191 ? source2Pipe[15:0] : 16'h0) | (compressDataVec_hitReq_1_191 ? source2Pipe[31:16] : 16'h0) | (compressDataVec_hitReq_2_191 ? source2Pipe[47:32] : 16'h0)
    | (compressDataVec_hitReq_3_191 ? source2Pipe[63:48] : 16'h0) | (compressDataVec_hitReq_4_191 ? source2Pipe[79:64] : 16'h0) | (compressDataVec_hitReq_5_191 ? source2Pipe[95:80] : 16'h0)
    | (compressDataVec_hitReq_6_191 ? source2Pipe[111:96] : 16'h0) | (compressDataVec_hitReq_7_191 ? source2Pipe[127:112] : 16'h0) | (compressDataVec_hitReq_8_191 ? source2Pipe[143:128] : 16'h0)
    | (compressDataVec_hitReq_9_191 ? source2Pipe[159:144] : 16'h0) | (compressDataVec_hitReq_10_191 ? source2Pipe[175:160] : 16'h0) | (compressDataVec_hitReq_11_191 ? source2Pipe[191:176] : 16'h0)
    | (compressDataVec_hitReq_12_191 ? source2Pipe[207:192] : 16'h0) | (compressDataVec_hitReq_13_191 ? source2Pipe[223:208] : 16'h0) | (compressDataVec_hitReq_14_191 ? source2Pipe[239:224] : 16'h0)
    | (compressDataVec_hitReq_15_191 ? source2Pipe[255:240] : 16'h0) | (compressDataVec_hitReq_16_191 ? source2Pipe[271:256] : 16'h0) | (compressDataVec_hitReq_17_191 ? source2Pipe[287:272] : 16'h0)
    | (compressDataVec_hitReq_18_191 ? source2Pipe[303:288] : 16'h0) | (compressDataVec_hitReq_19_191 ? source2Pipe[319:304] : 16'h0) | (compressDataVec_hitReq_20_191 ? source2Pipe[335:320] : 16'h0)
    | (compressDataVec_hitReq_21_191 ? source2Pipe[351:336] : 16'h0) | (compressDataVec_hitReq_22_191 ? source2Pipe[367:352] : 16'h0) | (compressDataVec_hitReq_23_191 ? source2Pipe[383:368] : 16'h0)
    | (compressDataVec_hitReq_24_191 ? source2Pipe[399:384] : 16'h0) | (compressDataVec_hitReq_25_191 ? source2Pipe[415:400] : 16'h0) | (compressDataVec_hitReq_26_191 ? source2Pipe[431:416] : 16'h0)
    | (compressDataVec_hitReq_27_191 ? source2Pipe[447:432] : 16'h0) | (compressDataVec_hitReq_28_191 ? source2Pipe[463:448] : 16'h0) | (compressDataVec_hitReq_29_191 ? source2Pipe[479:464] : 16'h0)
    | (compressDataVec_hitReq_30_191 ? source2Pipe[495:480] : 16'h0) | (compressDataVec_hitReq_31_191 ? source2Pipe[511:496] : 16'h0);
  wire [31:0]   compressDataVec_lo_lo_lo_lo_lo_1 = {compressDataVec_useTail_65 ? compressDataReg[31:16] : compressDataVec_selectReqData_129, compressDataVec_useTail_64 ? compressDataReg[15:0] : compressDataVec_selectReqData_128};
  wire [31:0]   compressDataVec_lo_lo_lo_lo_hi_1 = {compressDataVec_useTail_67 ? compressDataReg[63:48] : compressDataVec_selectReqData_131, compressDataVec_useTail_66 ? compressDataReg[47:32] : compressDataVec_selectReqData_130};
  wire [63:0]   compressDataVec_lo_lo_lo_lo_1 = {compressDataVec_lo_lo_lo_lo_hi_1, compressDataVec_lo_lo_lo_lo_lo_1};
  wire [31:0]   compressDataVec_lo_lo_lo_hi_lo_1 = {compressDataVec_useTail_69 ? compressDataReg[95:80] : compressDataVec_selectReqData_133, compressDataVec_useTail_68 ? compressDataReg[79:64] : compressDataVec_selectReqData_132};
  wire [31:0]   compressDataVec_lo_lo_lo_hi_hi_1 = {compressDataVec_useTail_71 ? compressDataReg[127:112] : compressDataVec_selectReqData_135, compressDataVec_useTail_70 ? compressDataReg[111:96] : compressDataVec_selectReqData_134};
  wire [63:0]   compressDataVec_lo_lo_lo_hi_1 = {compressDataVec_lo_lo_lo_hi_hi_1, compressDataVec_lo_lo_lo_hi_lo_1};
  wire [127:0]  compressDataVec_lo_lo_lo_1 = {compressDataVec_lo_lo_lo_hi_1, compressDataVec_lo_lo_lo_lo_1};
  wire [31:0]   compressDataVec_lo_lo_hi_lo_lo_1 = {compressDataVec_useTail_73 ? compressDataReg[159:144] : compressDataVec_selectReqData_137, compressDataVec_useTail_72 ? compressDataReg[143:128] : compressDataVec_selectReqData_136};
  wire [31:0]   compressDataVec_lo_lo_hi_lo_hi_1 = {compressDataVec_useTail_75 ? compressDataReg[191:176] : compressDataVec_selectReqData_139, compressDataVec_useTail_74 ? compressDataReg[175:160] : compressDataVec_selectReqData_138};
  wire [63:0]   compressDataVec_lo_lo_hi_lo_1 = {compressDataVec_lo_lo_hi_lo_hi_1, compressDataVec_lo_lo_hi_lo_lo_1};
  wire [31:0]   compressDataVec_lo_lo_hi_hi_lo_1 = {compressDataVec_useTail_77 ? compressDataReg[223:208] : compressDataVec_selectReqData_141, compressDataVec_useTail_76 ? compressDataReg[207:192] : compressDataVec_selectReqData_140};
  wire [31:0]   compressDataVec_lo_lo_hi_hi_hi_1 = {compressDataVec_useTail_79 ? compressDataReg[255:240] : compressDataVec_selectReqData_143, compressDataVec_useTail_78 ? compressDataReg[239:224] : compressDataVec_selectReqData_142};
  wire [63:0]   compressDataVec_lo_lo_hi_hi_1 = {compressDataVec_lo_lo_hi_hi_hi_1, compressDataVec_lo_lo_hi_hi_lo_1};
  wire [127:0]  compressDataVec_lo_lo_hi_1 = {compressDataVec_lo_lo_hi_hi_1, compressDataVec_lo_lo_hi_lo_1};
  wire [255:0]  compressDataVec_lo_lo_1 = {compressDataVec_lo_lo_hi_1, compressDataVec_lo_lo_lo_1};
  wire [31:0]   compressDataVec_lo_hi_lo_lo_lo_1 = {compressDataVec_useTail_81 ? compressDataReg[287:272] : compressDataVec_selectReqData_145, compressDataVec_useTail_80 ? compressDataReg[271:256] : compressDataVec_selectReqData_144};
  wire [31:0]   compressDataVec_lo_hi_lo_lo_hi_1 = {compressDataVec_useTail_83 ? compressDataReg[319:304] : compressDataVec_selectReqData_147, compressDataVec_useTail_82 ? compressDataReg[303:288] : compressDataVec_selectReqData_146};
  wire [63:0]   compressDataVec_lo_hi_lo_lo_1 = {compressDataVec_lo_hi_lo_lo_hi_1, compressDataVec_lo_hi_lo_lo_lo_1};
  wire [31:0]   compressDataVec_lo_hi_lo_hi_lo_1 = {compressDataVec_useTail_85 ? compressDataReg[351:336] : compressDataVec_selectReqData_149, compressDataVec_useTail_84 ? compressDataReg[335:320] : compressDataVec_selectReqData_148};
  wire [31:0]   compressDataVec_lo_hi_lo_hi_hi_1 = {compressDataVec_useTail_87 ? compressDataReg[383:368] : compressDataVec_selectReqData_151, compressDataVec_useTail_86 ? compressDataReg[367:352] : compressDataVec_selectReqData_150};
  wire [63:0]   compressDataVec_lo_hi_lo_hi_1 = {compressDataVec_lo_hi_lo_hi_hi_1, compressDataVec_lo_hi_lo_hi_lo_1};
  wire [127:0]  compressDataVec_lo_hi_lo_1 = {compressDataVec_lo_hi_lo_hi_1, compressDataVec_lo_hi_lo_lo_1};
  wire [31:0]   compressDataVec_lo_hi_hi_lo_lo_1 = {compressDataVec_useTail_89 ? compressDataReg[415:400] : compressDataVec_selectReqData_153, compressDataVec_useTail_88 ? compressDataReg[399:384] : compressDataVec_selectReqData_152};
  wire [31:0]   compressDataVec_lo_hi_hi_lo_hi_1 = {compressDataVec_useTail_91 ? compressDataReg[447:432] : compressDataVec_selectReqData_155, compressDataVec_useTail_90 ? compressDataReg[431:416] : compressDataVec_selectReqData_154};
  wire [63:0]   compressDataVec_lo_hi_hi_lo_1 = {compressDataVec_lo_hi_hi_lo_hi_1, compressDataVec_lo_hi_hi_lo_lo_1};
  wire [31:0]   compressDataVec_lo_hi_hi_hi_lo_1 = {compressDataVec_useTail_93 ? compressDataReg[479:464] : compressDataVec_selectReqData_157, compressDataVec_useTail_92 ? compressDataReg[463:448] : compressDataVec_selectReqData_156};
  wire [31:0]   compressDataVec_lo_hi_hi_hi_hi_1 = {compressDataVec_useTail_95 ? compressDataReg[511:496] : compressDataVec_selectReqData_159, compressDataVec_useTail_94 ? compressDataReg[495:480] : compressDataVec_selectReqData_158};
  wire [63:0]   compressDataVec_lo_hi_hi_hi_1 = {compressDataVec_lo_hi_hi_hi_hi_1, compressDataVec_lo_hi_hi_hi_lo_1};
  wire [127:0]  compressDataVec_lo_hi_hi_1 = {compressDataVec_lo_hi_hi_hi_1, compressDataVec_lo_hi_hi_lo_1};
  wire [255:0]  compressDataVec_lo_hi_1 = {compressDataVec_lo_hi_hi_1, compressDataVec_lo_hi_lo_1};
  wire [511:0]  compressDataVec_lo_1 = {compressDataVec_lo_hi_1, compressDataVec_lo_lo_1};
  wire [31:0]   compressDataVec_hi_lo_lo_lo_lo_1 = {compressDataVec_selectReqData_161, compressDataVec_selectReqData_160};
  wire [31:0]   compressDataVec_hi_lo_lo_lo_hi_1 = {compressDataVec_selectReqData_163, compressDataVec_selectReqData_162};
  wire [63:0]   compressDataVec_hi_lo_lo_lo_1 = {compressDataVec_hi_lo_lo_lo_hi_1, compressDataVec_hi_lo_lo_lo_lo_1};
  wire [31:0]   compressDataVec_hi_lo_lo_hi_lo_1 = {compressDataVec_selectReqData_165, compressDataVec_selectReqData_164};
  wire [31:0]   compressDataVec_hi_lo_lo_hi_hi_1 = {compressDataVec_selectReqData_167, compressDataVec_selectReqData_166};
  wire [63:0]   compressDataVec_hi_lo_lo_hi_1 = {compressDataVec_hi_lo_lo_hi_hi_1, compressDataVec_hi_lo_lo_hi_lo_1};
  wire [127:0]  compressDataVec_hi_lo_lo_1 = {compressDataVec_hi_lo_lo_hi_1, compressDataVec_hi_lo_lo_lo_1};
  wire [31:0]   compressDataVec_hi_lo_hi_lo_lo_1 = {compressDataVec_selectReqData_169, compressDataVec_selectReqData_168};
  wire [31:0]   compressDataVec_hi_lo_hi_lo_hi_1 = {compressDataVec_selectReqData_171, compressDataVec_selectReqData_170};
  wire [63:0]   compressDataVec_hi_lo_hi_lo_1 = {compressDataVec_hi_lo_hi_lo_hi_1, compressDataVec_hi_lo_hi_lo_lo_1};
  wire [31:0]   compressDataVec_hi_lo_hi_hi_lo_1 = {compressDataVec_selectReqData_173, compressDataVec_selectReqData_172};
  wire [31:0]   compressDataVec_hi_lo_hi_hi_hi_1 = {compressDataVec_selectReqData_175, compressDataVec_selectReqData_174};
  wire [63:0]   compressDataVec_hi_lo_hi_hi_1 = {compressDataVec_hi_lo_hi_hi_hi_1, compressDataVec_hi_lo_hi_hi_lo_1};
  wire [127:0]  compressDataVec_hi_lo_hi_1 = {compressDataVec_hi_lo_hi_hi_1, compressDataVec_hi_lo_hi_lo_1};
  wire [255:0]  compressDataVec_hi_lo_1 = {compressDataVec_hi_lo_hi_1, compressDataVec_hi_lo_lo_1};
  wire [31:0]   compressDataVec_hi_hi_lo_lo_lo_1 = {compressDataVec_selectReqData_177, compressDataVec_selectReqData_176};
  wire [31:0]   compressDataVec_hi_hi_lo_lo_hi_1 = {compressDataVec_selectReqData_179, compressDataVec_selectReqData_178};
  wire [63:0]   compressDataVec_hi_hi_lo_lo_1 = {compressDataVec_hi_hi_lo_lo_hi_1, compressDataVec_hi_hi_lo_lo_lo_1};
  wire [31:0]   compressDataVec_hi_hi_lo_hi_lo_1 = {compressDataVec_selectReqData_181, compressDataVec_selectReqData_180};
  wire [31:0]   compressDataVec_hi_hi_lo_hi_hi_1 = {compressDataVec_selectReqData_183, compressDataVec_selectReqData_182};
  wire [63:0]   compressDataVec_hi_hi_lo_hi_1 = {compressDataVec_hi_hi_lo_hi_hi_1, compressDataVec_hi_hi_lo_hi_lo_1};
  wire [127:0]  compressDataVec_hi_hi_lo_1 = {compressDataVec_hi_hi_lo_hi_1, compressDataVec_hi_hi_lo_lo_1};
  wire [31:0]   compressDataVec_hi_hi_hi_lo_lo_1 = {compressDataVec_selectReqData_185, compressDataVec_selectReqData_184};
  wire [31:0]   compressDataVec_hi_hi_hi_lo_hi_1 = {compressDataVec_selectReqData_187, compressDataVec_selectReqData_186};
  wire [63:0]   compressDataVec_hi_hi_hi_lo_1 = {compressDataVec_hi_hi_hi_lo_hi_1, compressDataVec_hi_hi_hi_lo_lo_1};
  wire [31:0]   compressDataVec_hi_hi_hi_hi_lo_1 = {compressDataVec_selectReqData_189, compressDataVec_selectReqData_188};
  wire [31:0]   compressDataVec_hi_hi_hi_hi_hi_1 = {compressDataVec_selectReqData_191, compressDataVec_selectReqData_190};
  wire [63:0]   compressDataVec_hi_hi_hi_hi_1 = {compressDataVec_hi_hi_hi_hi_hi_1, compressDataVec_hi_hi_hi_hi_lo_1};
  wire [127:0]  compressDataVec_hi_hi_hi_1 = {compressDataVec_hi_hi_hi_hi_1, compressDataVec_hi_hi_hi_lo_1};
  wire [255:0]  compressDataVec_hi_hi_1 = {compressDataVec_hi_hi_hi_1, compressDataVec_hi_hi_lo_1};
  wire [511:0]  compressDataVec_hi_1 = {compressDataVec_hi_hi_1, compressDataVec_hi_lo_1};
  wire [1023:0] compressDataVec_1 = {compressDataVec_hi_1, compressDataVec_lo_1};
  wire [31:0]   compressDataVec_selectReqData_192 =
    (compressDataVec_hitReq_0_192 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_192 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_192 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_192 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_192 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_192 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_192 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_192 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_192 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_192 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_192 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_192 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_192 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_192 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_192 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_192 ? source2Pipe[511:480] : 32'h0);
  wire          compressDataVec_useTail_96;
  assign compressDataVec_useTail_96 = |tailCount;
  wire [31:0]   compressDataVec_selectReqData_193 =
    (compressDataVec_hitReq_0_193 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_193 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_193 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_193 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_193 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_193 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_193 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_193 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_193 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_193 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_193 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_193 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_193 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_193 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_193 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_193 ? source2Pipe[511:480] : 32'h0);
  wire          compressDataVec_useTail_97;
  assign compressDataVec_useTail_97 = |(tailCount[5:1]);
  wire [31:0]   compressDataVec_selectReqData_194 =
    (compressDataVec_hitReq_0_194 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_194 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_194 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_194 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_194 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_194 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_194 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_194 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_194 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_194 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_194 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_194 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_194 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_194 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_194 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_194 ? source2Pipe[511:480] : 32'h0);
  wire [31:0]   compressDataVec_selectReqData_195 =
    (compressDataVec_hitReq_0_195 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_195 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_195 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_195 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_195 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_195 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_195 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_195 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_195 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_195 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_195 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_195 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_195 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_195 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_195 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_195 ? source2Pipe[511:480] : 32'h0);
  wire          compressDataVec_useTail_99;
  assign compressDataVec_useTail_99 = |(tailCount[5:2]);
  wire [31:0]   compressDataVec_selectReqData_196 =
    (compressDataVec_hitReq_0_196 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_196 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_196 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_196 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_196 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_196 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_196 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_196 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_196 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_196 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_196 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_196 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_196 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_196 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_196 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_196 ? source2Pipe[511:480] : 32'h0);
  wire [31:0]   compressDataVec_selectReqData_197 =
    (compressDataVec_hitReq_0_197 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_197 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_197 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_197 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_197 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_197 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_197 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_197 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_197 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_197 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_197 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_197 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_197 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_197 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_197 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_197 ? source2Pipe[511:480] : 32'h0);
  wire [31:0]   compressDataVec_selectReqData_198 =
    (compressDataVec_hitReq_0_198 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_198 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_198 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_198 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_198 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_198 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_198 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_198 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_198 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_198 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_198 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_198 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_198 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_198 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_198 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_198 ? source2Pipe[511:480] : 32'h0);
  wire [31:0]   compressDataVec_selectReqData_199 =
    (compressDataVec_hitReq_0_199 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_199 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_199 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_199 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_199 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_199 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_199 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_199 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_199 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_199 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_199 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_199 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_199 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_199 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_199 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_199 ? source2Pipe[511:480] : 32'h0);
  wire          compressDataVec_useTail_103;
  assign compressDataVec_useTail_103 = |(tailCount[5:3]);
  wire [31:0]   compressDataVec_selectReqData_200 =
    (compressDataVec_hitReq_0_200 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_200 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_200 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_200 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_200 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_200 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_200 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_200 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_200 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_200 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_200 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_200 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_200 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_200 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_200 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_200 ? source2Pipe[511:480] : 32'h0);
  wire [31:0]   compressDataVec_selectReqData_201 =
    (compressDataVec_hitReq_0_201 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_201 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_201 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_201 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_201 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_201 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_201 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_201 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_201 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_201 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_201 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_201 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_201 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_201 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_201 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_201 ? source2Pipe[511:480] : 32'h0);
  wire [31:0]   compressDataVec_selectReqData_202 =
    (compressDataVec_hitReq_0_202 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_202 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_202 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_202 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_202 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_202 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_202 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_202 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_202 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_202 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_202 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_202 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_202 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_202 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_202 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_202 ? source2Pipe[511:480] : 32'h0);
  wire [31:0]   compressDataVec_selectReqData_203 =
    (compressDataVec_hitReq_0_203 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_203 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_203 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_203 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_203 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_203 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_203 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_203 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_203 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_203 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_203 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_203 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_203 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_203 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_203 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_203 ? source2Pipe[511:480] : 32'h0);
  wire [31:0]   compressDataVec_selectReqData_204 =
    (compressDataVec_hitReq_0_204 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_204 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_204 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_204 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_204 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_204 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_204 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_204 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_204 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_204 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_204 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_204 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_204 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_204 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_204 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_204 ? source2Pipe[511:480] : 32'h0);
  wire [31:0]   compressDataVec_selectReqData_205 =
    (compressDataVec_hitReq_0_205 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_205 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_205 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_205 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_205 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_205 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_205 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_205 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_205 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_205 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_205 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_205 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_205 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_205 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_205 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_205 ? source2Pipe[511:480] : 32'h0);
  wire [31:0]   compressDataVec_selectReqData_206 =
    (compressDataVec_hitReq_0_206 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_206 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_206 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_206 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_206 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_206 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_206 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_206 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_206 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_206 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_206 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_206 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_206 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_206 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_206 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_206 ? source2Pipe[511:480] : 32'h0);
  wire [31:0]   compressDataVec_selectReqData_207 =
    (compressDataVec_hitReq_0_207 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_207 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_207 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_207 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_207 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_207 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_207 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_207 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_207 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_207 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_207 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_207 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_207 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_207 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_207 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_207 ? source2Pipe[511:480] : 32'h0);
  wire          compressDataVec_useTail_111;
  assign compressDataVec_useTail_111 = |(tailCount[5:4]);
  wire [31:0]   compressDataVec_selectReqData_208 =
    (compressDataVec_hitReq_0_208 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_208 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_208 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_208 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_208 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_208 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_208 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_208 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_208 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_208 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_208 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_208 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_208 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_208 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_208 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_208 ? source2Pipe[511:480] : 32'h0);
  wire [31:0]   compressDataVec_selectReqData_209 =
    (compressDataVec_hitReq_0_209 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_209 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_209 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_209 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_209 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_209 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_209 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_209 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_209 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_209 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_209 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_209 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_209 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_209 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_209 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_209 ? source2Pipe[511:480] : 32'h0);
  wire [31:0]   compressDataVec_selectReqData_210 =
    (compressDataVec_hitReq_0_210 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_210 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_210 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_210 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_210 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_210 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_210 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_210 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_210 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_210 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_210 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_210 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_210 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_210 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_210 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_210 ? source2Pipe[511:480] : 32'h0);
  wire [31:0]   compressDataVec_selectReqData_211 =
    (compressDataVec_hitReq_0_211 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_211 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_211 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_211 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_211 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_211 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_211 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_211 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_211 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_211 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_211 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_211 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_211 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_211 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_211 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_211 ? source2Pipe[511:480] : 32'h0);
  wire [31:0]   compressDataVec_selectReqData_212 =
    (compressDataVec_hitReq_0_212 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_212 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_212 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_212 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_212 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_212 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_212 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_212 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_212 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_212 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_212 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_212 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_212 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_212 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_212 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_212 ? source2Pipe[511:480] : 32'h0);
  wire [31:0]   compressDataVec_selectReqData_213 =
    (compressDataVec_hitReq_0_213 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_213 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_213 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_213 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_213 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_213 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_213 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_213 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_213 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_213 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_213 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_213 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_213 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_213 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_213 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_213 ? source2Pipe[511:480] : 32'h0);
  wire [31:0]   compressDataVec_selectReqData_214 =
    (compressDataVec_hitReq_0_214 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_214 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_214 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_214 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_214 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_214 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_214 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_214 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_214 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_214 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_214 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_214 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_214 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_214 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_214 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_214 ? source2Pipe[511:480] : 32'h0);
  wire [31:0]   compressDataVec_selectReqData_215 =
    (compressDataVec_hitReq_0_215 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_215 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_215 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_215 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_215 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_215 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_215 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_215 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_215 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_215 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_215 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_215 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_215 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_215 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_215 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_215 ? source2Pipe[511:480] : 32'h0);
  wire [31:0]   compressDataVec_selectReqData_216 =
    (compressDataVec_hitReq_0_216 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_216 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_216 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_216 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_216 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_216 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_216 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_216 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_216 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_216 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_216 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_216 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_216 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_216 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_216 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_216 ? source2Pipe[511:480] : 32'h0);
  wire [31:0]   compressDataVec_selectReqData_217 =
    (compressDataVec_hitReq_0_217 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_217 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_217 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_217 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_217 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_217 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_217 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_217 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_217 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_217 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_217 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_217 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_217 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_217 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_217 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_217 ? source2Pipe[511:480] : 32'h0);
  wire [31:0]   compressDataVec_selectReqData_218 =
    (compressDataVec_hitReq_0_218 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_218 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_218 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_218 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_218 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_218 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_218 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_218 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_218 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_218 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_218 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_218 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_218 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_218 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_218 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_218 ? source2Pipe[511:480] : 32'h0);
  wire [31:0]   compressDataVec_selectReqData_219 =
    (compressDataVec_hitReq_0_219 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_219 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_219 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_219 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_219 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_219 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_219 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_219 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_219 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_219 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_219 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_219 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_219 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_219 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_219 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_219 ? source2Pipe[511:480] : 32'h0);
  wire [31:0]   compressDataVec_selectReqData_220 =
    (compressDataVec_hitReq_0_220 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_220 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_220 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_220 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_220 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_220 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_220 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_220 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_220 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_220 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_220 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_220 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_220 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_220 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_220 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_220 ? source2Pipe[511:480] : 32'h0);
  wire [31:0]   compressDataVec_selectReqData_221 =
    (compressDataVec_hitReq_0_221 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_221 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_221 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_221 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_221 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_221 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_221 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_221 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_221 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_221 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_221 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_221 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_221 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_221 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_221 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_221 ? source2Pipe[511:480] : 32'h0);
  wire [31:0]   compressDataVec_selectReqData_222 =
    (compressDataVec_hitReq_0_222 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_222 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_222 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_222 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_222 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_222 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_222 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_222 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_222 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_222 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_222 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_222 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_222 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_222 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_222 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_222 ? source2Pipe[511:480] : 32'h0);
  wire [31:0]   compressDataVec_selectReqData_223 =
    (compressDataVec_hitReq_0_223 ? source2Pipe[31:0] : 32'h0) | (compressDataVec_hitReq_1_223 ? source2Pipe[63:32] : 32'h0) | (compressDataVec_hitReq_2_223 ? source2Pipe[95:64] : 32'h0)
    | (compressDataVec_hitReq_3_223 ? source2Pipe[127:96] : 32'h0) | (compressDataVec_hitReq_4_223 ? source2Pipe[159:128] : 32'h0) | (compressDataVec_hitReq_5_223 ? source2Pipe[191:160] : 32'h0)
    | (compressDataVec_hitReq_6_223 ? source2Pipe[223:192] : 32'h0) | (compressDataVec_hitReq_7_223 ? source2Pipe[255:224] : 32'h0) | (compressDataVec_hitReq_8_223 ? source2Pipe[287:256] : 32'h0)
    | (compressDataVec_hitReq_9_223 ? source2Pipe[319:288] : 32'h0) | (compressDataVec_hitReq_10_223 ? source2Pipe[351:320] : 32'h0) | (compressDataVec_hitReq_11_223 ? source2Pipe[383:352] : 32'h0)
    | (compressDataVec_hitReq_12_223 ? source2Pipe[415:384] : 32'h0) | (compressDataVec_hitReq_13_223 ? source2Pipe[447:416] : 32'h0) | (compressDataVec_hitReq_14_223 ? source2Pipe[479:448] : 32'h0)
    | (compressDataVec_hitReq_15_223 ? source2Pipe[511:480] : 32'h0);
  wire [63:0]   compressDataVec_lo_lo_lo_lo_2 = {compressDataVec_useTail_97 ? compressDataReg[63:32] : compressDataVec_selectReqData_193, compressDataVec_useTail_96 ? compressDataReg[31:0] : compressDataVec_selectReqData_192};
  wire [63:0]   compressDataVec_lo_lo_lo_hi_2 = {compressDataVec_useTail_99 ? compressDataReg[127:96] : compressDataVec_selectReqData_195, compressDataVec_useTail_98 ? compressDataReg[95:64] : compressDataVec_selectReqData_194};
  wire [127:0]  compressDataVec_lo_lo_lo_2 = {compressDataVec_lo_lo_lo_hi_2, compressDataVec_lo_lo_lo_lo_2};
  wire [63:0]   compressDataVec_lo_lo_hi_lo_2 = {compressDataVec_useTail_101 ? compressDataReg[191:160] : compressDataVec_selectReqData_197, compressDataVec_useTail_100 ? compressDataReg[159:128] : compressDataVec_selectReqData_196};
  wire [63:0]   compressDataVec_lo_lo_hi_hi_2 = {compressDataVec_useTail_103 ? compressDataReg[255:224] : compressDataVec_selectReqData_199, compressDataVec_useTail_102 ? compressDataReg[223:192] : compressDataVec_selectReqData_198};
  wire [127:0]  compressDataVec_lo_lo_hi_2 = {compressDataVec_lo_lo_hi_hi_2, compressDataVec_lo_lo_hi_lo_2};
  wire [255:0]  compressDataVec_lo_lo_2 = {compressDataVec_lo_lo_hi_2, compressDataVec_lo_lo_lo_2};
  wire [63:0]   compressDataVec_lo_hi_lo_lo_2 = {compressDataVec_useTail_105 ? compressDataReg[319:288] : compressDataVec_selectReqData_201, compressDataVec_useTail_104 ? compressDataReg[287:256] : compressDataVec_selectReqData_200};
  wire [63:0]   compressDataVec_lo_hi_lo_hi_2 = {compressDataVec_useTail_107 ? compressDataReg[383:352] : compressDataVec_selectReqData_203, compressDataVec_useTail_106 ? compressDataReg[351:320] : compressDataVec_selectReqData_202};
  wire [127:0]  compressDataVec_lo_hi_lo_2 = {compressDataVec_lo_hi_lo_hi_2, compressDataVec_lo_hi_lo_lo_2};
  wire [63:0]   compressDataVec_lo_hi_hi_lo_2 = {compressDataVec_useTail_109 ? compressDataReg[447:416] : compressDataVec_selectReqData_205, compressDataVec_useTail_108 ? compressDataReg[415:384] : compressDataVec_selectReqData_204};
  wire [63:0]   compressDataVec_lo_hi_hi_hi_2 = {compressDataVec_useTail_111 ? compressDataReg[511:480] : compressDataVec_selectReqData_207, compressDataVec_useTail_110 ? compressDataReg[479:448] : compressDataVec_selectReqData_206};
  wire [127:0]  compressDataVec_lo_hi_hi_2 = {compressDataVec_lo_hi_hi_hi_2, compressDataVec_lo_hi_hi_lo_2};
  wire [255:0]  compressDataVec_lo_hi_2 = {compressDataVec_lo_hi_hi_2, compressDataVec_lo_hi_lo_2};
  wire [511:0]  compressDataVec_lo_2 = {compressDataVec_lo_hi_2, compressDataVec_lo_lo_2};
  wire [63:0]   compressDataVec_hi_lo_lo_lo_2 = {compressDataVec_selectReqData_209, compressDataVec_selectReqData_208};
  wire [63:0]   compressDataVec_hi_lo_lo_hi_2 = {compressDataVec_selectReqData_211, compressDataVec_selectReqData_210};
  wire [127:0]  compressDataVec_hi_lo_lo_2 = {compressDataVec_hi_lo_lo_hi_2, compressDataVec_hi_lo_lo_lo_2};
  wire [63:0]   compressDataVec_hi_lo_hi_lo_2 = {compressDataVec_selectReqData_213, compressDataVec_selectReqData_212};
  wire [63:0]   compressDataVec_hi_lo_hi_hi_2 = {compressDataVec_selectReqData_215, compressDataVec_selectReqData_214};
  wire [127:0]  compressDataVec_hi_lo_hi_2 = {compressDataVec_hi_lo_hi_hi_2, compressDataVec_hi_lo_hi_lo_2};
  wire [255:0]  compressDataVec_hi_lo_2 = {compressDataVec_hi_lo_hi_2, compressDataVec_hi_lo_lo_2};
  wire [63:0]   compressDataVec_hi_hi_lo_lo_2 = {compressDataVec_selectReqData_217, compressDataVec_selectReqData_216};
  wire [63:0]   compressDataVec_hi_hi_lo_hi_2 = {compressDataVec_selectReqData_219, compressDataVec_selectReqData_218};
  wire [127:0]  compressDataVec_hi_hi_lo_2 = {compressDataVec_hi_hi_lo_hi_2, compressDataVec_hi_hi_lo_lo_2};
  wire [63:0]   compressDataVec_hi_hi_hi_lo_2 = {compressDataVec_selectReqData_221, compressDataVec_selectReqData_220};
  wire [63:0]   compressDataVec_hi_hi_hi_hi_2 = {compressDataVec_selectReqData_223, compressDataVec_selectReqData_222};
  wire [127:0]  compressDataVec_hi_hi_hi_2 = {compressDataVec_hi_hi_hi_hi_2, compressDataVec_hi_hi_hi_lo_2};
  wire [255:0]  compressDataVec_hi_hi_2 = {compressDataVec_hi_hi_hi_2, compressDataVec_hi_hi_lo_2};
  wire [511:0]  compressDataVec_hi_2 = {compressDataVec_hi_hi_2, compressDataVec_hi_lo_2};
  wire [1023:0] compressDataVec_2 = {compressDataVec_hi_2, compressDataVec_lo_2};
  wire [1023:0] compressResult = (eew1H[0] ? compressDataVec_0 : 1024'h0) | (eew1H[1] ? compressDataVec_1 : 1024'h0) | (eew1H[2] ? compressDataVec_2 : 1024'h0);
  wire          lastCompressEnq = stage2Valid & lastCompressPipe;
  wire [511:0]  splitCompressResult_0 = compressResult[511:0];
  wire [511:0]  splitCompressResult_1 = compressResult[1023:512];
  wire          compressTailMask_elementValid;
  assign compressTailMask_elementValid = |tailCountForMask;
  wire          compressTailMask_elementValid_1;
  assign compressTailMask_elementValid_1 = |(tailCountForMask[5:1]);
  wire          _GEN_2074 = tailCountForMask > 6'h2;
  wire          compressTailMask_elementValid_2;
  assign compressTailMask_elementValid_2 = _GEN_2074;
  wire          compressTailMask_elementValid_66;
  assign compressTailMask_elementValid_66 = _GEN_2074;
  wire          compressTailMask_elementValid_98;
  assign compressTailMask_elementValid_98 = _GEN_2074;
  wire          compressTailMask_elementValid_3;
  assign compressTailMask_elementValid_3 = |(tailCountForMask[5:2]);
  wire          _GEN_2075 = tailCountForMask > 6'h4;
  wire          compressTailMask_elementValid_4;
  assign compressTailMask_elementValid_4 = _GEN_2075;
  wire          compressTailMask_elementValid_68;
  assign compressTailMask_elementValid_68 = _GEN_2075;
  wire          compressTailMask_elementValid_100;
  assign compressTailMask_elementValid_100 = _GEN_2075;
  wire          _GEN_2076 = tailCountForMask > 6'h5;
  wire          compressTailMask_elementValid_5;
  assign compressTailMask_elementValid_5 = _GEN_2076;
  wire          compressTailMask_elementValid_69;
  assign compressTailMask_elementValid_69 = _GEN_2076;
  wire          compressTailMask_elementValid_101;
  assign compressTailMask_elementValid_101 = _GEN_2076;
  wire          _GEN_2077 = tailCountForMask > 6'h6;
  wire          compressTailMask_elementValid_6;
  assign compressTailMask_elementValid_6 = _GEN_2077;
  wire          compressTailMask_elementValid_70;
  assign compressTailMask_elementValid_70 = _GEN_2077;
  wire          compressTailMask_elementValid_102;
  assign compressTailMask_elementValid_102 = _GEN_2077;
  wire          compressTailMask_elementValid_7;
  assign compressTailMask_elementValid_7 = |(tailCountForMask[5:3]);
  wire          _GEN_2078 = tailCountForMask > 6'h8;
  wire          compressTailMask_elementValid_8;
  assign compressTailMask_elementValid_8 = _GEN_2078;
  wire          compressTailMask_elementValid_72;
  assign compressTailMask_elementValid_72 = _GEN_2078;
  wire          compressTailMask_elementValid_104;
  assign compressTailMask_elementValid_104 = _GEN_2078;
  wire          _GEN_2079 = tailCountForMask > 6'h9;
  wire          compressTailMask_elementValid_9;
  assign compressTailMask_elementValid_9 = _GEN_2079;
  wire          compressTailMask_elementValid_73;
  assign compressTailMask_elementValid_73 = _GEN_2079;
  wire          compressTailMask_elementValid_105;
  assign compressTailMask_elementValid_105 = _GEN_2079;
  wire          _GEN_2080 = tailCountForMask > 6'hA;
  wire          compressTailMask_elementValid_10;
  assign compressTailMask_elementValid_10 = _GEN_2080;
  wire          compressTailMask_elementValid_74;
  assign compressTailMask_elementValid_74 = _GEN_2080;
  wire          compressTailMask_elementValid_106;
  assign compressTailMask_elementValid_106 = _GEN_2080;
  wire          _GEN_2081 = tailCountForMask > 6'hB;
  wire          compressTailMask_elementValid_11;
  assign compressTailMask_elementValid_11 = _GEN_2081;
  wire          compressTailMask_elementValid_75;
  assign compressTailMask_elementValid_75 = _GEN_2081;
  wire          compressTailMask_elementValid_107;
  assign compressTailMask_elementValid_107 = _GEN_2081;
  wire          _GEN_2082 = tailCountForMask > 6'hC;
  wire          compressTailMask_elementValid_12;
  assign compressTailMask_elementValid_12 = _GEN_2082;
  wire          compressTailMask_elementValid_76;
  assign compressTailMask_elementValid_76 = _GEN_2082;
  wire          compressTailMask_elementValid_108;
  assign compressTailMask_elementValid_108 = _GEN_2082;
  wire          _GEN_2083 = tailCountForMask > 6'hD;
  wire          compressTailMask_elementValid_13;
  assign compressTailMask_elementValid_13 = _GEN_2083;
  wire          compressTailMask_elementValid_77;
  assign compressTailMask_elementValid_77 = _GEN_2083;
  wire          compressTailMask_elementValid_109;
  assign compressTailMask_elementValid_109 = _GEN_2083;
  wire          _GEN_2084 = tailCountForMask > 6'hE;
  wire          compressTailMask_elementValid_14;
  assign compressTailMask_elementValid_14 = _GEN_2084;
  wire          compressTailMask_elementValid_78;
  assign compressTailMask_elementValid_78 = _GEN_2084;
  wire          compressTailMask_elementValid_110;
  assign compressTailMask_elementValid_110 = _GEN_2084;
  wire          compressTailMask_elementValid_15;
  assign compressTailMask_elementValid_15 = |(tailCountForMask[5:4]);
  wire          _GEN_2085 = tailCountForMask > 6'h10;
  wire          compressTailMask_elementValid_16;
  assign compressTailMask_elementValid_16 = _GEN_2085;
  wire          compressTailMask_elementValid_80;
  assign compressTailMask_elementValid_80 = _GEN_2085;
  wire          _GEN_2086 = tailCountForMask > 6'h11;
  wire          compressTailMask_elementValid_17;
  assign compressTailMask_elementValid_17 = _GEN_2086;
  wire          compressTailMask_elementValid_81;
  assign compressTailMask_elementValid_81 = _GEN_2086;
  wire          _GEN_2087 = tailCountForMask > 6'h12;
  wire          compressTailMask_elementValid_18;
  assign compressTailMask_elementValid_18 = _GEN_2087;
  wire          compressTailMask_elementValid_82;
  assign compressTailMask_elementValid_82 = _GEN_2087;
  wire          _GEN_2088 = tailCountForMask > 6'h13;
  wire          compressTailMask_elementValid_19;
  assign compressTailMask_elementValid_19 = _GEN_2088;
  wire          compressTailMask_elementValid_83;
  assign compressTailMask_elementValid_83 = _GEN_2088;
  wire          _GEN_2089 = tailCountForMask > 6'h14;
  wire          compressTailMask_elementValid_20;
  assign compressTailMask_elementValid_20 = _GEN_2089;
  wire          compressTailMask_elementValid_84;
  assign compressTailMask_elementValid_84 = _GEN_2089;
  wire          _GEN_2090 = tailCountForMask > 6'h15;
  wire          compressTailMask_elementValid_21;
  assign compressTailMask_elementValid_21 = _GEN_2090;
  wire          compressTailMask_elementValid_85;
  assign compressTailMask_elementValid_85 = _GEN_2090;
  wire          _GEN_2091 = tailCountForMask > 6'h16;
  wire          compressTailMask_elementValid_22;
  assign compressTailMask_elementValid_22 = _GEN_2091;
  wire          compressTailMask_elementValid_86;
  assign compressTailMask_elementValid_86 = _GEN_2091;
  wire          _GEN_2092 = tailCountForMask > 6'h17;
  wire          compressTailMask_elementValid_23;
  assign compressTailMask_elementValid_23 = _GEN_2092;
  wire          compressTailMask_elementValid_87;
  assign compressTailMask_elementValid_87 = _GEN_2092;
  wire          _GEN_2093 = tailCountForMask > 6'h18;
  wire          compressTailMask_elementValid_24;
  assign compressTailMask_elementValid_24 = _GEN_2093;
  wire          compressTailMask_elementValid_88;
  assign compressTailMask_elementValid_88 = _GEN_2093;
  wire          _GEN_2094 = tailCountForMask > 6'h19;
  wire          compressTailMask_elementValid_25;
  assign compressTailMask_elementValid_25 = _GEN_2094;
  wire          compressTailMask_elementValid_89;
  assign compressTailMask_elementValid_89 = _GEN_2094;
  wire          _GEN_2095 = tailCountForMask > 6'h1A;
  wire          compressTailMask_elementValid_26;
  assign compressTailMask_elementValid_26 = _GEN_2095;
  wire          compressTailMask_elementValid_90;
  assign compressTailMask_elementValid_90 = _GEN_2095;
  wire          _GEN_2096 = tailCountForMask > 6'h1B;
  wire          compressTailMask_elementValid_27;
  assign compressTailMask_elementValid_27 = _GEN_2096;
  wire          compressTailMask_elementValid_91;
  assign compressTailMask_elementValid_91 = _GEN_2096;
  wire          _GEN_2097 = tailCountForMask > 6'h1C;
  wire          compressTailMask_elementValid_28;
  assign compressTailMask_elementValid_28 = _GEN_2097;
  wire          compressTailMask_elementValid_92;
  assign compressTailMask_elementValid_92 = _GEN_2097;
  wire          _GEN_2098 = tailCountForMask > 6'h1D;
  wire          compressTailMask_elementValid_29;
  assign compressTailMask_elementValid_29 = _GEN_2098;
  wire          compressTailMask_elementValid_93;
  assign compressTailMask_elementValid_93 = _GEN_2098;
  wire          _GEN_2099 = tailCountForMask > 6'h1E;
  wire          compressTailMask_elementValid_30;
  assign compressTailMask_elementValid_30 = _GEN_2099;
  wire          compressTailMask_elementValid_94;
  assign compressTailMask_elementValid_94 = _GEN_2099;
  wire          compressTailMask_elementValid_31 = tailCountForMask[5];
  wire          compressTailMask_elementValid_95 = tailCountForMask[5];
  wire          compressTailMask_elementValid_32 = tailCountForMask > 6'h20;
  wire          compressTailMask_elementValid_33 = tailCountForMask > 6'h21;
  wire          compressTailMask_elementValid_34 = tailCountForMask > 6'h22;
  wire          compressTailMask_elementValid_35 = tailCountForMask > 6'h23;
  wire          compressTailMask_elementValid_36 = tailCountForMask > 6'h24;
  wire          compressTailMask_elementValid_37 = tailCountForMask > 6'h25;
  wire          compressTailMask_elementValid_38 = tailCountForMask > 6'h26;
  wire          compressTailMask_elementValid_39 = tailCountForMask > 6'h27;
  wire          compressTailMask_elementValid_40 = tailCountForMask > 6'h28;
  wire          compressTailMask_elementValid_41 = tailCountForMask > 6'h29;
  wire          compressTailMask_elementValid_42 = tailCountForMask > 6'h2A;
  wire          compressTailMask_elementValid_43 = tailCountForMask > 6'h2B;
  wire          compressTailMask_elementValid_44 = tailCountForMask > 6'h2C;
  wire          compressTailMask_elementValid_45 = tailCountForMask > 6'h2D;
  wire          compressTailMask_elementValid_46 = tailCountForMask > 6'h2E;
  wire          compressTailMask_elementValid_47 = tailCountForMask > 6'h2F;
  wire          compressTailMask_elementValid_48 = tailCountForMask > 6'h30;
  wire          compressTailMask_elementValid_49 = tailCountForMask > 6'h31;
  wire          compressTailMask_elementValid_50 = tailCountForMask > 6'h32;
  wire          compressTailMask_elementValid_51 = tailCountForMask > 6'h33;
  wire          compressTailMask_elementValid_52 = tailCountForMask > 6'h34;
  wire          compressTailMask_elementValid_53 = tailCountForMask > 6'h35;
  wire          compressTailMask_elementValid_54 = tailCountForMask > 6'h36;
  wire          compressTailMask_elementValid_55 = tailCountForMask > 6'h37;
  wire          compressTailMask_elementValid_56 = tailCountForMask > 6'h38;
  wire          compressTailMask_elementValid_57 = tailCountForMask > 6'h39;
  wire          compressTailMask_elementValid_58 = tailCountForMask > 6'h3A;
  wire          compressTailMask_elementValid_59 = tailCountForMask > 6'h3B;
  wire          compressTailMask_elementValid_60 = tailCountForMask > 6'h3C;
  wire          compressTailMask_elementValid_61 = tailCountForMask > 6'h3D;
  wire          compressTailMask_elementValid_62 = &tailCountForMask;
  wire [1:0]    compressTailMask_lo_lo_lo_lo_lo = {compressTailMask_elementValid_1, compressTailMask_elementValid};
  wire [1:0]    compressTailMask_lo_lo_lo_lo_hi = {compressTailMask_elementValid_3, compressTailMask_elementValid_2};
  wire [3:0]    compressTailMask_lo_lo_lo_lo = {compressTailMask_lo_lo_lo_lo_hi, compressTailMask_lo_lo_lo_lo_lo};
  wire [1:0]    compressTailMask_lo_lo_lo_hi_lo = {compressTailMask_elementValid_5, compressTailMask_elementValid_4};
  wire [1:0]    compressTailMask_lo_lo_lo_hi_hi = {compressTailMask_elementValid_7, compressTailMask_elementValid_6};
  wire [3:0]    compressTailMask_lo_lo_lo_hi = {compressTailMask_lo_lo_lo_hi_hi, compressTailMask_lo_lo_lo_hi_lo};
  wire [7:0]    compressTailMask_lo_lo_lo = {compressTailMask_lo_lo_lo_hi, compressTailMask_lo_lo_lo_lo};
  wire [1:0]    compressTailMask_lo_lo_hi_lo_lo = {compressTailMask_elementValid_9, compressTailMask_elementValid_8};
  wire [1:0]    compressTailMask_lo_lo_hi_lo_hi = {compressTailMask_elementValid_11, compressTailMask_elementValid_10};
  wire [3:0]    compressTailMask_lo_lo_hi_lo = {compressTailMask_lo_lo_hi_lo_hi, compressTailMask_lo_lo_hi_lo_lo};
  wire [1:0]    compressTailMask_lo_lo_hi_hi_lo = {compressTailMask_elementValid_13, compressTailMask_elementValid_12};
  wire [1:0]    compressTailMask_lo_lo_hi_hi_hi = {compressTailMask_elementValid_15, compressTailMask_elementValid_14};
  wire [3:0]    compressTailMask_lo_lo_hi_hi = {compressTailMask_lo_lo_hi_hi_hi, compressTailMask_lo_lo_hi_hi_lo};
  wire [7:0]    compressTailMask_lo_lo_hi = {compressTailMask_lo_lo_hi_hi, compressTailMask_lo_lo_hi_lo};
  wire [15:0]   compressTailMask_lo_lo = {compressTailMask_lo_lo_hi, compressTailMask_lo_lo_lo};
  wire [1:0]    compressTailMask_lo_hi_lo_lo_lo = {compressTailMask_elementValid_17, compressTailMask_elementValid_16};
  wire [1:0]    compressTailMask_lo_hi_lo_lo_hi = {compressTailMask_elementValid_19, compressTailMask_elementValid_18};
  wire [3:0]    compressTailMask_lo_hi_lo_lo = {compressTailMask_lo_hi_lo_lo_hi, compressTailMask_lo_hi_lo_lo_lo};
  wire [1:0]    compressTailMask_lo_hi_lo_hi_lo = {compressTailMask_elementValid_21, compressTailMask_elementValid_20};
  wire [1:0]    compressTailMask_lo_hi_lo_hi_hi = {compressTailMask_elementValid_23, compressTailMask_elementValid_22};
  wire [3:0]    compressTailMask_lo_hi_lo_hi = {compressTailMask_lo_hi_lo_hi_hi, compressTailMask_lo_hi_lo_hi_lo};
  wire [7:0]    compressTailMask_lo_hi_lo = {compressTailMask_lo_hi_lo_hi, compressTailMask_lo_hi_lo_lo};
  wire [1:0]    compressTailMask_lo_hi_hi_lo_lo = {compressTailMask_elementValid_25, compressTailMask_elementValid_24};
  wire [1:0]    compressTailMask_lo_hi_hi_lo_hi = {compressTailMask_elementValid_27, compressTailMask_elementValid_26};
  wire [3:0]    compressTailMask_lo_hi_hi_lo = {compressTailMask_lo_hi_hi_lo_hi, compressTailMask_lo_hi_hi_lo_lo};
  wire [1:0]    compressTailMask_lo_hi_hi_hi_lo = {compressTailMask_elementValid_29, compressTailMask_elementValid_28};
  wire [1:0]    compressTailMask_lo_hi_hi_hi_hi = {compressTailMask_elementValid_31, compressTailMask_elementValid_30};
  wire [3:0]    compressTailMask_lo_hi_hi_hi = {compressTailMask_lo_hi_hi_hi_hi, compressTailMask_lo_hi_hi_hi_lo};
  wire [7:0]    compressTailMask_lo_hi_hi = {compressTailMask_lo_hi_hi_hi, compressTailMask_lo_hi_hi_lo};
  wire [15:0]   compressTailMask_lo_hi = {compressTailMask_lo_hi_hi, compressTailMask_lo_hi_lo};
  wire [31:0]   compressTailMask_lo = {compressTailMask_lo_hi, compressTailMask_lo_lo};
  wire [1:0]    compressTailMask_hi_lo_lo_lo_lo = {compressTailMask_elementValid_33, compressTailMask_elementValid_32};
  wire [1:0]    compressTailMask_hi_lo_lo_lo_hi = {compressTailMask_elementValid_35, compressTailMask_elementValid_34};
  wire [3:0]    compressTailMask_hi_lo_lo_lo = {compressTailMask_hi_lo_lo_lo_hi, compressTailMask_hi_lo_lo_lo_lo};
  wire [1:0]    compressTailMask_hi_lo_lo_hi_lo = {compressTailMask_elementValid_37, compressTailMask_elementValid_36};
  wire [1:0]    compressTailMask_hi_lo_lo_hi_hi = {compressTailMask_elementValid_39, compressTailMask_elementValid_38};
  wire [3:0]    compressTailMask_hi_lo_lo_hi = {compressTailMask_hi_lo_lo_hi_hi, compressTailMask_hi_lo_lo_hi_lo};
  wire [7:0]    compressTailMask_hi_lo_lo = {compressTailMask_hi_lo_lo_hi, compressTailMask_hi_lo_lo_lo};
  wire [1:0]    compressTailMask_hi_lo_hi_lo_lo = {compressTailMask_elementValid_41, compressTailMask_elementValid_40};
  wire [1:0]    compressTailMask_hi_lo_hi_lo_hi = {compressTailMask_elementValid_43, compressTailMask_elementValid_42};
  wire [3:0]    compressTailMask_hi_lo_hi_lo = {compressTailMask_hi_lo_hi_lo_hi, compressTailMask_hi_lo_hi_lo_lo};
  wire [1:0]    compressTailMask_hi_lo_hi_hi_lo = {compressTailMask_elementValid_45, compressTailMask_elementValid_44};
  wire [1:0]    compressTailMask_hi_lo_hi_hi_hi = {compressTailMask_elementValid_47, compressTailMask_elementValid_46};
  wire [3:0]    compressTailMask_hi_lo_hi_hi = {compressTailMask_hi_lo_hi_hi_hi, compressTailMask_hi_lo_hi_hi_lo};
  wire [7:0]    compressTailMask_hi_lo_hi = {compressTailMask_hi_lo_hi_hi, compressTailMask_hi_lo_hi_lo};
  wire [15:0]   compressTailMask_hi_lo = {compressTailMask_hi_lo_hi, compressTailMask_hi_lo_lo};
  wire [1:0]    compressTailMask_hi_hi_lo_lo_lo = {compressTailMask_elementValid_49, compressTailMask_elementValid_48};
  wire [1:0]    compressTailMask_hi_hi_lo_lo_hi = {compressTailMask_elementValid_51, compressTailMask_elementValid_50};
  wire [3:0]    compressTailMask_hi_hi_lo_lo = {compressTailMask_hi_hi_lo_lo_hi, compressTailMask_hi_hi_lo_lo_lo};
  wire [1:0]    compressTailMask_hi_hi_lo_hi_lo = {compressTailMask_elementValid_53, compressTailMask_elementValid_52};
  wire [1:0]    compressTailMask_hi_hi_lo_hi_hi = {compressTailMask_elementValid_55, compressTailMask_elementValid_54};
  wire [3:0]    compressTailMask_hi_hi_lo_hi = {compressTailMask_hi_hi_lo_hi_hi, compressTailMask_hi_hi_lo_hi_lo};
  wire [7:0]    compressTailMask_hi_hi_lo = {compressTailMask_hi_hi_lo_hi, compressTailMask_hi_hi_lo_lo};
  wire [1:0]    compressTailMask_hi_hi_hi_lo_lo = {compressTailMask_elementValid_57, compressTailMask_elementValid_56};
  wire [1:0]    compressTailMask_hi_hi_hi_lo_hi = {compressTailMask_elementValid_59, compressTailMask_elementValid_58};
  wire [3:0]    compressTailMask_hi_hi_hi_lo = {compressTailMask_hi_hi_hi_lo_hi, compressTailMask_hi_hi_hi_lo_lo};
  wire [1:0]    compressTailMask_hi_hi_hi_hi_lo = {compressTailMask_elementValid_61, compressTailMask_elementValid_60};
  wire [1:0]    compressTailMask_hi_hi_hi_hi_hi = {1'h0, compressTailMask_elementValid_62};
  wire [3:0]    compressTailMask_hi_hi_hi_hi = {compressTailMask_hi_hi_hi_hi_hi, compressTailMask_hi_hi_hi_hi_lo};
  wire [7:0]    compressTailMask_hi_hi_hi = {compressTailMask_hi_hi_hi_hi, compressTailMask_hi_hi_hi_lo};
  wire [15:0]   compressTailMask_hi_hi = {compressTailMask_hi_hi_hi, compressTailMask_hi_hi_lo};
  wire [31:0]   compressTailMask_hi = {compressTailMask_hi_hi, compressTailMask_hi_lo};
  wire          compressTailMask_elementValid_64;
  assign compressTailMask_elementValid_64 = |tailCountForMask;
  wire [1:0]    compressTailMask_elementMask = {2{compressTailMask_elementValid_64}};
  wire          compressTailMask_elementValid_65;
  assign compressTailMask_elementValid_65 = |(tailCountForMask[5:1]);
  wire [1:0]    compressTailMask_elementMask_1 = {2{compressTailMask_elementValid_65}};
  wire [1:0]    compressTailMask_elementMask_2 = {2{compressTailMask_elementValid_66}};
  wire          compressTailMask_elementValid_67;
  assign compressTailMask_elementValid_67 = |(tailCountForMask[5:2]);
  wire [1:0]    compressTailMask_elementMask_3 = {2{compressTailMask_elementValid_67}};
  wire [1:0]    compressTailMask_elementMask_4 = {2{compressTailMask_elementValid_68}};
  wire [1:0]    compressTailMask_elementMask_5 = {2{compressTailMask_elementValid_69}};
  wire [1:0]    compressTailMask_elementMask_6 = {2{compressTailMask_elementValid_70}};
  wire          compressTailMask_elementValid_71;
  assign compressTailMask_elementValid_71 = |(tailCountForMask[5:3]);
  wire [1:0]    compressTailMask_elementMask_7 = {2{compressTailMask_elementValid_71}};
  wire [1:0]    compressTailMask_elementMask_8 = {2{compressTailMask_elementValid_72}};
  wire [1:0]    compressTailMask_elementMask_9 = {2{compressTailMask_elementValid_73}};
  wire [1:0]    compressTailMask_elementMask_10 = {2{compressTailMask_elementValid_74}};
  wire [1:0]    compressTailMask_elementMask_11 = {2{compressTailMask_elementValid_75}};
  wire [1:0]    compressTailMask_elementMask_12 = {2{compressTailMask_elementValid_76}};
  wire [1:0]    compressTailMask_elementMask_13 = {2{compressTailMask_elementValid_77}};
  wire [1:0]    compressTailMask_elementMask_14 = {2{compressTailMask_elementValid_78}};
  wire          compressTailMask_elementValid_79;
  assign compressTailMask_elementValid_79 = |(tailCountForMask[5:4]);
  wire [1:0]    compressTailMask_elementMask_15 = {2{compressTailMask_elementValid_79}};
  wire [1:0]    compressTailMask_elementMask_16 = {2{compressTailMask_elementValid_80}};
  wire [1:0]    compressTailMask_elementMask_17 = {2{compressTailMask_elementValid_81}};
  wire [1:0]    compressTailMask_elementMask_18 = {2{compressTailMask_elementValid_82}};
  wire [1:0]    compressTailMask_elementMask_19 = {2{compressTailMask_elementValid_83}};
  wire [1:0]    compressTailMask_elementMask_20 = {2{compressTailMask_elementValid_84}};
  wire [1:0]    compressTailMask_elementMask_21 = {2{compressTailMask_elementValid_85}};
  wire [1:0]    compressTailMask_elementMask_22 = {2{compressTailMask_elementValid_86}};
  wire [1:0]    compressTailMask_elementMask_23 = {2{compressTailMask_elementValid_87}};
  wire [1:0]    compressTailMask_elementMask_24 = {2{compressTailMask_elementValid_88}};
  wire [1:0]    compressTailMask_elementMask_25 = {2{compressTailMask_elementValid_89}};
  wire [1:0]    compressTailMask_elementMask_26 = {2{compressTailMask_elementValid_90}};
  wire [1:0]    compressTailMask_elementMask_27 = {2{compressTailMask_elementValid_91}};
  wire [1:0]    compressTailMask_elementMask_28 = {2{compressTailMask_elementValid_92}};
  wire [1:0]    compressTailMask_elementMask_29 = {2{compressTailMask_elementValid_93}};
  wire [1:0]    compressTailMask_elementMask_30 = {2{compressTailMask_elementValid_94}};
  wire [1:0]    compressTailMask_elementMask_31 = {2{compressTailMask_elementValid_95}};
  wire [3:0]    compressTailMask_lo_lo_lo_lo_1 = {compressTailMask_elementMask_1, compressTailMask_elementMask};
  wire [3:0]    compressTailMask_lo_lo_lo_hi_1 = {compressTailMask_elementMask_3, compressTailMask_elementMask_2};
  wire [7:0]    compressTailMask_lo_lo_lo_1 = {compressTailMask_lo_lo_lo_hi_1, compressTailMask_lo_lo_lo_lo_1};
  wire [3:0]    compressTailMask_lo_lo_hi_lo_1 = {compressTailMask_elementMask_5, compressTailMask_elementMask_4};
  wire [3:0]    compressTailMask_lo_lo_hi_hi_1 = {compressTailMask_elementMask_7, compressTailMask_elementMask_6};
  wire [7:0]    compressTailMask_lo_lo_hi_1 = {compressTailMask_lo_lo_hi_hi_1, compressTailMask_lo_lo_hi_lo_1};
  wire [15:0]   compressTailMask_lo_lo_1 = {compressTailMask_lo_lo_hi_1, compressTailMask_lo_lo_lo_1};
  wire [3:0]    compressTailMask_lo_hi_lo_lo_1 = {compressTailMask_elementMask_9, compressTailMask_elementMask_8};
  wire [3:0]    compressTailMask_lo_hi_lo_hi_1 = {compressTailMask_elementMask_11, compressTailMask_elementMask_10};
  wire [7:0]    compressTailMask_lo_hi_lo_1 = {compressTailMask_lo_hi_lo_hi_1, compressTailMask_lo_hi_lo_lo_1};
  wire [3:0]    compressTailMask_lo_hi_hi_lo_1 = {compressTailMask_elementMask_13, compressTailMask_elementMask_12};
  wire [3:0]    compressTailMask_lo_hi_hi_hi_1 = {compressTailMask_elementMask_15, compressTailMask_elementMask_14};
  wire [7:0]    compressTailMask_lo_hi_hi_1 = {compressTailMask_lo_hi_hi_hi_1, compressTailMask_lo_hi_hi_lo_1};
  wire [15:0]   compressTailMask_lo_hi_1 = {compressTailMask_lo_hi_hi_1, compressTailMask_lo_hi_lo_1};
  wire [31:0]   compressTailMask_lo_1 = {compressTailMask_lo_hi_1, compressTailMask_lo_lo_1};
  wire [3:0]    compressTailMask_hi_lo_lo_lo_1 = {compressTailMask_elementMask_17, compressTailMask_elementMask_16};
  wire [3:0]    compressTailMask_hi_lo_lo_hi_1 = {compressTailMask_elementMask_19, compressTailMask_elementMask_18};
  wire [7:0]    compressTailMask_hi_lo_lo_1 = {compressTailMask_hi_lo_lo_hi_1, compressTailMask_hi_lo_lo_lo_1};
  wire [3:0]    compressTailMask_hi_lo_hi_lo_1 = {compressTailMask_elementMask_21, compressTailMask_elementMask_20};
  wire [3:0]    compressTailMask_hi_lo_hi_hi_1 = {compressTailMask_elementMask_23, compressTailMask_elementMask_22};
  wire [7:0]    compressTailMask_hi_lo_hi_1 = {compressTailMask_hi_lo_hi_hi_1, compressTailMask_hi_lo_hi_lo_1};
  wire [15:0]   compressTailMask_hi_lo_1 = {compressTailMask_hi_lo_hi_1, compressTailMask_hi_lo_lo_1};
  wire [3:0]    compressTailMask_hi_hi_lo_lo_1 = {compressTailMask_elementMask_25, compressTailMask_elementMask_24};
  wire [3:0]    compressTailMask_hi_hi_lo_hi_1 = {compressTailMask_elementMask_27, compressTailMask_elementMask_26};
  wire [7:0]    compressTailMask_hi_hi_lo_1 = {compressTailMask_hi_hi_lo_hi_1, compressTailMask_hi_hi_lo_lo_1};
  wire [3:0]    compressTailMask_hi_hi_hi_lo_1 = {compressTailMask_elementMask_29, compressTailMask_elementMask_28};
  wire [3:0]    compressTailMask_hi_hi_hi_hi_1 = {compressTailMask_elementMask_31, compressTailMask_elementMask_30};
  wire [7:0]    compressTailMask_hi_hi_hi_1 = {compressTailMask_hi_hi_hi_hi_1, compressTailMask_hi_hi_hi_lo_1};
  wire [15:0]   compressTailMask_hi_hi_1 = {compressTailMask_hi_hi_hi_1, compressTailMask_hi_hi_lo_1};
  wire [31:0]   compressTailMask_hi_1 = {compressTailMask_hi_hi_1, compressTailMask_hi_lo_1};
  wire          compressTailMask_elementValid_96;
  assign compressTailMask_elementValid_96 = |tailCountForMask;
  wire [3:0]    compressTailMask_elementMask_32 = {4{compressTailMask_elementValid_96}};
  wire          compressTailMask_elementValid_97;
  assign compressTailMask_elementValid_97 = |(tailCountForMask[5:1]);
  wire [3:0]    compressTailMask_elementMask_33 = {4{compressTailMask_elementValid_97}};
  wire [3:0]    compressTailMask_elementMask_34 = {4{compressTailMask_elementValid_98}};
  wire          compressTailMask_elementValid_99;
  assign compressTailMask_elementValid_99 = |(tailCountForMask[5:2]);
  wire [3:0]    compressTailMask_elementMask_35 = {4{compressTailMask_elementValid_99}};
  wire [3:0]    compressTailMask_elementMask_36 = {4{compressTailMask_elementValid_100}};
  wire [3:0]    compressTailMask_elementMask_37 = {4{compressTailMask_elementValid_101}};
  wire [3:0]    compressTailMask_elementMask_38 = {4{compressTailMask_elementValid_102}};
  wire          compressTailMask_elementValid_103;
  assign compressTailMask_elementValid_103 = |(tailCountForMask[5:3]);
  wire [3:0]    compressTailMask_elementMask_39 = {4{compressTailMask_elementValid_103}};
  wire [3:0]    compressTailMask_elementMask_40 = {4{compressTailMask_elementValid_104}};
  wire [3:0]    compressTailMask_elementMask_41 = {4{compressTailMask_elementValid_105}};
  wire [3:0]    compressTailMask_elementMask_42 = {4{compressTailMask_elementValid_106}};
  wire [3:0]    compressTailMask_elementMask_43 = {4{compressTailMask_elementValid_107}};
  wire [3:0]    compressTailMask_elementMask_44 = {4{compressTailMask_elementValid_108}};
  wire [3:0]    compressTailMask_elementMask_45 = {4{compressTailMask_elementValid_109}};
  wire [3:0]    compressTailMask_elementMask_46 = {4{compressTailMask_elementValid_110}};
  wire          compressTailMask_elementValid_111;
  assign compressTailMask_elementValid_111 = |(tailCountForMask[5:4]);
  wire [3:0]    compressTailMask_elementMask_47 = {4{compressTailMask_elementValid_111}};
  wire [7:0]    compressTailMask_lo_lo_lo_2 = {compressTailMask_elementMask_33, compressTailMask_elementMask_32};
  wire [7:0]    compressTailMask_lo_lo_hi_2 = {compressTailMask_elementMask_35, compressTailMask_elementMask_34};
  wire [15:0]   compressTailMask_lo_lo_2 = {compressTailMask_lo_lo_hi_2, compressTailMask_lo_lo_lo_2};
  wire [7:0]    compressTailMask_lo_hi_lo_2 = {compressTailMask_elementMask_37, compressTailMask_elementMask_36};
  wire [7:0]    compressTailMask_lo_hi_hi_2 = {compressTailMask_elementMask_39, compressTailMask_elementMask_38};
  wire [15:0]   compressTailMask_lo_hi_2 = {compressTailMask_lo_hi_hi_2, compressTailMask_lo_hi_lo_2};
  wire [31:0]   compressTailMask_lo_2 = {compressTailMask_lo_hi_2, compressTailMask_lo_lo_2};
  wire [7:0]    compressTailMask_hi_lo_lo_2 = {compressTailMask_elementMask_41, compressTailMask_elementMask_40};
  wire [7:0]    compressTailMask_hi_lo_hi_2 = {compressTailMask_elementMask_43, compressTailMask_elementMask_42};
  wire [15:0]   compressTailMask_hi_lo_2 = {compressTailMask_hi_lo_hi_2, compressTailMask_hi_lo_lo_2};
  wire [7:0]    compressTailMask_hi_hi_lo_2 = {compressTailMask_elementMask_45, compressTailMask_elementMask_44};
  wire [7:0]    compressTailMask_hi_hi_hi_2 = {compressTailMask_elementMask_47, compressTailMask_elementMask_46};
  wire [15:0]   compressTailMask_hi_hi_2 = {compressTailMask_hi_hi_hi_2, compressTailMask_hi_hi_lo_2};
  wire [31:0]   compressTailMask_hi_2 = {compressTailMask_hi_hi_2, compressTailMask_hi_lo_2};
  wire [63:0]   compressTailMask = (eew1H[0] ? {compressTailMask_hi, compressTailMask_lo} : 64'h0) | (eew1H[1] ? {compressTailMask_hi_1, compressTailMask_lo_1} : 64'h0) | (eew1H[2] ? {compressTailMask_hi_2, compressTailMask_lo_2} : 64'h0);
  wire [63:0]   compressMask = compressTailValid ? compressTailMask : 64'hFFFFFFFFFFFFFFFF;
  reg  [15:0]   validInputPipe;
  reg  [31:0]   readFromScalarPipe;
  wire [3:0]    mvMask = {2'h0, {1'h0, eew1H[0]} | {2{eew1H[1]}}} | {4{eew1H[2]}};
  wire [7:0]    ffoMask_lo_lo_lo = {{4{validInputPipe[1]}}, {4{validInputPipe[0]}}};
  wire [7:0]    ffoMask_lo_lo_hi = {{4{validInputPipe[3]}}, {4{validInputPipe[2]}}};
  wire [15:0]   ffoMask_lo_lo = {ffoMask_lo_lo_hi, ffoMask_lo_lo_lo};
  wire [7:0]    ffoMask_lo_hi_lo = {{4{validInputPipe[5]}}, {4{validInputPipe[4]}}};
  wire [7:0]    ffoMask_lo_hi_hi = {{4{validInputPipe[7]}}, {4{validInputPipe[6]}}};
  wire [15:0]   ffoMask_lo_hi = {ffoMask_lo_hi_hi, ffoMask_lo_hi_lo};
  wire [31:0]   ffoMask_lo = {ffoMask_lo_hi, ffoMask_lo_lo};
  wire [7:0]    ffoMask_hi_lo_lo = {{4{validInputPipe[9]}}, {4{validInputPipe[8]}}};
  wire [7:0]    ffoMask_hi_lo_hi = {{4{validInputPipe[11]}}, {4{validInputPipe[10]}}};
  wire [15:0]   ffoMask_hi_lo = {ffoMask_hi_lo_hi, ffoMask_hi_lo_lo};
  wire [7:0]    ffoMask_hi_hi_lo = {{4{validInputPipe[13]}}, {4{validInputPipe[12]}}};
  wire [7:0]    ffoMask_hi_hi_hi = {{4{validInputPipe[15]}}, {4{validInputPipe[14]}}};
  wire [15:0]   ffoMask_hi_hi = {ffoMask_hi_hi_hi, ffoMask_hi_hi_lo};
  wire [31:0]   ffoMask_hi = {ffoMask_hi_hi, ffoMask_hi_lo};
  wire [63:0]   ffoMask = {ffoMask_hi, ffoMask_lo};
  wire [15:0]   outWire_ffoOutput;
  wire [63:0]   ffoData_lo_lo_lo = {outWire_ffoOutput[1] ? in_1_bits_pipeData[63:32] : in_1_bits_source2[63:32], outWire_ffoOutput[0] ? in_1_bits_pipeData[31:0] : in_1_bits_source2[31:0]};
  wire [63:0]   ffoData_lo_lo_hi = {outWire_ffoOutput[3] ? in_1_bits_pipeData[127:96] : in_1_bits_source2[127:96], outWire_ffoOutput[2] ? in_1_bits_pipeData[95:64] : in_1_bits_source2[95:64]};
  wire [127:0]  ffoData_lo_lo = {ffoData_lo_lo_hi, ffoData_lo_lo_lo};
  wire [63:0]   ffoData_lo_hi_lo = {outWire_ffoOutput[5] ? in_1_bits_pipeData[191:160] : in_1_bits_source2[191:160], outWire_ffoOutput[4] ? in_1_bits_pipeData[159:128] : in_1_bits_source2[159:128]};
  wire [63:0]   ffoData_lo_hi_hi = {outWire_ffoOutput[7] ? in_1_bits_pipeData[255:224] : in_1_bits_source2[255:224], outWire_ffoOutput[6] ? in_1_bits_pipeData[223:192] : in_1_bits_source2[223:192]};
  wire [127:0]  ffoData_lo_hi = {ffoData_lo_hi_hi, ffoData_lo_hi_lo};
  wire [255:0]  ffoData_lo = {ffoData_lo_hi, ffoData_lo_lo};
  wire [63:0]   ffoData_hi_lo_lo = {outWire_ffoOutput[9] ? in_1_bits_pipeData[319:288] : in_1_bits_source2[319:288], outWire_ffoOutput[8] ? in_1_bits_pipeData[287:256] : in_1_bits_source2[287:256]};
  wire [63:0]   ffoData_hi_lo_hi = {outWire_ffoOutput[11] ? in_1_bits_pipeData[383:352] : in_1_bits_source2[383:352], outWire_ffoOutput[10] ? in_1_bits_pipeData[351:320] : in_1_bits_source2[351:320]};
  wire [127:0]  ffoData_hi_lo = {ffoData_hi_lo_hi, ffoData_hi_lo_lo};
  wire [63:0]   ffoData_hi_hi_lo = {outWire_ffoOutput[13] ? in_1_bits_pipeData[447:416] : in_1_bits_source2[447:416], outWire_ffoOutput[12] ? in_1_bits_pipeData[415:384] : in_1_bits_source2[415:384]};
  wire [63:0]   ffoData_hi_hi_hi = {outWire_ffoOutput[15] ? in_1_bits_pipeData[511:480] : in_1_bits_source2[511:480], outWire_ffoOutput[14] ? in_1_bits_pipeData[479:448] : in_1_bits_source2[479:448]};
  wire [127:0]  ffoData_hi_hi = {ffoData_hi_hi_hi, ffoData_hi_hi_lo};
  wire [255:0]  ffoData_hi = {ffoData_hi_hi, ffoData_hi_lo};
  wire [511:0]  ffoData = {ffoData_hi, ffoData_lo};
  wire [511:0]  _GEN_2100 = (compress ? compressResult[511:0] : 512'h0) | (viota ? viotaResult : 512'h0);
  wire [511:0]  outWire_data = {_GEN_2100[511:32], _GEN_2100[31:0] | (mv ? readFromScalarPipe : 32'h0)} | (ffoType ? ffoData : 512'h0);
  wire [63:0]   _outWire_mask_T_4 = (compress ? compressMask : 64'h0) | (viota ? viotaMask : 64'h0);
  wire [63:0]   outWire_mask = {_outWire_mask_T_4[63:4], _outWire_mask_T_4[3:0] | (mv ? mvMask : 4'h0)} | (ffoType ? ffoMask : 64'h0);
  wire          outWire_compressValid = (compressTailValid | compressDeqValidPipe & stage2Valid) & ~writeRD;
  wire [5:0]    outWire_groupCounter = compress ? compressWriteGroupCount : groupCounterPipe;
  wire [14:0]   _completedLeftOr_T_2 = in_1_bits_ffoInput[14:0] | {in_1_bits_ffoInput[13:0], 1'h0};
  wire [14:0]   _GEN_2101 = {_completedLeftOr_T_2[12:0], 2'h0};
  wire [14:0]   _firstLane_T_5 = _completedLeftOr_T_2 | _GEN_2101;
  wire [14:0]   _firstLane_T_8 = _firstLane_T_5 | {_firstLane_T_5[10:0], 4'h0};
  wire [15:0]   firstLane = {~(_firstLane_T_8 | {_firstLane_T_8[6:0], 8'h0}), 1'h1} & in_1_bits_ffoInput;
  wire [7:0]    firstLaneIndex_hi = firstLane[15:8];
  wire [7:0]    firstLaneIndex_lo = firstLane[7:0];
  wire [7:0]    _firstLaneIndex_T_1 = firstLaneIndex_hi | firstLaneIndex_lo;
  wire [3:0]    firstLaneIndex_hi_1 = _firstLaneIndex_T_1[7:4];
  wire [3:0]    firstLaneIndex_lo_1 = _firstLaneIndex_T_1[3:0];
  wire [3:0]    _firstLaneIndex_T_3 = firstLaneIndex_hi_1 | firstLaneIndex_lo_1;
  wire [1:0]    firstLaneIndex_hi_2 = _firstLaneIndex_T_3[3:2];
  wire [1:0]    firstLaneIndex_lo_2 = _firstLaneIndex_T_3[1:0];
  wire [3:0]    firstLaneIndex = {|firstLaneIndex_hi, |firstLaneIndex_hi_1, |firstLaneIndex_hi_2, firstLaneIndex_hi_2[1] | firstLaneIndex_lo_2[1]};
  wire [31:0]   source1SigExtend = (eew1H[0] ? {{24{in_1_bits_source1[7]}}, in_1_bits_source1[7:0]} : 32'h0) | (eew1H[1] ? {{16{in_1_bits_source1[15]}}, in_1_bits_source1[15:0]} : 32'h0) | (eew1H[2] ? in_1_bits_source1 : 32'h0);
  wire [14:0]   _completedLeftOr_T_5 = _completedLeftOr_T_2 | _GEN_2101;
  wire [14:0]   _completedLeftOr_T_8 = _completedLeftOr_T_5 | {_completedLeftOr_T_5[10:0], 4'h0};
  wire [15:0]   completedLeftOr = {_completedLeftOr_T_8 | {_completedLeftOr_T_8[6:0], 8'h0}, 1'h0};
  reg  [15:0]   ffoOutPipe;
  assign outWire_ffoOutput = ffoOutPipe;
  reg  [511:0]  view__out_REG_data;
  reg  [63:0]   view__out_REG_mask;
  reg  [5:0]    view__out_REG_groupCounter;
  reg  [15:0]   view__out_REG_ffoOutput;
  reg           view__out_REG_compressValid;
  always @(posedge clock) begin
    if (reset) begin
      in_1_valid <= 1'h0;
      in_1_bits_maskType <= 1'h0;
      in_1_bits_eew <= 2'h0;
      in_1_bits_uop <= 3'h0;
      in_1_bits_readFromScalar <= 32'h0;
      in_1_bits_source1 <= 32'h0;
      in_1_bits_mask <= 32'h0;
      in_1_bits_source2 <= 512'h0;
      in_1_bits_pipeData <= 512'h0;
      in_1_bits_groupCounter <= 6'h0;
      in_1_bits_ffoInput <= 16'h0;
      in_1_bits_validInput <= 16'h0;
      in_1_bits_lastCompress <= 1'h0;
      compressInit <= 11'h0;
      ffoIndex <= 32'h0;
      ffoValid <= 1'h0;
      compressVecPipe_0 <= 11'h0;
      compressVecPipe_1 <= 11'h0;
      compressVecPipe_2 <= 11'h0;
      compressVecPipe_3 <= 11'h0;
      compressVecPipe_4 <= 11'h0;
      compressVecPipe_5 <= 11'h0;
      compressVecPipe_6 <= 11'h0;
      compressVecPipe_7 <= 11'h0;
      compressVecPipe_8 <= 11'h0;
      compressVecPipe_9 <= 11'h0;
      compressVecPipe_10 <= 11'h0;
      compressVecPipe_11 <= 11'h0;
      compressVecPipe_12 <= 11'h0;
      compressVecPipe_13 <= 11'h0;
      compressVecPipe_14 <= 11'h0;
      compressVecPipe_15 <= 11'h0;
      compressVecPipe_16 <= 11'h0;
      compressVecPipe_17 <= 11'h0;
      compressVecPipe_18 <= 11'h0;
      compressVecPipe_19 <= 11'h0;
      compressVecPipe_20 <= 11'h0;
      compressVecPipe_21 <= 11'h0;
      compressVecPipe_22 <= 11'h0;
      compressVecPipe_23 <= 11'h0;
      compressVecPipe_24 <= 11'h0;
      compressVecPipe_25 <= 11'h0;
      compressVecPipe_26 <= 11'h0;
      compressVecPipe_27 <= 11'h0;
      compressVecPipe_28 <= 11'h0;
      compressVecPipe_29 <= 11'h0;
      compressVecPipe_30 <= 11'h0;
      compressVecPipe_31 <= 11'h0;
      compressVecPipe_32 <= 11'h0;
      compressVecPipe_33 <= 11'h0;
      compressVecPipe_34 <= 11'h0;
      compressVecPipe_35 <= 11'h0;
      compressVecPipe_36 <= 11'h0;
      compressVecPipe_37 <= 11'h0;
      compressVecPipe_38 <= 11'h0;
      compressVecPipe_39 <= 11'h0;
      compressVecPipe_40 <= 11'h0;
      compressVecPipe_41 <= 11'h0;
      compressVecPipe_42 <= 11'h0;
      compressVecPipe_43 <= 11'h0;
      compressVecPipe_44 <= 11'h0;
      compressVecPipe_45 <= 11'h0;
      compressVecPipe_46 <= 11'h0;
      compressVecPipe_47 <= 11'h0;
      compressVecPipe_48 <= 11'h0;
      compressVecPipe_49 <= 11'h0;
      compressVecPipe_50 <= 11'h0;
      compressVecPipe_51 <= 11'h0;
      compressVecPipe_52 <= 11'h0;
      compressVecPipe_53 <= 11'h0;
      compressVecPipe_54 <= 11'h0;
      compressVecPipe_55 <= 11'h0;
      compressVecPipe_56 <= 11'h0;
      compressVecPipe_57 <= 11'h0;
      compressVecPipe_58 <= 11'h0;
      compressVecPipe_59 <= 11'h0;
      compressVecPipe_60 <= 11'h0;
      compressVecPipe_61 <= 11'h0;
      compressVecPipe_62 <= 11'h0;
      compressVecPipe_63 <= 11'h0;
      compressMaskVecPipe_0 <= 1'h0;
      compressMaskVecPipe_1 <= 1'h0;
      compressMaskVecPipe_2 <= 1'h0;
      compressMaskVecPipe_3 <= 1'h0;
      compressMaskVecPipe_4 <= 1'h0;
      compressMaskVecPipe_5 <= 1'h0;
      compressMaskVecPipe_6 <= 1'h0;
      compressMaskVecPipe_7 <= 1'h0;
      compressMaskVecPipe_8 <= 1'h0;
      compressMaskVecPipe_9 <= 1'h0;
      compressMaskVecPipe_10 <= 1'h0;
      compressMaskVecPipe_11 <= 1'h0;
      compressMaskVecPipe_12 <= 1'h0;
      compressMaskVecPipe_13 <= 1'h0;
      compressMaskVecPipe_14 <= 1'h0;
      compressMaskVecPipe_15 <= 1'h0;
      compressMaskVecPipe_16 <= 1'h0;
      compressMaskVecPipe_17 <= 1'h0;
      compressMaskVecPipe_18 <= 1'h0;
      compressMaskVecPipe_19 <= 1'h0;
      compressMaskVecPipe_20 <= 1'h0;
      compressMaskVecPipe_21 <= 1'h0;
      compressMaskVecPipe_22 <= 1'h0;
      compressMaskVecPipe_23 <= 1'h0;
      compressMaskVecPipe_24 <= 1'h0;
      compressMaskVecPipe_25 <= 1'h0;
      compressMaskVecPipe_26 <= 1'h0;
      compressMaskVecPipe_27 <= 1'h0;
      compressMaskVecPipe_28 <= 1'h0;
      compressMaskVecPipe_29 <= 1'h0;
      compressMaskVecPipe_30 <= 1'h0;
      compressMaskVecPipe_31 <= 1'h0;
      compressMaskVecPipe_32 <= 1'h0;
      compressMaskVecPipe_33 <= 1'h0;
      compressMaskVecPipe_34 <= 1'h0;
      compressMaskVecPipe_35 <= 1'h0;
      compressMaskVecPipe_36 <= 1'h0;
      compressMaskVecPipe_37 <= 1'h0;
      compressMaskVecPipe_38 <= 1'h0;
      compressMaskVecPipe_39 <= 1'h0;
      compressMaskVecPipe_40 <= 1'h0;
      compressMaskVecPipe_41 <= 1'h0;
      compressMaskVecPipe_42 <= 1'h0;
      compressMaskVecPipe_43 <= 1'h0;
      compressMaskVecPipe_44 <= 1'h0;
      compressMaskVecPipe_45 <= 1'h0;
      compressMaskVecPipe_46 <= 1'h0;
      compressMaskVecPipe_47 <= 1'h0;
      compressMaskVecPipe_48 <= 1'h0;
      compressMaskVecPipe_49 <= 1'h0;
      compressMaskVecPipe_50 <= 1'h0;
      compressMaskVecPipe_51 <= 1'h0;
      compressMaskVecPipe_52 <= 1'h0;
      compressMaskVecPipe_53 <= 1'h0;
      compressMaskVecPipe_54 <= 1'h0;
      compressMaskVecPipe_55 <= 1'h0;
      compressMaskVecPipe_56 <= 1'h0;
      compressMaskVecPipe_57 <= 1'h0;
      compressMaskVecPipe_58 <= 1'h0;
      compressMaskVecPipe_59 <= 1'h0;
      compressMaskVecPipe_60 <= 1'h0;
      compressMaskVecPipe_61 <= 1'h0;
      compressMaskVecPipe_62 <= 1'h0;
      compressMaskVecPipe_63 <= 1'h0;
      maskPipe <= 32'h0;
      source2Pipe <= 512'h0;
      lastCompressPipe <= 1'h0;
      stage2Valid <= 1'h0;
      newInstructionPipe <= 1'h0;
      compressInitPipe <= 11'h0;
      compressDeqValidPipe <= 1'h0;
      groupCounterPipe <= 6'h0;
      compressDataReg <= 512'h0;
      compressTailValid <= 1'h0;
      compressWriteGroupCount <= 6'h0;
      validInputPipe <= 16'h0;
      readFromScalarPipe <= 32'h0;
      ffoOutPipe <= 16'h0;
      view__out_REG_data <= 512'h0;
      view__out_REG_mask <= 64'h0;
      view__out_REG_groupCounter <= 6'h0;
      view__out_REG_ffoOutput <= 16'h0;
      view__out_REG_compressValid <= 1'h0;
    end
    else begin
      automatic logic _GEN_2102;
      automatic logic _GEN_2103;
      _GEN_2102 = newInstruction & ffoInstruction;
      _GEN_2103 = in_1_valid & (|in_1_bits_ffoInput) & ffoType;
      in_1_valid <= in_valid;
      in_1_bits_maskType <= in_bits_maskType;
      in_1_bits_eew <= in_bits_eew;
      in_1_bits_uop <= in_bits_uop;
      in_1_bits_readFromScalar <= in_bits_readFromScalar;
      in_1_bits_source1 <= in_bits_source1;
      in_1_bits_mask <= in_bits_mask;
      in_1_bits_source2 <= in_bits_source2;
      in_1_bits_pipeData <= in_bits_pipeData;
      in_1_bits_groupCounter <= in_bits_groupCounter;
      in_1_bits_ffoInput <= in_bits_ffoInput;
      in_1_bits_validInput <= in_bits_validInput;
      in_1_bits_lastCompress <= in_bits_lastCompress;
      if (in_1_valid) begin
        compressInit <= viota ? compressCount : {5'h0, compressCountSelect};
        compressVecPipe_0 <= compressVec_0;
        compressVecPipe_1 <= compressVec_1;
        compressVecPipe_2 <= compressVec_2;
        compressVecPipe_3 <= compressVec_3;
        compressVecPipe_4 <= compressVec_4;
        compressVecPipe_5 <= compressVec_5;
        compressVecPipe_6 <= compressVec_6;
        compressVecPipe_7 <= compressVec_7;
        compressVecPipe_8 <= compressVec_8;
        compressVecPipe_9 <= compressVec_9;
        compressVecPipe_10 <= compressVec_10;
        compressVecPipe_11 <= compressVec_11;
        compressVecPipe_12 <= compressVec_12;
        compressVecPipe_13 <= compressVec_13;
        compressVecPipe_14 <= compressVec_14;
        compressVecPipe_15 <= compressVec_15;
        compressVecPipe_16 <= compressVec_16;
        compressVecPipe_17 <= compressVec_17;
        compressVecPipe_18 <= compressVec_18;
        compressVecPipe_19 <= compressVec_19;
        compressVecPipe_20 <= compressVec_20;
        compressVecPipe_21 <= compressVec_21;
        compressVecPipe_22 <= compressVec_22;
        compressVecPipe_23 <= compressVec_23;
        compressVecPipe_24 <= compressVec_24;
        compressVecPipe_25 <= compressVec_25;
        compressVecPipe_26 <= compressVec_26;
        compressVecPipe_27 <= compressVec_27;
        compressVecPipe_28 <= compressVec_28;
        compressVecPipe_29 <= compressVec_29;
        compressVecPipe_30 <= compressVec_30;
        compressVecPipe_31 <= compressVec_31;
        compressVecPipe_32 <= compressVec_32;
        compressVecPipe_33 <= compressVec_33;
        compressVecPipe_34 <= compressVec_34;
        compressVecPipe_35 <= compressVec_35;
        compressVecPipe_36 <= compressVec_36;
        compressVecPipe_37 <= compressVec_37;
        compressVecPipe_38 <= compressVec_38;
        compressVecPipe_39 <= compressVec_39;
        compressVecPipe_40 <= compressVec_40;
        compressVecPipe_41 <= compressVec_41;
        compressVecPipe_42 <= compressVec_42;
        compressVecPipe_43 <= compressVec_43;
        compressVecPipe_44 <= compressVec_44;
        compressVecPipe_45 <= compressVec_45;
        compressVecPipe_46 <= compressVec_46;
        compressVecPipe_47 <= compressVec_47;
        compressVecPipe_48 <= compressVec_48;
        compressVecPipe_49 <= compressVec_49;
        compressVecPipe_50 <= compressVec_50;
        compressVecPipe_51 <= compressVec_51;
        compressVecPipe_52 <= compressVec_52;
        compressVecPipe_53 <= compressVec_53;
        compressVecPipe_54 <= compressVec_54;
        compressVecPipe_55 <= compressVec_55;
        compressVecPipe_56 <= compressVec_56;
        compressVecPipe_57 <= compressVec_57;
        compressVecPipe_58 <= compressVec_58;
        compressVecPipe_59 <= compressVec_59;
        compressVecPipe_60 <= compressVec_60;
        compressVecPipe_61 <= compressVec_61;
        compressVecPipe_62 <= compressVec_62;
        compressVecPipe_63 <= compressVec_63;
        compressMaskVecPipe_0 <= compressMaskVec_0;
        compressMaskVecPipe_1 <= compressMaskVec_1;
        compressMaskVecPipe_2 <= compressMaskVec_2;
        compressMaskVecPipe_3 <= compressMaskVec_3;
        compressMaskVecPipe_4 <= compressMaskVec_4;
        compressMaskVecPipe_5 <= compressMaskVec_5;
        compressMaskVecPipe_6 <= compressMaskVec_6;
        compressMaskVecPipe_7 <= compressMaskVec_7;
        compressMaskVecPipe_8 <= compressMaskVec_8;
        compressMaskVecPipe_9 <= compressMaskVec_9;
        compressMaskVecPipe_10 <= compressMaskVec_10;
        compressMaskVecPipe_11 <= compressMaskVec_11;
        compressMaskVecPipe_12 <= compressMaskVec_12;
        compressMaskVecPipe_13 <= compressMaskVec_13;
        compressMaskVecPipe_14 <= compressMaskVec_14;
        compressMaskVecPipe_15 <= compressMaskVec_15;
        compressMaskVecPipe_16 <= compressMaskVec_16;
        compressMaskVecPipe_17 <= compressMaskVec_17;
        compressMaskVecPipe_18 <= compressMaskVec_18;
        compressMaskVecPipe_19 <= compressMaskVec_19;
        compressMaskVecPipe_20 <= compressMaskVec_20;
        compressMaskVecPipe_21 <= compressMaskVec_21;
        compressMaskVecPipe_22 <= compressMaskVec_22;
        compressMaskVecPipe_23 <= compressMaskVec_23;
        compressMaskVecPipe_24 <= compressMaskVec_24;
        compressMaskVecPipe_25 <= compressMaskVec_25;
        compressMaskVecPipe_26 <= compressMaskVec_26;
        compressMaskVecPipe_27 <= compressMaskVec_27;
        compressMaskVecPipe_28 <= compressMaskVec_28;
        compressMaskVecPipe_29 <= compressMaskVec_29;
        compressMaskVecPipe_30 <= compressMaskVec_30;
        compressMaskVecPipe_31 <= compressMaskVec_31;
        compressMaskVecPipe_32 <= compressMaskVec_32;
        compressMaskVecPipe_33 <= compressMaskVec_33;
        compressMaskVecPipe_34 <= compressMaskVec_34;
        compressMaskVecPipe_35 <= compressMaskVec_35;
        compressMaskVecPipe_36 <= compressMaskVec_36;
        compressMaskVecPipe_37 <= compressMaskVec_37;
        compressMaskVecPipe_38 <= compressMaskVec_38;
        compressMaskVecPipe_39 <= compressMaskVec_39;
        compressMaskVecPipe_40 <= compressMaskVec_40;
        compressMaskVecPipe_41 <= compressMaskVec_41;
        compressMaskVecPipe_42 <= compressMaskVec_42;
        compressMaskVecPipe_43 <= compressMaskVec_43;
        compressMaskVecPipe_44 <= compressMaskVec_44;
        compressMaskVecPipe_45 <= compressMaskVec_45;
        compressMaskVecPipe_46 <= compressMaskVec_46;
        compressMaskVecPipe_47 <= compressMaskVec_47;
        compressMaskVecPipe_48 <= compressMaskVec_48;
        compressMaskVecPipe_49 <= compressMaskVec_49;
        compressMaskVecPipe_50 <= compressMaskVec_50;
        compressMaskVecPipe_51 <= compressMaskVec_51;
        compressMaskVecPipe_52 <= compressMaskVec_52;
        compressMaskVecPipe_53 <= compressMaskVec_53;
        compressMaskVecPipe_54 <= compressMaskVec_54;
        compressMaskVecPipe_55 <= compressMaskVec_55;
        compressMaskVecPipe_56 <= compressMaskVec_56;
        compressMaskVecPipe_57 <= compressMaskVec_57;
        compressMaskVecPipe_58 <= compressMaskVec_58;
        compressMaskVecPipe_59 <= compressMaskVec_59;
        compressMaskVecPipe_60 <= compressMaskVec_60;
        compressMaskVecPipe_61 <= compressMaskVec_61;
        compressMaskVecPipe_62 <= compressMaskVec_62;
        compressMaskVecPipe_63 <= compressMaskVec_63;
        maskPipe <= in_1_bits_mask;
        source2Pipe <= in_1_bits_source2;
        lastCompressPipe <= in_1_bits_lastCompress;
        compressInitPipe <= compressInit;
        compressDeqValidPipe <= compressDeqValid;
        groupCounterPipe <= in_1_bits_groupCounter;
        validInputPipe <= in_1_bits_validInput;
        readFromScalarPipe <= in_1_bits_readFromScalar;
        ffoOutPipe <= completedLeftOr | {16{ffoValid}};
      end
      else if (newInstruction)
        compressInit <= 11'h0;
      if (_GEN_2103) begin
        if (ffoValid) begin
          if (_GEN_2102)
            ffoIndex <= 32'hFFFFFFFF;
        end
        else
          ffoIndex <=
            (firstLane[0] ? {in_1_bits_source2[27:5], firstLaneIndex, in_1_bits_source2[4:0]} : 32'h0) | (firstLane[1] ? {in_1_bits_source2[59:37], firstLaneIndex, in_1_bits_source2[36:32]} : 32'h0)
            | (firstLane[2] ? {in_1_bits_source2[91:69], firstLaneIndex, in_1_bits_source2[68:64]} : 32'h0) | (firstLane[3] ? {in_1_bits_source2[123:101], firstLaneIndex, in_1_bits_source2[100:96]} : 32'h0)
            | (firstLane[4] ? {in_1_bits_source2[155:133], firstLaneIndex, in_1_bits_source2[132:128]} : 32'h0) | (firstLane[5] ? {in_1_bits_source2[187:165], firstLaneIndex, in_1_bits_source2[164:160]} : 32'h0)
            | (firstLane[6] ? {in_1_bits_source2[219:197], firstLaneIndex, in_1_bits_source2[196:192]} : 32'h0) | (firstLane[7] ? {in_1_bits_source2[251:229], firstLaneIndex, in_1_bits_source2[228:224]} : 32'h0)
            | (firstLane[8] ? {in_1_bits_source2[283:261], firstLaneIndex, in_1_bits_source2[260:256]} : 32'h0) | (firstLane[9] ? {in_1_bits_source2[315:293], firstLaneIndex, in_1_bits_source2[292:288]} : 32'h0)
            | (firstLane[10] ? {in_1_bits_source2[347:325], firstLaneIndex, in_1_bits_source2[324:320]} : 32'h0) | (firstLane[11] ? {in_1_bits_source2[379:357], firstLaneIndex, in_1_bits_source2[356:352]} : 32'h0)
            | (firstLane[12] ? {in_1_bits_source2[411:389], firstLaneIndex, in_1_bits_source2[388:384]} : 32'h0) | (firstLane[13] ? {in_1_bits_source2[443:421], firstLaneIndex, in_1_bits_source2[420:416]} : 32'h0)
            | (firstLane[14] ? {in_1_bits_source2[475:453], firstLaneIndex, in_1_bits_source2[452:448]} : 32'h0) | (firstLane[15] ? {in_1_bits_source2[507:485], firstLaneIndex, in_1_bits_source2[484:480]} : 32'h0);
      end
      else if (mvRd)
        ffoIndex <= source1SigExtend;
      else if (_GEN_2102)
        ffoIndex <= 32'hFFFFFFFF;
      ffoValid <= _GEN_2103 | ~_GEN_2102 & ffoValid;
      stage2Valid <= in_1_valid;
      newInstructionPipe <= newInstruction;
      if (stage2Valid)
        compressDataReg <= compressDeqValidPipe ? splitCompressResult_1 : splitCompressResult_0;
      if (newInstructionPipe | lastCompressEnq | outWire_compressValid)
        compressTailValid <= lastCompressEnq & compress;
      if (newInstructionPipe | outWire_compressValid)
        compressWriteGroupCount <= newInstructionPipe ? 6'h0 : compressWriteGroupCount + 6'h1;
      view__out_REG_data <= outWire_data;
      view__out_REG_mask <= outWire_mask;
      view__out_REG_groupCounter <= outWire_groupCounter;
      view__out_REG_ffoOutput <= outWire_ffoOutput;
      view__out_REG_compressValid <= outWire_compressValid;
    end
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:116];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [6:0] i = 7'h0; i < 7'h75; i += 7'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        in_1_valid = _RANDOM[7'h0][0];
        in_1_bits_maskType = _RANDOM[7'h0][1];
        in_1_bits_eew = _RANDOM[7'h0][3:2];
        in_1_bits_uop = _RANDOM[7'h0][6:4];
        in_1_bits_readFromScalar = {_RANDOM[7'h0][31:7], _RANDOM[7'h1][6:0]};
        in_1_bits_source1 = {_RANDOM[7'h1][31:7], _RANDOM[7'h2][6:0]};
        in_1_bits_mask = {_RANDOM[7'h2][31:7], _RANDOM[7'h3][6:0]};
        in_1_bits_source2 =
          {_RANDOM[7'h3][31:7],
           _RANDOM[7'h4],
           _RANDOM[7'h5],
           _RANDOM[7'h6],
           _RANDOM[7'h7],
           _RANDOM[7'h8],
           _RANDOM[7'h9],
           _RANDOM[7'hA],
           _RANDOM[7'hB],
           _RANDOM[7'hC],
           _RANDOM[7'hD],
           _RANDOM[7'hE],
           _RANDOM[7'hF],
           _RANDOM[7'h10],
           _RANDOM[7'h11],
           _RANDOM[7'h12],
           _RANDOM[7'h13][6:0]};
        in_1_bits_pipeData =
          {_RANDOM[7'h13][31:7],
           _RANDOM[7'h14],
           _RANDOM[7'h15],
           _RANDOM[7'h16],
           _RANDOM[7'h17],
           _RANDOM[7'h18],
           _RANDOM[7'h19],
           _RANDOM[7'h1A],
           _RANDOM[7'h1B],
           _RANDOM[7'h1C],
           _RANDOM[7'h1D],
           _RANDOM[7'h1E],
           _RANDOM[7'h1F],
           _RANDOM[7'h20],
           _RANDOM[7'h21],
           _RANDOM[7'h22],
           _RANDOM[7'h23][6:0]};
        in_1_bits_groupCounter = _RANDOM[7'h23][12:7];
        in_1_bits_ffoInput = _RANDOM[7'h23][28:13];
        in_1_bits_validInput = {_RANDOM[7'h23][31:29], _RANDOM[7'h24][12:0]};
        in_1_bits_lastCompress = _RANDOM[7'h24][13];
        compressInit = _RANDOM[7'h24][24:14];
        ffoIndex = {_RANDOM[7'h24][31:25], _RANDOM[7'h25][24:0]};
        ffoValid = _RANDOM[7'h25][25];
        compressVecPipe_0 = {_RANDOM[7'h25][31:26], _RANDOM[7'h26][4:0]};
        compressVecPipe_1 = _RANDOM[7'h26][15:5];
        compressVecPipe_2 = _RANDOM[7'h26][26:16];
        compressVecPipe_3 = {_RANDOM[7'h26][31:27], _RANDOM[7'h27][5:0]};
        compressVecPipe_4 = _RANDOM[7'h27][16:6];
        compressVecPipe_5 = _RANDOM[7'h27][27:17];
        compressVecPipe_6 = {_RANDOM[7'h27][31:28], _RANDOM[7'h28][6:0]};
        compressVecPipe_7 = _RANDOM[7'h28][17:7];
        compressVecPipe_8 = _RANDOM[7'h28][28:18];
        compressVecPipe_9 = {_RANDOM[7'h28][31:29], _RANDOM[7'h29][7:0]};
        compressVecPipe_10 = _RANDOM[7'h29][18:8];
        compressVecPipe_11 = _RANDOM[7'h29][29:19];
        compressVecPipe_12 = {_RANDOM[7'h29][31:30], _RANDOM[7'h2A][8:0]};
        compressVecPipe_13 = _RANDOM[7'h2A][19:9];
        compressVecPipe_14 = _RANDOM[7'h2A][30:20];
        compressVecPipe_15 = {_RANDOM[7'h2A][31], _RANDOM[7'h2B][9:0]};
        compressVecPipe_16 = _RANDOM[7'h2B][20:10];
        compressVecPipe_17 = _RANDOM[7'h2B][31:21];
        compressVecPipe_18 = _RANDOM[7'h2C][10:0];
        compressVecPipe_19 = _RANDOM[7'h2C][21:11];
        compressVecPipe_20 = {_RANDOM[7'h2C][31:22], _RANDOM[7'h2D][0]};
        compressVecPipe_21 = _RANDOM[7'h2D][11:1];
        compressVecPipe_22 = _RANDOM[7'h2D][22:12];
        compressVecPipe_23 = {_RANDOM[7'h2D][31:23], _RANDOM[7'h2E][1:0]};
        compressVecPipe_24 = _RANDOM[7'h2E][12:2];
        compressVecPipe_25 = _RANDOM[7'h2E][23:13];
        compressVecPipe_26 = {_RANDOM[7'h2E][31:24], _RANDOM[7'h2F][2:0]};
        compressVecPipe_27 = _RANDOM[7'h2F][13:3];
        compressVecPipe_28 = _RANDOM[7'h2F][24:14];
        compressVecPipe_29 = {_RANDOM[7'h2F][31:25], _RANDOM[7'h30][3:0]};
        compressVecPipe_30 = _RANDOM[7'h30][14:4];
        compressVecPipe_31 = _RANDOM[7'h30][25:15];
        compressVecPipe_32 = {_RANDOM[7'h30][31:26], _RANDOM[7'h31][4:0]};
        compressVecPipe_33 = _RANDOM[7'h31][15:5];
        compressVecPipe_34 = _RANDOM[7'h31][26:16];
        compressVecPipe_35 = {_RANDOM[7'h31][31:27], _RANDOM[7'h32][5:0]};
        compressVecPipe_36 = _RANDOM[7'h32][16:6];
        compressVecPipe_37 = _RANDOM[7'h32][27:17];
        compressVecPipe_38 = {_RANDOM[7'h32][31:28], _RANDOM[7'h33][6:0]};
        compressVecPipe_39 = _RANDOM[7'h33][17:7];
        compressVecPipe_40 = _RANDOM[7'h33][28:18];
        compressVecPipe_41 = {_RANDOM[7'h33][31:29], _RANDOM[7'h34][7:0]};
        compressVecPipe_42 = _RANDOM[7'h34][18:8];
        compressVecPipe_43 = _RANDOM[7'h34][29:19];
        compressVecPipe_44 = {_RANDOM[7'h34][31:30], _RANDOM[7'h35][8:0]};
        compressVecPipe_45 = _RANDOM[7'h35][19:9];
        compressVecPipe_46 = _RANDOM[7'h35][30:20];
        compressVecPipe_47 = {_RANDOM[7'h35][31], _RANDOM[7'h36][9:0]};
        compressVecPipe_48 = _RANDOM[7'h36][20:10];
        compressVecPipe_49 = _RANDOM[7'h36][31:21];
        compressVecPipe_50 = _RANDOM[7'h37][10:0];
        compressVecPipe_51 = _RANDOM[7'h37][21:11];
        compressVecPipe_52 = {_RANDOM[7'h37][31:22], _RANDOM[7'h38][0]};
        compressVecPipe_53 = _RANDOM[7'h38][11:1];
        compressVecPipe_54 = _RANDOM[7'h38][22:12];
        compressVecPipe_55 = {_RANDOM[7'h38][31:23], _RANDOM[7'h39][1:0]};
        compressVecPipe_56 = _RANDOM[7'h39][12:2];
        compressVecPipe_57 = _RANDOM[7'h39][23:13];
        compressVecPipe_58 = {_RANDOM[7'h39][31:24], _RANDOM[7'h3A][2:0]};
        compressVecPipe_59 = _RANDOM[7'h3A][13:3];
        compressVecPipe_60 = _RANDOM[7'h3A][24:14];
        compressVecPipe_61 = {_RANDOM[7'h3A][31:25], _RANDOM[7'h3B][3:0]};
        compressVecPipe_62 = _RANDOM[7'h3B][14:4];
        compressVecPipe_63 = _RANDOM[7'h3B][25:15];
        compressMaskVecPipe_0 = _RANDOM[7'h3B][26];
        compressMaskVecPipe_1 = _RANDOM[7'h3B][27];
        compressMaskVecPipe_2 = _RANDOM[7'h3B][28];
        compressMaskVecPipe_3 = _RANDOM[7'h3B][29];
        compressMaskVecPipe_4 = _RANDOM[7'h3B][30];
        compressMaskVecPipe_5 = _RANDOM[7'h3B][31];
        compressMaskVecPipe_6 = _RANDOM[7'h3C][0];
        compressMaskVecPipe_7 = _RANDOM[7'h3C][1];
        compressMaskVecPipe_8 = _RANDOM[7'h3C][2];
        compressMaskVecPipe_9 = _RANDOM[7'h3C][3];
        compressMaskVecPipe_10 = _RANDOM[7'h3C][4];
        compressMaskVecPipe_11 = _RANDOM[7'h3C][5];
        compressMaskVecPipe_12 = _RANDOM[7'h3C][6];
        compressMaskVecPipe_13 = _RANDOM[7'h3C][7];
        compressMaskVecPipe_14 = _RANDOM[7'h3C][8];
        compressMaskVecPipe_15 = _RANDOM[7'h3C][9];
        compressMaskVecPipe_16 = _RANDOM[7'h3C][10];
        compressMaskVecPipe_17 = _RANDOM[7'h3C][11];
        compressMaskVecPipe_18 = _RANDOM[7'h3C][12];
        compressMaskVecPipe_19 = _RANDOM[7'h3C][13];
        compressMaskVecPipe_20 = _RANDOM[7'h3C][14];
        compressMaskVecPipe_21 = _RANDOM[7'h3C][15];
        compressMaskVecPipe_22 = _RANDOM[7'h3C][16];
        compressMaskVecPipe_23 = _RANDOM[7'h3C][17];
        compressMaskVecPipe_24 = _RANDOM[7'h3C][18];
        compressMaskVecPipe_25 = _RANDOM[7'h3C][19];
        compressMaskVecPipe_26 = _RANDOM[7'h3C][20];
        compressMaskVecPipe_27 = _RANDOM[7'h3C][21];
        compressMaskVecPipe_28 = _RANDOM[7'h3C][22];
        compressMaskVecPipe_29 = _RANDOM[7'h3C][23];
        compressMaskVecPipe_30 = _RANDOM[7'h3C][24];
        compressMaskVecPipe_31 = _RANDOM[7'h3C][25];
        compressMaskVecPipe_32 = _RANDOM[7'h3C][26];
        compressMaskVecPipe_33 = _RANDOM[7'h3C][27];
        compressMaskVecPipe_34 = _RANDOM[7'h3C][28];
        compressMaskVecPipe_35 = _RANDOM[7'h3C][29];
        compressMaskVecPipe_36 = _RANDOM[7'h3C][30];
        compressMaskVecPipe_37 = _RANDOM[7'h3C][31];
        compressMaskVecPipe_38 = _RANDOM[7'h3D][0];
        compressMaskVecPipe_39 = _RANDOM[7'h3D][1];
        compressMaskVecPipe_40 = _RANDOM[7'h3D][2];
        compressMaskVecPipe_41 = _RANDOM[7'h3D][3];
        compressMaskVecPipe_42 = _RANDOM[7'h3D][4];
        compressMaskVecPipe_43 = _RANDOM[7'h3D][5];
        compressMaskVecPipe_44 = _RANDOM[7'h3D][6];
        compressMaskVecPipe_45 = _RANDOM[7'h3D][7];
        compressMaskVecPipe_46 = _RANDOM[7'h3D][8];
        compressMaskVecPipe_47 = _RANDOM[7'h3D][9];
        compressMaskVecPipe_48 = _RANDOM[7'h3D][10];
        compressMaskVecPipe_49 = _RANDOM[7'h3D][11];
        compressMaskVecPipe_50 = _RANDOM[7'h3D][12];
        compressMaskVecPipe_51 = _RANDOM[7'h3D][13];
        compressMaskVecPipe_52 = _RANDOM[7'h3D][14];
        compressMaskVecPipe_53 = _RANDOM[7'h3D][15];
        compressMaskVecPipe_54 = _RANDOM[7'h3D][16];
        compressMaskVecPipe_55 = _RANDOM[7'h3D][17];
        compressMaskVecPipe_56 = _RANDOM[7'h3D][18];
        compressMaskVecPipe_57 = _RANDOM[7'h3D][19];
        compressMaskVecPipe_58 = _RANDOM[7'h3D][20];
        compressMaskVecPipe_59 = _RANDOM[7'h3D][21];
        compressMaskVecPipe_60 = _RANDOM[7'h3D][22];
        compressMaskVecPipe_61 = _RANDOM[7'h3D][23];
        compressMaskVecPipe_62 = _RANDOM[7'h3D][24];
        compressMaskVecPipe_63 = _RANDOM[7'h3D][25];
        maskPipe = {_RANDOM[7'h3D][31:26], _RANDOM[7'h3E][25:0]};
        source2Pipe =
          {_RANDOM[7'h3E][31:26],
           _RANDOM[7'h3F],
           _RANDOM[7'h40],
           _RANDOM[7'h41],
           _RANDOM[7'h42],
           _RANDOM[7'h43],
           _RANDOM[7'h44],
           _RANDOM[7'h45],
           _RANDOM[7'h46],
           _RANDOM[7'h47],
           _RANDOM[7'h48],
           _RANDOM[7'h49],
           _RANDOM[7'h4A],
           _RANDOM[7'h4B],
           _RANDOM[7'h4C],
           _RANDOM[7'h4D],
           _RANDOM[7'h4E][25:0]};
        lastCompressPipe = _RANDOM[7'h4E][26];
        stage2Valid = _RANDOM[7'h4E][27];
        newInstructionPipe = _RANDOM[7'h4E][28];
        compressInitPipe = {_RANDOM[7'h4E][31:29], _RANDOM[7'h4F][7:0]};
        compressDeqValidPipe = _RANDOM[7'h4F][8];
        groupCounterPipe = _RANDOM[7'h4F][14:9];
        compressDataReg =
          {_RANDOM[7'h4F][31:15],
           _RANDOM[7'h50],
           _RANDOM[7'h51],
           _RANDOM[7'h52],
           _RANDOM[7'h53],
           _RANDOM[7'h54],
           _RANDOM[7'h55],
           _RANDOM[7'h56],
           _RANDOM[7'h57],
           _RANDOM[7'h58],
           _RANDOM[7'h59],
           _RANDOM[7'h5A],
           _RANDOM[7'h5B],
           _RANDOM[7'h5C],
           _RANDOM[7'h5D],
           _RANDOM[7'h5E],
           _RANDOM[7'h5F][14:0]};
        compressTailValid = _RANDOM[7'h5F][15];
        compressWriteGroupCount = _RANDOM[7'h5F][21:16];
        validInputPipe = {_RANDOM[7'h5F][31:22], _RANDOM[7'h60][5:0]};
        readFromScalarPipe = {_RANDOM[7'h60][31:6], _RANDOM[7'h61][5:0]};
        ffoOutPipe = _RANDOM[7'h61][21:6];
        view__out_REG_data =
          {_RANDOM[7'h61][31:22],
           _RANDOM[7'h62],
           _RANDOM[7'h63],
           _RANDOM[7'h64],
           _RANDOM[7'h65],
           _RANDOM[7'h66],
           _RANDOM[7'h67],
           _RANDOM[7'h68],
           _RANDOM[7'h69],
           _RANDOM[7'h6A],
           _RANDOM[7'h6B],
           _RANDOM[7'h6C],
           _RANDOM[7'h6D],
           _RANDOM[7'h6E],
           _RANDOM[7'h6F],
           _RANDOM[7'h70],
           _RANDOM[7'h71][21:0]};
        view__out_REG_mask = {_RANDOM[7'h71][31:22], _RANDOM[7'h72], _RANDOM[7'h73][21:0]};
        view__out_REG_groupCounter = _RANDOM[7'h73][27:22];
        view__out_REG_ffoOutput = {_RANDOM[7'h73][31:28], _RANDOM[7'h74][11:0]};
        view__out_REG_compressValid = _RANDOM[7'h74][12];
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  assign out_data = view__out_REG_data;
  assign out_mask = view__out_REG_mask;
  assign out_groupCounter = view__out_REG_groupCounter;
  assign out_ffoOutput = view__out_REG_ffoOutput;
  assign out_compressValid = view__out_REG_compressValid;
  assign writeData = ffoIndex;
  assign stageValid = stage2Valid | in_1_valid | compressTailValid;
endmodule

