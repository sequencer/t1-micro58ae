
// Include register initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for register randomization.

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_
module LSU(
  input          clock,
                 reset,
  output         request_ready,
  input          request_valid,
  input  [2:0]   request_bits_instructionInformation_nf,
  input          request_bits_instructionInformation_mew,
  input  [1:0]   request_bits_instructionInformation_mop,
  input  [4:0]   request_bits_instructionInformation_lumop,
  input  [1:0]   request_bits_instructionInformation_eew,
  input  [4:0]   request_bits_instructionInformation_vs3,
  input          request_bits_instructionInformation_isStore,
                 request_bits_instructionInformation_maskedLoadStore,
  input  [31:0]  request_bits_rs1Data,
                 request_bits_rs2Data,
  input  [2:0]   request_bits_instructionIndex,
  input          v0UpdateVec_0_valid,
  input  [31:0]  v0UpdateVec_0_bits_data,
  input  [5:0]   v0UpdateVec_0_bits_offset,
  input  [3:0]   v0UpdateVec_0_bits_mask,
  input          v0UpdateVec_1_valid,
  input  [31:0]  v0UpdateVec_1_bits_data,
  input  [5:0]   v0UpdateVec_1_bits_offset,
  input  [3:0]   v0UpdateVec_1_bits_mask,
  input          v0UpdateVec_2_valid,
  input  [31:0]  v0UpdateVec_2_bits_data,
  input  [5:0]   v0UpdateVec_2_bits_offset,
  input  [3:0]   v0UpdateVec_2_bits_mask,
  input          v0UpdateVec_3_valid,
  input  [31:0]  v0UpdateVec_3_bits_data,
  input  [5:0]   v0UpdateVec_3_bits_offset,
  input  [3:0]   v0UpdateVec_3_bits_mask,
  input          axi4Port_aw_ready,
  output         axi4Port_aw_valid,
  output [1:0]   axi4Port_aw_bits_id,
  output [31:0]  axi4Port_aw_bits_addr,
  input          axi4Port_w_ready,
  output         axi4Port_w_valid,
  output [127:0] axi4Port_w_bits_data,
  output [15:0]  axi4Port_w_bits_strb,
  input          axi4Port_b_valid,
  input  [1:0]   axi4Port_b_bits_id,
                 axi4Port_b_bits_resp,
  input          axi4Port_ar_ready,
  output         axi4Port_ar_valid,
  output [31:0]  axi4Port_ar_bits_addr,
  output         axi4Port_r_ready,
  input          axi4Port_r_valid,
  input  [1:0]   axi4Port_r_bits_id,
  input  [127:0] axi4Port_r_bits_data,
  input  [1:0]   axi4Port_r_bits_resp,
  input          axi4Port_r_bits_last,
                 simpleAccessPorts_aw_ready,
  output         simpleAccessPorts_aw_valid,
  output [1:0]   simpleAccessPorts_aw_bits_id,
  output [31:0]  simpleAccessPorts_aw_bits_addr,
  output [2:0]   simpleAccessPorts_aw_bits_size,
  input          simpleAccessPorts_w_ready,
  output         simpleAccessPorts_w_valid,
  output [31:0]  simpleAccessPorts_w_bits_data,
  output [3:0]   simpleAccessPorts_w_bits_strb,
  input          simpleAccessPorts_b_valid,
  input  [1:0]   simpleAccessPorts_b_bits_id,
                 simpleAccessPorts_b_bits_resp,
  input          simpleAccessPorts_ar_ready,
  output         simpleAccessPorts_ar_valid,
  output [31:0]  simpleAccessPorts_ar_bits_addr,
  output         simpleAccessPorts_r_ready,
  input          simpleAccessPorts_r_valid,
  input  [1:0]   simpleAccessPorts_r_bits_id,
  input  [31:0]  simpleAccessPorts_r_bits_data,
  input  [1:0]   simpleAccessPorts_r_bits_resp,
  input          simpleAccessPorts_r_bits_last,
                 vrfReadDataPorts_0_ready,
  output         vrfReadDataPorts_0_valid,
  output [4:0]   vrfReadDataPorts_0_bits_vs,
  output [5:0]   vrfReadDataPorts_0_bits_offset,
  output [2:0]   vrfReadDataPorts_0_bits_instructionIndex,
  input          vrfReadDataPorts_1_ready,
  output         vrfReadDataPorts_1_valid,
  output [4:0]   vrfReadDataPorts_1_bits_vs,
  output [5:0]   vrfReadDataPorts_1_bits_offset,
  output [2:0]   vrfReadDataPorts_1_bits_instructionIndex,
  input          vrfReadDataPorts_2_ready,
  output         vrfReadDataPorts_2_valid,
  output [4:0]   vrfReadDataPorts_2_bits_vs,
  output [5:0]   vrfReadDataPorts_2_bits_offset,
  output [2:0]   vrfReadDataPorts_2_bits_instructionIndex,
  input          vrfReadDataPorts_3_ready,
  output         vrfReadDataPorts_3_valid,
  output [4:0]   vrfReadDataPorts_3_bits_vs,
  output [5:0]   vrfReadDataPorts_3_bits_offset,
  output [2:0]   vrfReadDataPorts_3_bits_instructionIndex,
  input          vrfReadResults_0_valid,
  input  [31:0]  vrfReadResults_0_bits,
  input          vrfReadResults_1_valid,
  input  [31:0]  vrfReadResults_1_bits,
  input          vrfReadResults_2_valid,
  input  [31:0]  vrfReadResults_2_bits,
  input          vrfReadResults_3_valid,
  input  [31:0]  vrfReadResults_3_bits,
  input          vrfWritePort_0_ready,
  output         vrfWritePort_0_valid,
  output [4:0]   vrfWritePort_0_bits_vd,
  output [5:0]   vrfWritePort_0_bits_offset,
  output [3:0]   vrfWritePort_0_bits_mask,
  output [31:0]  vrfWritePort_0_bits_data,
  output         vrfWritePort_0_bits_last,
  output [2:0]   vrfWritePort_0_bits_instructionIndex,
  input          vrfWritePort_1_ready,
  output         vrfWritePort_1_valid,
  output [4:0]   vrfWritePort_1_bits_vd,
  output [5:0]   vrfWritePort_1_bits_offset,
  output [3:0]   vrfWritePort_1_bits_mask,
  output [31:0]  vrfWritePort_1_bits_data,
  output         vrfWritePort_1_bits_last,
  output [2:0]   vrfWritePort_1_bits_instructionIndex,
  input          vrfWritePort_2_ready,
  output         vrfWritePort_2_valid,
  output [4:0]   vrfWritePort_2_bits_vd,
  output [5:0]   vrfWritePort_2_bits_offset,
  output [3:0]   vrfWritePort_2_bits_mask,
  output [31:0]  vrfWritePort_2_bits_data,
  output         vrfWritePort_2_bits_last,
  output [2:0]   vrfWritePort_2_bits_instructionIndex,
  input          vrfWritePort_3_ready,
  output         vrfWritePort_3_valid,
  output [4:0]   vrfWritePort_3_bits_vd,
  output [5:0]   vrfWritePort_3_bits_offset,
  output [3:0]   vrfWritePort_3_bits_mask,
  output [31:0]  vrfWritePort_3_bits_data,
  output         vrfWritePort_3_bits_last,
  output [2:0]   vrfWritePort_3_bits_instructionIndex,
  input          writeRelease_0,
                 writeRelease_1,
                 writeRelease_2,
                 writeRelease_3,
  output [7:0]   dataInWriteQueue_0,
                 dataInWriteQueue_1,
                 dataInWriteQueue_2,
                 dataInWriteQueue_3,
  input  [13:0]  csrInterface_vl,
                 csrInterface_vStart,
  input  [2:0]   csrInterface_vlmul,
  input  [1:0]   csrInterface_vSew,
                 csrInterface_vxrm,
  input          csrInterface_vta,
                 csrInterface_vma,
                 offsetReadResult_0_valid,
  input  [31:0]  offsetReadResult_0_bits,
  input          offsetReadResult_1_valid,
  input  [31:0]  offsetReadResult_1_bits,
  input          offsetReadResult_2_valid,
  input  [31:0]  offsetReadResult_2_bits,
  input          offsetReadResult_3_valid,
  input  [31:0]  offsetReadResult_3_bits,
  output [7:0]   lastReport,
  output [3:0]   tokenIO_offsetGroupRelease
);

  wire               _simpleDataQueue_fifo_empty;
  wire               _simpleDataQueue_fifo_full;
  wire               _simpleDataQueue_fifo_error;
  wire [77:0]        _simpleDataQueue_fifo_data_out;
  wire               _simpleSourceQueue_fifo_empty;
  wire               _simpleSourceQueue_fifo_full;
  wire               _simpleSourceQueue_fifo_error;
  wire               _dataQueue_fifo_empty;
  wire               _dataQueue_fifo_full;
  wire               _dataQueue_fifo_error;
  wire [185:0]       _dataQueue_fifo_data_out;
  wire               _sourceQueue_fifo_empty;
  wire               _sourceQueue_fifo_full;
  wire               _sourceQueue_fifo_error;
  wire               _writeIndexQueue_fifo_3_empty;
  wire               _writeIndexQueue_fifo_3_full;
  wire               _writeIndexQueue_fifo_3_error;
  wire               _writeIndexQueue_fifo_2_empty;
  wire               _writeIndexQueue_fifo_2_full;
  wire               _writeIndexQueue_fifo_2_error;
  wire               _writeIndexQueue_fifo_1_empty;
  wire               _writeIndexQueue_fifo_1_full;
  wire               _writeIndexQueue_fifo_1_error;
  wire               _writeIndexQueue_fifo_empty;
  wire               _writeIndexQueue_fifo_full;
  wire               _writeIndexQueue_fifo_error;
  wire               _otherUnitDataQueueVec_fifo_3_empty;
  wire               _otherUnitDataQueueVec_fifo_3_full;
  wire               _otherUnitDataQueueVec_fifo_3_error;
  wire [31:0]        _otherUnitDataQueueVec_fifo_3_data_out;
  wire               _otherUnitDataQueueVec_fifo_2_empty;
  wire               _otherUnitDataQueueVec_fifo_2_full;
  wire               _otherUnitDataQueueVec_fifo_2_error;
  wire [31:0]        _otherUnitDataQueueVec_fifo_2_data_out;
  wire               _otherUnitDataQueueVec_fifo_1_empty;
  wire               _otherUnitDataQueueVec_fifo_1_full;
  wire               _otherUnitDataQueueVec_fifo_1_error;
  wire [31:0]        _otherUnitDataQueueVec_fifo_1_data_out;
  wire               _otherUnitDataQueueVec_fifo_empty;
  wire               _otherUnitDataQueueVec_fifo_full;
  wire               _otherUnitDataQueueVec_fifo_error;
  wire [31:0]        _otherUnitDataQueueVec_fifo_data_out;
  wire               _otherUnitTargetQueue_fifo_empty;
  wire               _otherUnitTargetQueue_fifo_full;
  wire               _otherUnitTargetQueue_fifo_error;
  wire               _writeQueueVec_fifo_3_empty;
  wire               _writeQueueVec_fifo_3_full;
  wire               _writeQueueVec_fifo_3_error;
  wire [54:0]        _writeQueueVec_fifo_3_data_out;
  wire               _writeQueueVec_fifo_2_empty;
  wire               _writeQueueVec_fifo_2_full;
  wire               _writeQueueVec_fifo_2_error;
  wire [54:0]        _writeQueueVec_fifo_2_data_out;
  wire               _writeQueueVec_fifo_1_empty;
  wire               _writeQueueVec_fifo_1_full;
  wire               _writeQueueVec_fifo_1_error;
  wire [54:0]        _writeQueueVec_fifo_1_data_out;
  wire               _writeQueueVec_fifo_empty;
  wire               _writeQueueVec_fifo_full;
  wire               _writeQueueVec_fifo_error;
  wire [54:0]        _writeQueueVec_fifo_data_out;
  wire               _otherUnit_vrfReadDataPorts_valid;
  wire [4:0]         _otherUnit_vrfReadDataPorts_bits_vs;
  wire [5:0]         _otherUnit_vrfReadDataPorts_bits_offset;
  wire [2:0]         _otherUnit_vrfReadDataPorts_bits_instructionIndex;
  wire               _otherUnit_maskSelect_valid;
  wire [8:0]         _otherUnit_maskSelect_bits;
  wire               _otherUnit_memReadRequest_valid;
  wire               _otherUnit_memWriteRequest_valid;
  wire [7:0]         _otherUnit_memWriteRequest_bits_source;
  wire [31:0]        _otherUnit_memWriteRequest_bits_address;
  wire [1:0]         _otherUnit_memWriteRequest_bits_size;
  wire               _otherUnit_vrfWritePort_valid;
  wire [4:0]         _otherUnit_vrfWritePort_bits_vd;
  wire [5:0]         _otherUnit_vrfWritePort_bits_offset;
  wire [3:0]         _otherUnit_vrfWritePort_bits_mask;
  wire [31:0]        _otherUnit_vrfWritePort_bits_data;
  wire               _otherUnit_vrfWritePort_bits_last;
  wire [2:0]         _otherUnit_vrfWritePort_bits_instructionIndex;
  wire               _otherUnit_status_idle;
  wire               _otherUnit_status_last;
  wire [2:0]         _otherUnit_status_instructionIndex;
  wire [3:0]         _otherUnit_status_targetLane;
  wire               _otherUnit_status_isStore;
  wire               _otherUnit_offsetRelease_0;
  wire               _otherUnit_offsetRelease_1;
  wire               _otherUnit_offsetRelease_2;
  wire               _otherUnit_offsetRelease_3;
  wire               _storeUnit_maskSelect_valid;
  wire [8:0]         _storeUnit_maskSelect_bits;
  wire               _storeUnit_memRequest_valid;
  wire [9:0]         _storeUnit_memRequest_bits_index;
  wire [31:0]        _storeUnit_memRequest_bits_address;
  wire               _storeUnit_status_idle;
  wire               _storeUnit_status_last;
  wire [2:0]         _storeUnit_status_instructionIndex;
  wire [31:0]        _storeUnit_status_startAddress;
  wire [31:0]        _storeUnit_status_endAddress;
  wire               _storeUnit_vrfReadDataPorts_0_valid;
  wire [4:0]         _storeUnit_vrfReadDataPorts_0_bits_vs;
  wire [5:0]         _storeUnit_vrfReadDataPorts_0_bits_offset;
  wire [2:0]         _storeUnit_vrfReadDataPorts_0_bits_instructionIndex;
  wire               _storeUnit_vrfReadDataPorts_1_valid;
  wire [4:0]         _storeUnit_vrfReadDataPorts_1_bits_vs;
  wire [5:0]         _storeUnit_vrfReadDataPorts_1_bits_offset;
  wire [2:0]         _storeUnit_vrfReadDataPorts_1_bits_instructionIndex;
  wire               _storeUnit_vrfReadDataPorts_2_valid;
  wire [4:0]         _storeUnit_vrfReadDataPorts_2_bits_vs;
  wire [5:0]         _storeUnit_vrfReadDataPorts_2_bits_offset;
  wire [2:0]         _storeUnit_vrfReadDataPorts_2_bits_instructionIndex;
  wire               _storeUnit_vrfReadDataPorts_3_valid;
  wire [4:0]         _storeUnit_vrfReadDataPorts_3_bits_vs;
  wire [5:0]         _storeUnit_vrfReadDataPorts_3_bits_offset;
  wire [2:0]         _storeUnit_vrfReadDataPorts_3_bits_instructionIndex;
  wire               _loadUnit_maskSelect_valid;
  wire [8:0]         _loadUnit_maskSelect_bits;
  wire               _loadUnit_memRequest_valid;
  wire               _loadUnit_status_idle;
  wire               _loadUnit_status_last;
  wire [2:0]         _loadUnit_status_instructionIndex;
  wire [31:0]        _loadUnit_status_startAddress;
  wire [31:0]        _loadUnit_status_endAddress;
  wire               _loadUnit_vrfWritePort_0_valid;
  wire [4:0]         _loadUnit_vrfWritePort_0_bits_vd;
  wire [5:0]         _loadUnit_vrfWritePort_0_bits_offset;
  wire [3:0]         _loadUnit_vrfWritePort_0_bits_mask;
  wire [31:0]        _loadUnit_vrfWritePort_0_bits_data;
  wire [2:0]         _loadUnit_vrfWritePort_0_bits_instructionIndex;
  wire               _loadUnit_vrfWritePort_1_valid;
  wire [4:0]         _loadUnit_vrfWritePort_1_bits_vd;
  wire [5:0]         _loadUnit_vrfWritePort_1_bits_offset;
  wire [3:0]         _loadUnit_vrfWritePort_1_bits_mask;
  wire [31:0]        _loadUnit_vrfWritePort_1_bits_data;
  wire [2:0]         _loadUnit_vrfWritePort_1_bits_instructionIndex;
  wire               _loadUnit_vrfWritePort_2_valid;
  wire [4:0]         _loadUnit_vrfWritePort_2_bits_vd;
  wire [5:0]         _loadUnit_vrfWritePort_2_bits_offset;
  wire [3:0]         _loadUnit_vrfWritePort_2_bits_mask;
  wire [31:0]        _loadUnit_vrfWritePort_2_bits_data;
  wire [2:0]         _loadUnit_vrfWritePort_2_bits_instructionIndex;
  wire               _loadUnit_vrfWritePort_3_valid;
  wire [4:0]         _loadUnit_vrfWritePort_3_bits_vd;
  wire [5:0]         _loadUnit_vrfWritePort_3_bits_offset;
  wire [3:0]         _loadUnit_vrfWritePort_3_bits_mask;
  wire [31:0]        _loadUnit_vrfWritePort_3_bits_data;
  wire [2:0]         _loadUnit_vrfWritePort_3_bits_instructionIndex;
  wire               simpleDataQueue_almostFull;
  wire               simpleDataQueue_almostEmpty;
  wire               simpleSourceQueue_almostFull;
  wire               simpleSourceQueue_almostEmpty;
  wire               dataQueue_almostFull;
  wire               dataQueue_almostEmpty;
  wire               sourceQueue_almostFull;
  wire               sourceQueue_almostEmpty;
  wire               writeIndexQueue_3_almostFull;
  wire               writeIndexQueue_3_almostEmpty;
  wire               writeIndexQueue_2_almostFull;
  wire               writeIndexQueue_2_almostEmpty;
  wire               writeIndexQueue_1_almostFull;
  wire               writeIndexQueue_1_almostEmpty;
  wire               writeIndexQueue_almostFull;
  wire               writeIndexQueue_almostEmpty;
  wire               otherUnitDataQueueVec_3_almostFull;
  wire               otherUnitDataQueueVec_3_almostEmpty;
  wire               otherUnitDataQueueVec_2_almostFull;
  wire               otherUnitDataQueueVec_2_almostEmpty;
  wire               otherUnitDataQueueVec_1_almostFull;
  wire               otherUnitDataQueueVec_1_almostEmpty;
  wire               otherUnitDataQueueVec_0_almostFull;
  wire               otherUnitDataQueueVec_0_almostEmpty;
  wire               otherUnitTargetQueue_almostFull;
  wire               otherUnitTargetQueue_almostEmpty;
  wire               writeQueueVec_3_almostFull;
  wire               writeQueueVec_3_almostEmpty;
  wire               writeQueueVec_2_almostFull;
  wire               writeQueueVec_2_almostEmpty;
  wire               writeQueueVec_1_almostFull;
  wire               writeQueueVec_1_almostEmpty;
  wire               writeQueueVec_0_almostFull;
  wire               writeQueueVec_0_almostEmpty;
  wire [6:0]         simpleSourceQueue_enq_bits;
  wire [31:0]        simpleAccessPorts_ar_bits_addr_0;
  wire [9:0]         sourceQueue_enq_bits;
  wire [31:0]        axi4Port_ar_bits_addr_0;
  wire               request_valid_0 = request_valid;
  wire [2:0]         request_bits_instructionInformation_nf_0 = request_bits_instructionInformation_nf;
  wire               request_bits_instructionInformation_mew_0 = request_bits_instructionInformation_mew;
  wire [1:0]         request_bits_instructionInformation_mop_0 = request_bits_instructionInformation_mop;
  wire [4:0]         request_bits_instructionInformation_lumop_0 = request_bits_instructionInformation_lumop;
  wire [1:0]         request_bits_instructionInformation_eew_0 = request_bits_instructionInformation_eew;
  wire [4:0]         request_bits_instructionInformation_vs3_0 = request_bits_instructionInformation_vs3;
  wire               request_bits_instructionInformation_isStore_0 = request_bits_instructionInformation_isStore;
  wire               request_bits_instructionInformation_maskedLoadStore_0 = request_bits_instructionInformation_maskedLoadStore;
  wire [31:0]        request_bits_rs1Data_0 = request_bits_rs1Data;
  wire [31:0]        request_bits_rs2Data_0 = request_bits_rs2Data;
  wire [2:0]         request_bits_instructionIndex_0 = request_bits_instructionIndex;
  wire               axi4Port_aw_ready_0 = axi4Port_aw_ready;
  wire               axi4Port_w_ready_0 = axi4Port_w_ready;
  wire               axi4Port_b_valid_0 = axi4Port_b_valid;
  wire [1:0]         axi4Port_b_bits_id_0 = axi4Port_b_bits_id;
  wire [1:0]         axi4Port_b_bits_resp_0 = axi4Port_b_bits_resp;
  wire               axi4Port_ar_ready_0 = axi4Port_ar_ready;
  wire               axi4Port_r_valid_0 = axi4Port_r_valid;
  wire [1:0]         axi4Port_r_bits_id_0 = axi4Port_r_bits_id;
  wire [127:0]       axi4Port_r_bits_data_0 = axi4Port_r_bits_data;
  wire [1:0]         axi4Port_r_bits_resp_0 = axi4Port_r_bits_resp;
  wire               axi4Port_r_bits_last_0 = axi4Port_r_bits_last;
  wire               simpleAccessPorts_aw_ready_0 = simpleAccessPorts_aw_ready;
  wire               simpleAccessPorts_w_ready_0 = simpleAccessPorts_w_ready;
  wire               simpleAccessPorts_b_valid_0 = simpleAccessPorts_b_valid;
  wire [1:0]         simpleAccessPorts_b_bits_id_0 = simpleAccessPorts_b_bits_id;
  wire [1:0]         simpleAccessPorts_b_bits_resp_0 = simpleAccessPorts_b_bits_resp;
  wire               simpleAccessPorts_ar_ready_0 = simpleAccessPorts_ar_ready;
  wire               simpleAccessPorts_r_valid_0 = simpleAccessPorts_r_valid;
  wire [1:0]         simpleAccessPorts_r_bits_id_0 = simpleAccessPorts_r_bits_id;
  wire [31:0]        simpleAccessPorts_r_bits_data_0 = simpleAccessPorts_r_bits_data;
  wire [1:0]         simpleAccessPorts_r_bits_resp_0 = simpleAccessPorts_r_bits_resp;
  wire               simpleAccessPorts_r_bits_last_0 = simpleAccessPorts_r_bits_last;
  wire               vrfReadDataPorts_0_ready_0 = vrfReadDataPorts_0_ready;
  wire               vrfReadDataPorts_1_ready_0 = vrfReadDataPorts_1_ready;
  wire               vrfReadDataPorts_2_ready_0 = vrfReadDataPorts_2_ready;
  wire               vrfReadDataPorts_3_ready_0 = vrfReadDataPorts_3_ready;
  wire               vrfWritePort_0_ready_0 = vrfWritePort_0_ready;
  wire               vrfWritePort_1_ready_0 = vrfWritePort_1_ready;
  wire               vrfWritePort_2_ready_0 = vrfWritePort_2_ready;
  wire               vrfWritePort_3_ready_0 = vrfWritePort_3_ready;
  wire [31:0]        otherUnitDataQueueVec_0_enq_bits = vrfReadResults_0_bits;
  wire [31:0]        otherUnitDataQueueVec_1_enq_bits = vrfReadResults_1_bits;
  wire [31:0]        otherUnitDataQueueVec_2_enq_bits = vrfReadResults_2_bits;
  wire [31:0]        otherUnitDataQueueVec_3_enq_bits = vrfReadResults_3_bits;
  wire               writeIndexQueue_deq_ready = writeRelease_0;
  wire               writeIndexQueue_1_deq_ready = writeRelease_1;
  wire               writeIndexQueue_2_deq_ready = writeRelease_2;
  wire               writeIndexQueue_3_deq_ready = writeRelease_3;
  wire [1:0]         vrfReadDataPorts_0_bits_readSource = 2'h2;
  wire [1:0]         vrfReadDataPorts_1_bits_readSource = 2'h2;
  wire [1:0]         vrfReadDataPorts_2_bits_readSource = 2'h2;
  wire [1:0]         vrfReadDataPorts_3_bits_readSource = 2'h2;
  wire [1:0]         axi4Port_ar_bits_id = 2'h0;
  wire [1:0]         simpleAccessPorts_ar_bits_id = 2'h0;
  wire [1:0]         axi4Port_aw_bits_burst = 2'h1;
  wire [1:0]         axi4Port_ar_bits_burst = 2'h1;
  wire [1:0]         simpleAccessPorts_aw_bits_burst = 2'h1;
  wire [1:0]         simpleAccessPorts_ar_bits_burst = 2'h1;
  wire [3:0]         writeQueueVec_0_enq_bits_targetLane = 4'h1;
  wire [3:0]         writeQueueVec_1_enq_bits_targetLane = 4'h2;
  wire [3:0]         writeQueueVec_2_enq_bits_targetLane = 4'h4;
  wire [3:0]         writeQueueVec_3_enq_bits_targetLane = 4'h8;
  wire [7:0]         axi4Port_aw_bits_len = 8'h0;
  wire [7:0]         axi4Port_ar_bits_len = 8'h0;
  wire [7:0]         simpleAccessPorts_aw_bits_len = 8'h0;
  wire [7:0]         simpleAccessPorts_ar_bits_len = 8'h0;
  wire [2:0]         axi4Port_aw_bits_size = 3'h4;
  wire [2:0]         axi4Port_ar_bits_size = 3'h4;
  wire               axi4Port_aw_bits_lock = 1'h0;
  wire               axi4Port_ar_bits_lock = 1'h0;
  wire               simpleAccessPorts_aw_bits_lock = 1'h0;
  wire               simpleAccessPorts_ar_bits_lock = 1'h0;
  wire [3:0]         axi4Port_aw_bits_cache = 4'h0;
  wire [3:0]         axi4Port_aw_bits_qos = 4'h0;
  wire [3:0]         axi4Port_aw_bits_region = 4'h0;
  wire [3:0]         axi4Port_ar_bits_cache = 4'h0;
  wire [3:0]         axi4Port_ar_bits_qos = 4'h0;
  wire [3:0]         axi4Port_ar_bits_region = 4'h0;
  wire [3:0]         simpleAccessPorts_aw_bits_cache = 4'h0;
  wire [3:0]         simpleAccessPorts_aw_bits_qos = 4'h0;
  wire [3:0]         simpleAccessPorts_aw_bits_region = 4'h0;
  wire [3:0]         simpleAccessPorts_ar_bits_cache = 4'h0;
  wire [3:0]         simpleAccessPorts_ar_bits_qos = 4'h0;
  wire [3:0]         simpleAccessPorts_ar_bits_region = 4'h0;
  wire [2:0]         axi4Port_aw_bits_prot = 3'h0;
  wire [2:0]         axi4Port_ar_bits_prot = 3'h0;
  wire [2:0]         simpleAccessPorts_aw_bits_prot = 3'h0;
  wire [2:0]         simpleAccessPorts_ar_bits_prot = 3'h0;
  wire               axi4Port_w_bits_last = 1'h1;
  wire               axi4Port_b_ready = 1'h1;
  wire               simpleAccessPorts_w_bits_last = 1'h1;
  wire               simpleAccessPorts_b_ready = 1'h1;
  wire [2:0]         simpleAccessPorts_ar_bits_size = 3'h2;
  wire               dataQueue_deq_ready = axi4Port_w_ready_0;
  wire               dataQueue_deq_valid;
  wire [127:0]       dataQueue_deq_bits_data;
  wire [15:0]        dataQueue_deq_bits_mask;
  wire               simpleDataQueue_deq_ready = simpleAccessPorts_w_ready_0;
  wire               simpleDataQueue_deq_valid;
  wire [31:0]        simpleDataQueue_deq_bits_data;
  wire [3:0]         simpleDataQueue_deq_bits_mask;
  wire               writeQueueVec_0_deq_ready = vrfWritePort_0_ready_0;
  wire               writeQueueVec_0_deq_valid;
  wire [4:0]         writeQueueVec_0_deq_bits_data_vd;
  wire [5:0]         writeQueueVec_0_deq_bits_data_offset;
  wire [3:0]         writeQueueVec_0_deq_bits_data_mask;
  wire [31:0]        writeQueueVec_0_deq_bits_data_data;
  wire               writeQueueVec_0_deq_bits_data_last;
  wire [2:0]         writeQueueVec_0_deq_bits_data_instructionIndex;
  wire               writeQueueVec_1_deq_ready = vrfWritePort_1_ready_0;
  wire               writeQueueVec_1_deq_valid;
  wire [4:0]         writeQueueVec_1_deq_bits_data_vd;
  wire [5:0]         writeQueueVec_1_deq_bits_data_offset;
  wire [3:0]         writeQueueVec_1_deq_bits_data_mask;
  wire [31:0]        writeQueueVec_1_deq_bits_data_data;
  wire               writeQueueVec_1_deq_bits_data_last;
  wire [2:0]         writeQueueVec_1_deq_bits_data_instructionIndex;
  wire               writeQueueVec_2_deq_ready = vrfWritePort_2_ready_0;
  wire               writeQueueVec_2_deq_valid;
  wire [4:0]         writeQueueVec_2_deq_bits_data_vd;
  wire [5:0]         writeQueueVec_2_deq_bits_data_offset;
  wire [3:0]         writeQueueVec_2_deq_bits_data_mask;
  wire [31:0]        writeQueueVec_2_deq_bits_data_data;
  wire               writeQueueVec_2_deq_bits_data_last;
  wire [2:0]         writeQueueVec_2_deq_bits_data_instructionIndex;
  wire               writeQueueVec_3_deq_ready = vrfWritePort_3_ready_0;
  wire               writeQueueVec_3_deq_valid;
  wire [4:0]         writeQueueVec_3_deq_bits_data_vd;
  wire [5:0]         writeQueueVec_3_deq_bits_data_offset;
  wire [3:0]         writeQueueVec_3_deq_bits_data_mask;
  wire [31:0]        writeQueueVec_3_deq_bits_data_data;
  wire               writeQueueVec_3_deq_bits_data_last;
  wire [2:0]         writeQueueVec_3_deq_bits_data_instructionIndex;
  reg  [31:0]        v0_0;
  reg  [31:0]        v0_1;
  reg  [31:0]        v0_2;
  reg  [31:0]        v0_3;
  reg  [31:0]        v0_4;
  reg  [31:0]        v0_5;
  reg  [31:0]        v0_6;
  reg  [31:0]        v0_7;
  reg  [31:0]        v0_8;
  reg  [31:0]        v0_9;
  reg  [31:0]        v0_10;
  reg  [31:0]        v0_11;
  reg  [31:0]        v0_12;
  reg  [31:0]        v0_13;
  reg  [31:0]        v0_14;
  reg  [31:0]        v0_15;
  reg  [31:0]        v0_16;
  reg  [31:0]        v0_17;
  reg  [31:0]        v0_18;
  reg  [31:0]        v0_19;
  reg  [31:0]        v0_20;
  reg  [31:0]        v0_21;
  reg  [31:0]        v0_22;
  reg  [31:0]        v0_23;
  reg  [31:0]        v0_24;
  reg  [31:0]        v0_25;
  reg  [31:0]        v0_26;
  reg  [31:0]        v0_27;
  reg  [31:0]        v0_28;
  reg  [31:0]        v0_29;
  reg  [31:0]        v0_30;
  reg  [31:0]        v0_31;
  reg  [31:0]        v0_32;
  reg  [31:0]        v0_33;
  reg  [31:0]        v0_34;
  reg  [31:0]        v0_35;
  reg  [31:0]        v0_36;
  reg  [31:0]        v0_37;
  reg  [31:0]        v0_38;
  reg  [31:0]        v0_39;
  reg  [31:0]        v0_40;
  reg  [31:0]        v0_41;
  reg  [31:0]        v0_42;
  reg  [31:0]        v0_43;
  reg  [31:0]        v0_44;
  reg  [31:0]        v0_45;
  reg  [31:0]        v0_46;
  reg  [31:0]        v0_47;
  reg  [31:0]        v0_48;
  reg  [31:0]        v0_49;
  reg  [31:0]        v0_50;
  reg  [31:0]        v0_51;
  reg  [31:0]        v0_52;
  reg  [31:0]        v0_53;
  reg  [31:0]        v0_54;
  reg  [31:0]        v0_55;
  reg  [31:0]        v0_56;
  reg  [31:0]        v0_57;
  reg  [31:0]        v0_58;
  reg  [31:0]        v0_59;
  reg  [31:0]        v0_60;
  reg  [31:0]        v0_61;
  reg  [31:0]        v0_62;
  reg  [31:0]        v0_63;
  reg  [31:0]        v0_64;
  reg  [31:0]        v0_65;
  reg  [31:0]        v0_66;
  reg  [31:0]        v0_67;
  reg  [31:0]        v0_68;
  reg  [31:0]        v0_69;
  reg  [31:0]        v0_70;
  reg  [31:0]        v0_71;
  reg  [31:0]        v0_72;
  reg  [31:0]        v0_73;
  reg  [31:0]        v0_74;
  reg  [31:0]        v0_75;
  reg  [31:0]        v0_76;
  reg  [31:0]        v0_77;
  reg  [31:0]        v0_78;
  reg  [31:0]        v0_79;
  reg  [31:0]        v0_80;
  reg  [31:0]        v0_81;
  reg  [31:0]        v0_82;
  reg  [31:0]        v0_83;
  reg  [31:0]        v0_84;
  reg  [31:0]        v0_85;
  reg  [31:0]        v0_86;
  reg  [31:0]        v0_87;
  reg  [31:0]        v0_88;
  reg  [31:0]        v0_89;
  reg  [31:0]        v0_90;
  reg  [31:0]        v0_91;
  reg  [31:0]        v0_92;
  reg  [31:0]        v0_93;
  reg  [31:0]        v0_94;
  reg  [31:0]        v0_95;
  reg  [31:0]        v0_96;
  reg  [31:0]        v0_97;
  reg  [31:0]        v0_98;
  reg  [31:0]        v0_99;
  reg  [31:0]        v0_100;
  reg  [31:0]        v0_101;
  reg  [31:0]        v0_102;
  reg  [31:0]        v0_103;
  reg  [31:0]        v0_104;
  reg  [31:0]        v0_105;
  reg  [31:0]        v0_106;
  reg  [31:0]        v0_107;
  reg  [31:0]        v0_108;
  reg  [31:0]        v0_109;
  reg  [31:0]        v0_110;
  reg  [31:0]        v0_111;
  reg  [31:0]        v0_112;
  reg  [31:0]        v0_113;
  reg  [31:0]        v0_114;
  reg  [31:0]        v0_115;
  reg  [31:0]        v0_116;
  reg  [31:0]        v0_117;
  reg  [31:0]        v0_118;
  reg  [31:0]        v0_119;
  reg  [31:0]        v0_120;
  reg  [31:0]        v0_121;
  reg  [31:0]        v0_122;
  reg  [31:0]        v0_123;
  reg  [31:0]        v0_124;
  reg  [31:0]        v0_125;
  reg  [31:0]        v0_126;
  reg  [31:0]        v0_127;
  reg  [31:0]        v0_128;
  reg  [31:0]        v0_129;
  reg  [31:0]        v0_130;
  reg  [31:0]        v0_131;
  reg  [31:0]        v0_132;
  reg  [31:0]        v0_133;
  reg  [31:0]        v0_134;
  reg  [31:0]        v0_135;
  reg  [31:0]        v0_136;
  reg  [31:0]        v0_137;
  reg  [31:0]        v0_138;
  reg  [31:0]        v0_139;
  reg  [31:0]        v0_140;
  reg  [31:0]        v0_141;
  reg  [31:0]        v0_142;
  reg  [31:0]        v0_143;
  reg  [31:0]        v0_144;
  reg  [31:0]        v0_145;
  reg  [31:0]        v0_146;
  reg  [31:0]        v0_147;
  reg  [31:0]        v0_148;
  reg  [31:0]        v0_149;
  reg  [31:0]        v0_150;
  reg  [31:0]        v0_151;
  reg  [31:0]        v0_152;
  reg  [31:0]        v0_153;
  reg  [31:0]        v0_154;
  reg  [31:0]        v0_155;
  reg  [31:0]        v0_156;
  reg  [31:0]        v0_157;
  reg  [31:0]        v0_158;
  reg  [31:0]        v0_159;
  reg  [31:0]        v0_160;
  reg  [31:0]        v0_161;
  reg  [31:0]        v0_162;
  reg  [31:0]        v0_163;
  reg  [31:0]        v0_164;
  reg  [31:0]        v0_165;
  reg  [31:0]        v0_166;
  reg  [31:0]        v0_167;
  reg  [31:0]        v0_168;
  reg  [31:0]        v0_169;
  reg  [31:0]        v0_170;
  reg  [31:0]        v0_171;
  reg  [31:0]        v0_172;
  reg  [31:0]        v0_173;
  reg  [31:0]        v0_174;
  reg  [31:0]        v0_175;
  reg  [31:0]        v0_176;
  reg  [31:0]        v0_177;
  reg  [31:0]        v0_178;
  reg  [31:0]        v0_179;
  reg  [31:0]        v0_180;
  reg  [31:0]        v0_181;
  reg  [31:0]        v0_182;
  reg  [31:0]        v0_183;
  reg  [31:0]        v0_184;
  reg  [31:0]        v0_185;
  reg  [31:0]        v0_186;
  reg  [31:0]        v0_187;
  reg  [31:0]        v0_188;
  reg  [31:0]        v0_189;
  reg  [31:0]        v0_190;
  reg  [31:0]        v0_191;
  reg  [31:0]        v0_192;
  reg  [31:0]        v0_193;
  reg  [31:0]        v0_194;
  reg  [31:0]        v0_195;
  reg  [31:0]        v0_196;
  reg  [31:0]        v0_197;
  reg  [31:0]        v0_198;
  reg  [31:0]        v0_199;
  reg  [31:0]        v0_200;
  reg  [31:0]        v0_201;
  reg  [31:0]        v0_202;
  reg  [31:0]        v0_203;
  reg  [31:0]        v0_204;
  reg  [31:0]        v0_205;
  reg  [31:0]        v0_206;
  reg  [31:0]        v0_207;
  reg  [31:0]        v0_208;
  reg  [31:0]        v0_209;
  reg  [31:0]        v0_210;
  reg  [31:0]        v0_211;
  reg  [31:0]        v0_212;
  reg  [31:0]        v0_213;
  reg  [31:0]        v0_214;
  reg  [31:0]        v0_215;
  reg  [31:0]        v0_216;
  reg  [31:0]        v0_217;
  reg  [31:0]        v0_218;
  reg  [31:0]        v0_219;
  reg  [31:0]        v0_220;
  reg  [31:0]        v0_221;
  reg  [31:0]        v0_222;
  reg  [31:0]        v0_223;
  reg  [31:0]        v0_224;
  reg  [31:0]        v0_225;
  reg  [31:0]        v0_226;
  reg  [31:0]        v0_227;
  reg  [31:0]        v0_228;
  reg  [31:0]        v0_229;
  reg  [31:0]        v0_230;
  reg  [31:0]        v0_231;
  reg  [31:0]        v0_232;
  reg  [31:0]        v0_233;
  reg  [31:0]        v0_234;
  reg  [31:0]        v0_235;
  reg  [31:0]        v0_236;
  reg  [31:0]        v0_237;
  reg  [31:0]        v0_238;
  reg  [31:0]        v0_239;
  reg  [31:0]        v0_240;
  reg  [31:0]        v0_241;
  reg  [31:0]        v0_242;
  reg  [31:0]        v0_243;
  reg  [31:0]        v0_244;
  reg  [31:0]        v0_245;
  reg  [31:0]        v0_246;
  reg  [31:0]        v0_247;
  reg  [31:0]        v0_248;
  reg  [31:0]        v0_249;
  reg  [31:0]        v0_250;
  reg  [31:0]        v0_251;
  reg  [31:0]        v0_252;
  reg  [31:0]        v0_253;
  reg  [31:0]        v0_254;
  reg  [31:0]        v0_255;
  wire [15:0]        maskExt_lo = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt = {maskExt_hi, maskExt_lo};
  wire [15:0]        maskExt_lo_1 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_1 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_1 = {maskExt_hi_1, maskExt_lo_1};
  wire [15:0]        maskExt_lo_2 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_2 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_2 = {maskExt_hi_2, maskExt_lo_2};
  wire [15:0]        maskExt_lo_3 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_3 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_3 = {maskExt_hi_3, maskExt_lo_3};
  wire [15:0]        maskExt_lo_4 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_4 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_4 = {maskExt_hi_4, maskExt_lo_4};
  wire [15:0]        maskExt_lo_5 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_5 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_5 = {maskExt_hi_5, maskExt_lo_5};
  wire [15:0]        maskExt_lo_6 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_6 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_6 = {maskExt_hi_6, maskExt_lo_6};
  wire [15:0]        maskExt_lo_7 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_7 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_7 = {maskExt_hi_7, maskExt_lo_7};
  wire [15:0]        maskExt_lo_8 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_8 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_8 = {maskExt_hi_8, maskExt_lo_8};
  wire [15:0]        maskExt_lo_9 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_9 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_9 = {maskExt_hi_9, maskExt_lo_9};
  wire [15:0]        maskExt_lo_10 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_10 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_10 = {maskExt_hi_10, maskExt_lo_10};
  wire [15:0]        maskExt_lo_11 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_11 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_11 = {maskExt_hi_11, maskExt_lo_11};
  wire [15:0]        maskExt_lo_12 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_12 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_12 = {maskExt_hi_12, maskExt_lo_12};
  wire [15:0]        maskExt_lo_13 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_13 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_13 = {maskExt_hi_13, maskExt_lo_13};
  wire [15:0]        maskExt_lo_14 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_14 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_14 = {maskExt_hi_14, maskExt_lo_14};
  wire [15:0]        maskExt_lo_15 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_15 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_15 = {maskExt_hi_15, maskExt_lo_15};
  wire [15:0]        maskExt_lo_16 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_16 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_16 = {maskExt_hi_16, maskExt_lo_16};
  wire [15:0]        maskExt_lo_17 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_17 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_17 = {maskExt_hi_17, maskExt_lo_17};
  wire [15:0]        maskExt_lo_18 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_18 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_18 = {maskExt_hi_18, maskExt_lo_18};
  wire [15:0]        maskExt_lo_19 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_19 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_19 = {maskExt_hi_19, maskExt_lo_19};
  wire [15:0]        maskExt_lo_20 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_20 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_20 = {maskExt_hi_20, maskExt_lo_20};
  wire [15:0]        maskExt_lo_21 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_21 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_21 = {maskExt_hi_21, maskExt_lo_21};
  wire [15:0]        maskExt_lo_22 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_22 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_22 = {maskExt_hi_22, maskExt_lo_22};
  wire [15:0]        maskExt_lo_23 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_23 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_23 = {maskExt_hi_23, maskExt_lo_23};
  wire [15:0]        maskExt_lo_24 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_24 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_24 = {maskExt_hi_24, maskExt_lo_24};
  wire [15:0]        maskExt_lo_25 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_25 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_25 = {maskExt_hi_25, maskExt_lo_25};
  wire [15:0]        maskExt_lo_26 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_26 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_26 = {maskExt_hi_26, maskExt_lo_26};
  wire [15:0]        maskExt_lo_27 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_27 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_27 = {maskExt_hi_27, maskExt_lo_27};
  wire [15:0]        maskExt_lo_28 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_28 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_28 = {maskExt_hi_28, maskExt_lo_28};
  wire [15:0]        maskExt_lo_29 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_29 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_29 = {maskExt_hi_29, maskExt_lo_29};
  wire [15:0]        maskExt_lo_30 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_30 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_30 = {maskExt_hi_30, maskExt_lo_30};
  wire [15:0]        maskExt_lo_31 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_31 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_31 = {maskExt_hi_31, maskExt_lo_31};
  wire [15:0]        maskExt_lo_32 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_32 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_32 = {maskExt_hi_32, maskExt_lo_32};
  wire [15:0]        maskExt_lo_33 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_33 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_33 = {maskExt_hi_33, maskExt_lo_33};
  wire [15:0]        maskExt_lo_34 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_34 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_34 = {maskExt_hi_34, maskExt_lo_34};
  wire [15:0]        maskExt_lo_35 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_35 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_35 = {maskExt_hi_35, maskExt_lo_35};
  wire [15:0]        maskExt_lo_36 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_36 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_36 = {maskExt_hi_36, maskExt_lo_36};
  wire [15:0]        maskExt_lo_37 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_37 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_37 = {maskExt_hi_37, maskExt_lo_37};
  wire [15:0]        maskExt_lo_38 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_38 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_38 = {maskExt_hi_38, maskExt_lo_38};
  wire [15:0]        maskExt_lo_39 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_39 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_39 = {maskExt_hi_39, maskExt_lo_39};
  wire [15:0]        maskExt_lo_40 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_40 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_40 = {maskExt_hi_40, maskExt_lo_40};
  wire [15:0]        maskExt_lo_41 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_41 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_41 = {maskExt_hi_41, maskExt_lo_41};
  wire [15:0]        maskExt_lo_42 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_42 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_42 = {maskExt_hi_42, maskExt_lo_42};
  wire [15:0]        maskExt_lo_43 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_43 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_43 = {maskExt_hi_43, maskExt_lo_43};
  wire [15:0]        maskExt_lo_44 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_44 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_44 = {maskExt_hi_44, maskExt_lo_44};
  wire [15:0]        maskExt_lo_45 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_45 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_45 = {maskExt_hi_45, maskExt_lo_45};
  wire [15:0]        maskExt_lo_46 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_46 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_46 = {maskExt_hi_46, maskExt_lo_46};
  wire [15:0]        maskExt_lo_47 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_47 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_47 = {maskExt_hi_47, maskExt_lo_47};
  wire [15:0]        maskExt_lo_48 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_48 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_48 = {maskExt_hi_48, maskExt_lo_48};
  wire [15:0]        maskExt_lo_49 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_49 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_49 = {maskExt_hi_49, maskExt_lo_49};
  wire [15:0]        maskExt_lo_50 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_50 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_50 = {maskExt_hi_50, maskExt_lo_50};
  wire [15:0]        maskExt_lo_51 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_51 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_51 = {maskExt_hi_51, maskExt_lo_51};
  wire [15:0]        maskExt_lo_52 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_52 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_52 = {maskExt_hi_52, maskExt_lo_52};
  wire [15:0]        maskExt_lo_53 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_53 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_53 = {maskExt_hi_53, maskExt_lo_53};
  wire [15:0]        maskExt_lo_54 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_54 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_54 = {maskExt_hi_54, maskExt_lo_54};
  wire [15:0]        maskExt_lo_55 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_55 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_55 = {maskExt_hi_55, maskExt_lo_55};
  wire [15:0]        maskExt_lo_56 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_56 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_56 = {maskExt_hi_56, maskExt_lo_56};
  wire [15:0]        maskExt_lo_57 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_57 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_57 = {maskExt_hi_57, maskExt_lo_57};
  wire [15:0]        maskExt_lo_58 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_58 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_58 = {maskExt_hi_58, maskExt_lo_58};
  wire [15:0]        maskExt_lo_59 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_59 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_59 = {maskExt_hi_59, maskExt_lo_59};
  wire [15:0]        maskExt_lo_60 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_60 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_60 = {maskExt_hi_60, maskExt_lo_60};
  wire [15:0]        maskExt_lo_61 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_61 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_61 = {maskExt_hi_61, maskExt_lo_61};
  wire [15:0]        maskExt_lo_62 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_62 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_62 = {maskExt_hi_62, maskExt_lo_62};
  wire [15:0]        maskExt_lo_63 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_63 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_63 = {maskExt_hi_63, maskExt_lo_63};
  wire [15:0]        maskExt_lo_64 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_64 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_64 = {maskExt_hi_64, maskExt_lo_64};
  wire [15:0]        maskExt_lo_65 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_65 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_65 = {maskExt_hi_65, maskExt_lo_65};
  wire [15:0]        maskExt_lo_66 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_66 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_66 = {maskExt_hi_66, maskExt_lo_66};
  wire [15:0]        maskExt_lo_67 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_67 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_67 = {maskExt_hi_67, maskExt_lo_67};
  wire [15:0]        maskExt_lo_68 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_68 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_68 = {maskExt_hi_68, maskExt_lo_68};
  wire [15:0]        maskExt_lo_69 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_69 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_69 = {maskExt_hi_69, maskExt_lo_69};
  wire [15:0]        maskExt_lo_70 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_70 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_70 = {maskExt_hi_70, maskExt_lo_70};
  wire [15:0]        maskExt_lo_71 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_71 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_71 = {maskExt_hi_71, maskExt_lo_71};
  wire [15:0]        maskExt_lo_72 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_72 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_72 = {maskExt_hi_72, maskExt_lo_72};
  wire [15:0]        maskExt_lo_73 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_73 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_73 = {maskExt_hi_73, maskExt_lo_73};
  wire [15:0]        maskExt_lo_74 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_74 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_74 = {maskExt_hi_74, maskExt_lo_74};
  wire [15:0]        maskExt_lo_75 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_75 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_75 = {maskExt_hi_75, maskExt_lo_75};
  wire [15:0]        maskExt_lo_76 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_76 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_76 = {maskExt_hi_76, maskExt_lo_76};
  wire [15:0]        maskExt_lo_77 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_77 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_77 = {maskExt_hi_77, maskExt_lo_77};
  wire [15:0]        maskExt_lo_78 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_78 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_78 = {maskExt_hi_78, maskExt_lo_78};
  wire [15:0]        maskExt_lo_79 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_79 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_79 = {maskExt_hi_79, maskExt_lo_79};
  wire [15:0]        maskExt_lo_80 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_80 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_80 = {maskExt_hi_80, maskExt_lo_80};
  wire [15:0]        maskExt_lo_81 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_81 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_81 = {maskExt_hi_81, maskExt_lo_81};
  wire [15:0]        maskExt_lo_82 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_82 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_82 = {maskExt_hi_82, maskExt_lo_82};
  wire [15:0]        maskExt_lo_83 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_83 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_83 = {maskExt_hi_83, maskExt_lo_83};
  wire [15:0]        maskExt_lo_84 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_84 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_84 = {maskExt_hi_84, maskExt_lo_84};
  wire [15:0]        maskExt_lo_85 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_85 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_85 = {maskExt_hi_85, maskExt_lo_85};
  wire [15:0]        maskExt_lo_86 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_86 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_86 = {maskExt_hi_86, maskExt_lo_86};
  wire [15:0]        maskExt_lo_87 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_87 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_87 = {maskExt_hi_87, maskExt_lo_87};
  wire [15:0]        maskExt_lo_88 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_88 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_88 = {maskExt_hi_88, maskExt_lo_88};
  wire [15:0]        maskExt_lo_89 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_89 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_89 = {maskExt_hi_89, maskExt_lo_89};
  wire [15:0]        maskExt_lo_90 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_90 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_90 = {maskExt_hi_90, maskExt_lo_90};
  wire [15:0]        maskExt_lo_91 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_91 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_91 = {maskExt_hi_91, maskExt_lo_91};
  wire [15:0]        maskExt_lo_92 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_92 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_92 = {maskExt_hi_92, maskExt_lo_92};
  wire [15:0]        maskExt_lo_93 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_93 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_93 = {maskExt_hi_93, maskExt_lo_93};
  wire [15:0]        maskExt_lo_94 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_94 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_94 = {maskExt_hi_94, maskExt_lo_94};
  wire [15:0]        maskExt_lo_95 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_95 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_95 = {maskExt_hi_95, maskExt_lo_95};
  wire [15:0]        maskExt_lo_96 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_96 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_96 = {maskExt_hi_96, maskExt_lo_96};
  wire [15:0]        maskExt_lo_97 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_97 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_97 = {maskExt_hi_97, maskExt_lo_97};
  wire [15:0]        maskExt_lo_98 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_98 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_98 = {maskExt_hi_98, maskExt_lo_98};
  wire [15:0]        maskExt_lo_99 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_99 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_99 = {maskExt_hi_99, maskExt_lo_99};
  wire [15:0]        maskExt_lo_100 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_100 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_100 = {maskExt_hi_100, maskExt_lo_100};
  wire [15:0]        maskExt_lo_101 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_101 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_101 = {maskExt_hi_101, maskExt_lo_101};
  wire [15:0]        maskExt_lo_102 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_102 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_102 = {maskExt_hi_102, maskExt_lo_102};
  wire [15:0]        maskExt_lo_103 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_103 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_103 = {maskExt_hi_103, maskExt_lo_103};
  wire [15:0]        maskExt_lo_104 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_104 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_104 = {maskExt_hi_104, maskExt_lo_104};
  wire [15:0]        maskExt_lo_105 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_105 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_105 = {maskExt_hi_105, maskExt_lo_105};
  wire [15:0]        maskExt_lo_106 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_106 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_106 = {maskExt_hi_106, maskExt_lo_106};
  wire [15:0]        maskExt_lo_107 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_107 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_107 = {maskExt_hi_107, maskExt_lo_107};
  wire [15:0]        maskExt_lo_108 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_108 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_108 = {maskExt_hi_108, maskExt_lo_108};
  wire [15:0]        maskExt_lo_109 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_109 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_109 = {maskExt_hi_109, maskExt_lo_109};
  wire [15:0]        maskExt_lo_110 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_110 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_110 = {maskExt_hi_110, maskExt_lo_110};
  wire [15:0]        maskExt_lo_111 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_111 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_111 = {maskExt_hi_111, maskExt_lo_111};
  wire [15:0]        maskExt_lo_112 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_112 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_112 = {maskExt_hi_112, maskExt_lo_112};
  wire [15:0]        maskExt_lo_113 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_113 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_113 = {maskExt_hi_113, maskExt_lo_113};
  wire [15:0]        maskExt_lo_114 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_114 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_114 = {maskExt_hi_114, maskExt_lo_114};
  wire [15:0]        maskExt_lo_115 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_115 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_115 = {maskExt_hi_115, maskExt_lo_115};
  wire [15:0]        maskExt_lo_116 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_116 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_116 = {maskExt_hi_116, maskExt_lo_116};
  wire [15:0]        maskExt_lo_117 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_117 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_117 = {maskExt_hi_117, maskExt_lo_117};
  wire [15:0]        maskExt_lo_118 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_118 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_118 = {maskExt_hi_118, maskExt_lo_118};
  wire [15:0]        maskExt_lo_119 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_119 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_119 = {maskExt_hi_119, maskExt_lo_119};
  wire [15:0]        maskExt_lo_120 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_120 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_120 = {maskExt_hi_120, maskExt_lo_120};
  wire [15:0]        maskExt_lo_121 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_121 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_121 = {maskExt_hi_121, maskExt_lo_121};
  wire [15:0]        maskExt_lo_122 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_122 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_122 = {maskExt_hi_122, maskExt_lo_122};
  wire [15:0]        maskExt_lo_123 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_123 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_123 = {maskExt_hi_123, maskExt_lo_123};
  wire [15:0]        maskExt_lo_124 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_124 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_124 = {maskExt_hi_124, maskExt_lo_124};
  wire [15:0]        maskExt_lo_125 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_125 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_125 = {maskExt_hi_125, maskExt_lo_125};
  wire [15:0]        maskExt_lo_126 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_126 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_126 = {maskExt_hi_126, maskExt_lo_126};
  wire [15:0]        maskExt_lo_127 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_127 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_127 = {maskExt_hi_127, maskExt_lo_127};
  wire [15:0]        maskExt_lo_128 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_128 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_128 = {maskExt_hi_128, maskExt_lo_128};
  wire [15:0]        maskExt_lo_129 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_129 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_129 = {maskExt_hi_129, maskExt_lo_129};
  wire [15:0]        maskExt_lo_130 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_130 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_130 = {maskExt_hi_130, maskExt_lo_130};
  wire [15:0]        maskExt_lo_131 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_131 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_131 = {maskExt_hi_131, maskExt_lo_131};
  wire [15:0]        maskExt_lo_132 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_132 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_132 = {maskExt_hi_132, maskExt_lo_132};
  wire [15:0]        maskExt_lo_133 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_133 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_133 = {maskExt_hi_133, maskExt_lo_133};
  wire [15:0]        maskExt_lo_134 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_134 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_134 = {maskExt_hi_134, maskExt_lo_134};
  wire [15:0]        maskExt_lo_135 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_135 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_135 = {maskExt_hi_135, maskExt_lo_135};
  wire [15:0]        maskExt_lo_136 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_136 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_136 = {maskExt_hi_136, maskExt_lo_136};
  wire [15:0]        maskExt_lo_137 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_137 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_137 = {maskExt_hi_137, maskExt_lo_137};
  wire [15:0]        maskExt_lo_138 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_138 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_138 = {maskExt_hi_138, maskExt_lo_138};
  wire [15:0]        maskExt_lo_139 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_139 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_139 = {maskExt_hi_139, maskExt_lo_139};
  wire [15:0]        maskExt_lo_140 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_140 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_140 = {maskExt_hi_140, maskExt_lo_140};
  wire [15:0]        maskExt_lo_141 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_141 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_141 = {maskExt_hi_141, maskExt_lo_141};
  wire [15:0]        maskExt_lo_142 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_142 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_142 = {maskExt_hi_142, maskExt_lo_142};
  wire [15:0]        maskExt_lo_143 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_143 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_143 = {maskExt_hi_143, maskExt_lo_143};
  wire [15:0]        maskExt_lo_144 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_144 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_144 = {maskExt_hi_144, maskExt_lo_144};
  wire [15:0]        maskExt_lo_145 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_145 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_145 = {maskExt_hi_145, maskExt_lo_145};
  wire [15:0]        maskExt_lo_146 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_146 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_146 = {maskExt_hi_146, maskExt_lo_146};
  wire [15:0]        maskExt_lo_147 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_147 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_147 = {maskExt_hi_147, maskExt_lo_147};
  wire [15:0]        maskExt_lo_148 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_148 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_148 = {maskExt_hi_148, maskExt_lo_148};
  wire [15:0]        maskExt_lo_149 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_149 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_149 = {maskExt_hi_149, maskExt_lo_149};
  wire [15:0]        maskExt_lo_150 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_150 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_150 = {maskExt_hi_150, maskExt_lo_150};
  wire [15:0]        maskExt_lo_151 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_151 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_151 = {maskExt_hi_151, maskExt_lo_151};
  wire [15:0]        maskExt_lo_152 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_152 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_152 = {maskExt_hi_152, maskExt_lo_152};
  wire [15:0]        maskExt_lo_153 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_153 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_153 = {maskExt_hi_153, maskExt_lo_153};
  wire [15:0]        maskExt_lo_154 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_154 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_154 = {maskExt_hi_154, maskExt_lo_154};
  wire [15:0]        maskExt_lo_155 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_155 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_155 = {maskExt_hi_155, maskExt_lo_155};
  wire [15:0]        maskExt_lo_156 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_156 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_156 = {maskExt_hi_156, maskExt_lo_156};
  wire [15:0]        maskExt_lo_157 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_157 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_157 = {maskExt_hi_157, maskExt_lo_157};
  wire [15:0]        maskExt_lo_158 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_158 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_158 = {maskExt_hi_158, maskExt_lo_158};
  wire [15:0]        maskExt_lo_159 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_159 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_159 = {maskExt_hi_159, maskExt_lo_159};
  wire [15:0]        maskExt_lo_160 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_160 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_160 = {maskExt_hi_160, maskExt_lo_160};
  wire [15:0]        maskExt_lo_161 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_161 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_161 = {maskExt_hi_161, maskExt_lo_161};
  wire [15:0]        maskExt_lo_162 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_162 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_162 = {maskExt_hi_162, maskExt_lo_162};
  wire [15:0]        maskExt_lo_163 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_163 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_163 = {maskExt_hi_163, maskExt_lo_163};
  wire [15:0]        maskExt_lo_164 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_164 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_164 = {maskExt_hi_164, maskExt_lo_164};
  wire [15:0]        maskExt_lo_165 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_165 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_165 = {maskExt_hi_165, maskExt_lo_165};
  wire [15:0]        maskExt_lo_166 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_166 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_166 = {maskExt_hi_166, maskExt_lo_166};
  wire [15:0]        maskExt_lo_167 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_167 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_167 = {maskExt_hi_167, maskExt_lo_167};
  wire [15:0]        maskExt_lo_168 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_168 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_168 = {maskExt_hi_168, maskExt_lo_168};
  wire [15:0]        maskExt_lo_169 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_169 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_169 = {maskExt_hi_169, maskExt_lo_169};
  wire [15:0]        maskExt_lo_170 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_170 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_170 = {maskExt_hi_170, maskExt_lo_170};
  wire [15:0]        maskExt_lo_171 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_171 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_171 = {maskExt_hi_171, maskExt_lo_171};
  wire [15:0]        maskExt_lo_172 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_172 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_172 = {maskExt_hi_172, maskExt_lo_172};
  wire [15:0]        maskExt_lo_173 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_173 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_173 = {maskExt_hi_173, maskExt_lo_173};
  wire [15:0]        maskExt_lo_174 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_174 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_174 = {maskExt_hi_174, maskExt_lo_174};
  wire [15:0]        maskExt_lo_175 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_175 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_175 = {maskExt_hi_175, maskExt_lo_175};
  wire [15:0]        maskExt_lo_176 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_176 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_176 = {maskExt_hi_176, maskExt_lo_176};
  wire [15:0]        maskExt_lo_177 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_177 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_177 = {maskExt_hi_177, maskExt_lo_177};
  wire [15:0]        maskExt_lo_178 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_178 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_178 = {maskExt_hi_178, maskExt_lo_178};
  wire [15:0]        maskExt_lo_179 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_179 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_179 = {maskExt_hi_179, maskExt_lo_179};
  wire [15:0]        maskExt_lo_180 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_180 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_180 = {maskExt_hi_180, maskExt_lo_180};
  wire [15:0]        maskExt_lo_181 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_181 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_181 = {maskExt_hi_181, maskExt_lo_181};
  wire [15:0]        maskExt_lo_182 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_182 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_182 = {maskExt_hi_182, maskExt_lo_182};
  wire [15:0]        maskExt_lo_183 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_183 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_183 = {maskExt_hi_183, maskExt_lo_183};
  wire [15:0]        maskExt_lo_184 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_184 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_184 = {maskExt_hi_184, maskExt_lo_184};
  wire [15:0]        maskExt_lo_185 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_185 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_185 = {maskExt_hi_185, maskExt_lo_185};
  wire [15:0]        maskExt_lo_186 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_186 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_186 = {maskExt_hi_186, maskExt_lo_186};
  wire [15:0]        maskExt_lo_187 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_187 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_187 = {maskExt_hi_187, maskExt_lo_187};
  wire [15:0]        maskExt_lo_188 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_188 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_188 = {maskExt_hi_188, maskExt_lo_188};
  wire [15:0]        maskExt_lo_189 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_189 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_189 = {maskExt_hi_189, maskExt_lo_189};
  wire [15:0]        maskExt_lo_190 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_190 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_190 = {maskExt_hi_190, maskExt_lo_190};
  wire [15:0]        maskExt_lo_191 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_191 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_191 = {maskExt_hi_191, maskExt_lo_191};
  wire [15:0]        maskExt_lo_192 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_192 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_192 = {maskExt_hi_192, maskExt_lo_192};
  wire [15:0]        maskExt_lo_193 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_193 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_193 = {maskExt_hi_193, maskExt_lo_193};
  wire [15:0]        maskExt_lo_194 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_194 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_194 = {maskExt_hi_194, maskExt_lo_194};
  wire [15:0]        maskExt_lo_195 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_195 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_195 = {maskExt_hi_195, maskExt_lo_195};
  wire [15:0]        maskExt_lo_196 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_196 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_196 = {maskExt_hi_196, maskExt_lo_196};
  wire [15:0]        maskExt_lo_197 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_197 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_197 = {maskExt_hi_197, maskExt_lo_197};
  wire [15:0]        maskExt_lo_198 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_198 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_198 = {maskExt_hi_198, maskExt_lo_198};
  wire [15:0]        maskExt_lo_199 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_199 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_199 = {maskExt_hi_199, maskExt_lo_199};
  wire [15:0]        maskExt_lo_200 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_200 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_200 = {maskExt_hi_200, maskExt_lo_200};
  wire [15:0]        maskExt_lo_201 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_201 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_201 = {maskExt_hi_201, maskExt_lo_201};
  wire [15:0]        maskExt_lo_202 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_202 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_202 = {maskExt_hi_202, maskExt_lo_202};
  wire [15:0]        maskExt_lo_203 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_203 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_203 = {maskExt_hi_203, maskExt_lo_203};
  wire [15:0]        maskExt_lo_204 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_204 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_204 = {maskExt_hi_204, maskExt_lo_204};
  wire [15:0]        maskExt_lo_205 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_205 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_205 = {maskExt_hi_205, maskExt_lo_205};
  wire [15:0]        maskExt_lo_206 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_206 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_206 = {maskExt_hi_206, maskExt_lo_206};
  wire [15:0]        maskExt_lo_207 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_207 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_207 = {maskExt_hi_207, maskExt_lo_207};
  wire [15:0]        maskExt_lo_208 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_208 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_208 = {maskExt_hi_208, maskExt_lo_208};
  wire [15:0]        maskExt_lo_209 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_209 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_209 = {maskExt_hi_209, maskExt_lo_209};
  wire [15:0]        maskExt_lo_210 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_210 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_210 = {maskExt_hi_210, maskExt_lo_210};
  wire [15:0]        maskExt_lo_211 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_211 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_211 = {maskExt_hi_211, maskExt_lo_211};
  wire [15:0]        maskExt_lo_212 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_212 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_212 = {maskExt_hi_212, maskExt_lo_212};
  wire [15:0]        maskExt_lo_213 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_213 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_213 = {maskExt_hi_213, maskExt_lo_213};
  wire [15:0]        maskExt_lo_214 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_214 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_214 = {maskExt_hi_214, maskExt_lo_214};
  wire [15:0]        maskExt_lo_215 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_215 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_215 = {maskExt_hi_215, maskExt_lo_215};
  wire [15:0]        maskExt_lo_216 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_216 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_216 = {maskExt_hi_216, maskExt_lo_216};
  wire [15:0]        maskExt_lo_217 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_217 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_217 = {maskExt_hi_217, maskExt_lo_217};
  wire [15:0]        maskExt_lo_218 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_218 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_218 = {maskExt_hi_218, maskExt_lo_218};
  wire [15:0]        maskExt_lo_219 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_219 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_219 = {maskExt_hi_219, maskExt_lo_219};
  wire [15:0]        maskExt_lo_220 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_220 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_220 = {maskExt_hi_220, maskExt_lo_220};
  wire [15:0]        maskExt_lo_221 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_221 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_221 = {maskExt_hi_221, maskExt_lo_221};
  wire [15:0]        maskExt_lo_222 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_222 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_222 = {maskExt_hi_222, maskExt_lo_222};
  wire [15:0]        maskExt_lo_223 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_223 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_223 = {maskExt_hi_223, maskExt_lo_223};
  wire [15:0]        maskExt_lo_224 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_224 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_224 = {maskExt_hi_224, maskExt_lo_224};
  wire [15:0]        maskExt_lo_225 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_225 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_225 = {maskExt_hi_225, maskExt_lo_225};
  wire [15:0]        maskExt_lo_226 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_226 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_226 = {maskExt_hi_226, maskExt_lo_226};
  wire [15:0]        maskExt_lo_227 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_227 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_227 = {maskExt_hi_227, maskExt_lo_227};
  wire [15:0]        maskExt_lo_228 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_228 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_228 = {maskExt_hi_228, maskExt_lo_228};
  wire [15:0]        maskExt_lo_229 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_229 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_229 = {maskExt_hi_229, maskExt_lo_229};
  wire [15:0]        maskExt_lo_230 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_230 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_230 = {maskExt_hi_230, maskExt_lo_230};
  wire [15:0]        maskExt_lo_231 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_231 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_231 = {maskExt_hi_231, maskExt_lo_231};
  wire [15:0]        maskExt_lo_232 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_232 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_232 = {maskExt_hi_232, maskExt_lo_232};
  wire [15:0]        maskExt_lo_233 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_233 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_233 = {maskExt_hi_233, maskExt_lo_233};
  wire [15:0]        maskExt_lo_234 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_234 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_234 = {maskExt_hi_234, maskExt_lo_234};
  wire [15:0]        maskExt_lo_235 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_235 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_235 = {maskExt_hi_235, maskExt_lo_235};
  wire [15:0]        maskExt_lo_236 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_236 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_236 = {maskExt_hi_236, maskExt_lo_236};
  wire [15:0]        maskExt_lo_237 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_237 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_237 = {maskExt_hi_237, maskExt_lo_237};
  wire [15:0]        maskExt_lo_238 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_238 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_238 = {maskExt_hi_238, maskExt_lo_238};
  wire [15:0]        maskExt_lo_239 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_239 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_239 = {maskExt_hi_239, maskExt_lo_239};
  wire [15:0]        maskExt_lo_240 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_240 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_240 = {maskExt_hi_240, maskExt_lo_240};
  wire [15:0]        maskExt_lo_241 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_241 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_241 = {maskExt_hi_241, maskExt_lo_241};
  wire [15:0]        maskExt_lo_242 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_242 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_242 = {maskExt_hi_242, maskExt_lo_242};
  wire [15:0]        maskExt_lo_243 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_243 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_243 = {maskExt_hi_243, maskExt_lo_243};
  wire [15:0]        maskExt_lo_244 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_244 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_244 = {maskExt_hi_244, maskExt_lo_244};
  wire [15:0]        maskExt_lo_245 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_245 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_245 = {maskExt_hi_245, maskExt_lo_245};
  wire [15:0]        maskExt_lo_246 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_246 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_246 = {maskExt_hi_246, maskExt_lo_246};
  wire [15:0]        maskExt_lo_247 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_247 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_247 = {maskExt_hi_247, maskExt_lo_247};
  wire [15:0]        maskExt_lo_248 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_248 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_248 = {maskExt_hi_248, maskExt_lo_248};
  wire [15:0]        maskExt_lo_249 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_249 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_249 = {maskExt_hi_249, maskExt_lo_249};
  wire [15:0]        maskExt_lo_250 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_250 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_250 = {maskExt_hi_250, maskExt_lo_250};
  wire [15:0]        maskExt_lo_251 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_251 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_251 = {maskExt_hi_251, maskExt_lo_251};
  wire [15:0]        maskExt_lo_252 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_252 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_252 = {maskExt_hi_252, maskExt_lo_252};
  wire [15:0]        maskExt_lo_253 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_253 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_253 = {maskExt_hi_253, maskExt_lo_253};
  wire [15:0]        maskExt_lo_254 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_254 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_254 = {maskExt_hi_254, maskExt_lo_254};
  wire [15:0]        maskExt_lo_255 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_255 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_255 = {maskExt_hi_255, maskExt_lo_255};
  wire               alwaysMerge = {request_bits_instructionInformation_mop_0, request_bits_instructionInformation_lumop_0[2:0], request_bits_instructionInformation_lumop_0[4]} == 6'h0;
  wire               useLoadUnit = alwaysMerge & ~request_bits_instructionInformation_isStore_0;
  wire               useStoreUnit = alwaysMerge & request_bits_instructionInformation_isStore_0;
  wire               useOtherUnit = ~alwaysMerge;
  wire               addressCheck = _otherUnit_status_idle & (~useOtherUnit | _loadUnit_status_idle & _storeUnit_status_idle);
  wire               unitReady = useLoadUnit & _loadUnit_status_idle | useStoreUnit & _storeUnit_status_idle | useOtherUnit & _otherUnit_status_idle;
  wire               request_ready_0 = unitReady & addressCheck;
  wire               requestFire = request_ready_0 & request_valid_0;
  wire               reqEnq_0 = useLoadUnit & requestFire;
  wire               reqEnq_1 = useStoreUnit & requestFire;
  wire               reqEnq_2 = useOtherUnit & requestFire;
  wire [8:0]         maskSelect = _loadUnit_maskSelect_valid ? _loadUnit_maskSelect_bits : 9'h0;
  wire [63:0]        _GEN = {v0_1, v0_0};
  wire [63:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo = _GEN;
  wire [63:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo = _GEN;
  wire [63:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo = _GEN;
  wire [63:0]        _GEN_0 = {v0_3, v0_2};
  wire [63:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi = _GEN_0;
  wire [63:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi = _GEN_0;
  wire [63:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi = _GEN_0;
  wire [127:0]       loadUnit_maskInput_lo_lo_lo_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo};
  wire [63:0]        _GEN_1 = {v0_5, v0_4};
  wire [63:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo = _GEN_1;
  wire [63:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo = _GEN_1;
  wire [63:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo = _GEN_1;
  wire [63:0]        _GEN_2 = {v0_7, v0_6};
  wire [63:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi = _GEN_2;
  wire [63:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi = _GEN_2;
  wire [63:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi = _GEN_2;
  wire [127:0]       loadUnit_maskInput_lo_lo_lo_lo_lo_hi = {loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]       loadUnit_maskInput_lo_lo_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_lo};
  wire [63:0]        _GEN_3 = {v0_9, v0_8};
  wire [63:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo = _GEN_3;
  wire [63:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo = _GEN_3;
  wire [63:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo = _GEN_3;
  wire [63:0]        _GEN_4 = {v0_11, v0_10};
  wire [63:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi = _GEN_4;
  wire [63:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi = _GEN_4;
  wire [63:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi = _GEN_4;
  wire [127:0]       loadUnit_maskInput_lo_lo_lo_lo_hi_lo = {loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo};
  wire [63:0]        _GEN_5 = {v0_13, v0_12};
  wire [63:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo = _GEN_5;
  wire [63:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo = _GEN_5;
  wire [63:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo = _GEN_5;
  wire [63:0]        _GEN_6 = {v0_15, v0_14};
  wire [63:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi = _GEN_6;
  wire [63:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi = _GEN_6;
  wire [63:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi = _GEN_6;
  wire [127:0]       loadUnit_maskInput_lo_lo_lo_lo_hi_hi = {loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]       loadUnit_maskInput_lo_lo_lo_lo_hi = {loadUnit_maskInput_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_lo};
  wire [511:0]       loadUnit_maskInput_lo_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_lo};
  wire [63:0]        _GEN_7 = {v0_17, v0_16};
  wire [63:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo = _GEN_7;
  wire [63:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo = _GEN_7;
  wire [63:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo = _GEN_7;
  wire [63:0]        _GEN_8 = {v0_19, v0_18};
  wire [63:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi = _GEN_8;
  wire [63:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi = _GEN_8;
  wire [63:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi = _GEN_8;
  wire [127:0]       loadUnit_maskInput_lo_lo_lo_hi_lo_lo = {loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo};
  wire [63:0]        _GEN_9 = {v0_21, v0_20};
  wire [63:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo = _GEN_9;
  wire [63:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo = _GEN_9;
  wire [63:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo = _GEN_9;
  wire [63:0]        _GEN_10 = {v0_23, v0_22};
  wire [63:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi = _GEN_10;
  wire [63:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi = _GEN_10;
  wire [63:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi = _GEN_10;
  wire [127:0]       loadUnit_maskInput_lo_lo_lo_hi_lo_hi = {loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]       loadUnit_maskInput_lo_lo_lo_hi_lo = {loadUnit_maskInput_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_lo};
  wire [63:0]        _GEN_11 = {v0_25, v0_24};
  wire [63:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo = _GEN_11;
  wire [63:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo = _GEN_11;
  wire [63:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo = _GEN_11;
  wire [63:0]        _GEN_12 = {v0_27, v0_26};
  wire [63:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi = _GEN_12;
  wire [63:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi = _GEN_12;
  wire [63:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi = _GEN_12;
  wire [127:0]       loadUnit_maskInput_lo_lo_lo_hi_hi_lo = {loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo};
  wire [63:0]        _GEN_13 = {v0_29, v0_28};
  wire [63:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo = _GEN_13;
  wire [63:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo = _GEN_13;
  wire [63:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo = _GEN_13;
  wire [63:0]        _GEN_14 = {v0_31, v0_30};
  wire [63:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi = _GEN_14;
  wire [63:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi = _GEN_14;
  wire [63:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi = _GEN_14;
  wire [127:0]       loadUnit_maskInput_lo_lo_lo_hi_hi_hi = {loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]       loadUnit_maskInput_lo_lo_lo_hi_hi = {loadUnit_maskInput_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_lo};
  wire [511:0]       loadUnit_maskInput_lo_lo_lo_hi = {loadUnit_maskInput_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_lo};
  wire [1023:0]      loadUnit_maskInput_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo};
  wire [63:0]        _GEN_15 = {v0_33, v0_32};
  wire [63:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo = _GEN_15;
  wire [63:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo = _GEN_15;
  wire [63:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo = _GEN_15;
  wire [63:0]        _GEN_16 = {v0_35, v0_34};
  wire [63:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi = _GEN_16;
  wire [63:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi = _GEN_16;
  wire [63:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi = _GEN_16;
  wire [127:0]       loadUnit_maskInput_lo_lo_hi_lo_lo_lo = {loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo};
  wire [63:0]        _GEN_17 = {v0_37, v0_36};
  wire [63:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo = _GEN_17;
  wire [63:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo = _GEN_17;
  wire [63:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo = _GEN_17;
  wire [63:0]        _GEN_18 = {v0_39, v0_38};
  wire [63:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi = _GEN_18;
  wire [63:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi = _GEN_18;
  wire [63:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi = _GEN_18;
  wire [127:0]       loadUnit_maskInput_lo_lo_hi_lo_lo_hi = {loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]       loadUnit_maskInput_lo_lo_hi_lo_lo = {loadUnit_maskInput_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_lo};
  wire [63:0]        _GEN_19 = {v0_41, v0_40};
  wire [63:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo = _GEN_19;
  wire [63:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo = _GEN_19;
  wire [63:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo = _GEN_19;
  wire [63:0]        _GEN_20 = {v0_43, v0_42};
  wire [63:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi = _GEN_20;
  wire [63:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi = _GEN_20;
  wire [63:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi = _GEN_20;
  wire [127:0]       loadUnit_maskInput_lo_lo_hi_lo_hi_lo = {loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo};
  wire [63:0]        _GEN_21 = {v0_45, v0_44};
  wire [63:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo = _GEN_21;
  wire [63:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo = _GEN_21;
  wire [63:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo = _GEN_21;
  wire [63:0]        _GEN_22 = {v0_47, v0_46};
  wire [63:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi = _GEN_22;
  wire [63:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi = _GEN_22;
  wire [63:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi = _GEN_22;
  wire [127:0]       loadUnit_maskInput_lo_lo_hi_lo_hi_hi = {loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]       loadUnit_maskInput_lo_lo_hi_lo_hi = {loadUnit_maskInput_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_lo};
  wire [511:0]       loadUnit_maskInput_lo_lo_hi_lo = {loadUnit_maskInput_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_lo};
  wire [63:0]        _GEN_23 = {v0_49, v0_48};
  wire [63:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo = _GEN_23;
  wire [63:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo = _GEN_23;
  wire [63:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo = _GEN_23;
  wire [63:0]        _GEN_24 = {v0_51, v0_50};
  wire [63:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi = _GEN_24;
  wire [63:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi = _GEN_24;
  wire [63:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi = _GEN_24;
  wire [127:0]       loadUnit_maskInput_lo_lo_hi_hi_lo_lo = {loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo};
  wire [63:0]        _GEN_25 = {v0_53, v0_52};
  wire [63:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo = _GEN_25;
  wire [63:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo = _GEN_25;
  wire [63:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo = _GEN_25;
  wire [63:0]        _GEN_26 = {v0_55, v0_54};
  wire [63:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi = _GEN_26;
  wire [63:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi = _GEN_26;
  wire [63:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi = _GEN_26;
  wire [127:0]       loadUnit_maskInput_lo_lo_hi_hi_lo_hi = {loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]       loadUnit_maskInput_lo_lo_hi_hi_lo = {loadUnit_maskInput_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_lo};
  wire [63:0]        _GEN_27 = {v0_57, v0_56};
  wire [63:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo = _GEN_27;
  wire [63:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo = _GEN_27;
  wire [63:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo = _GEN_27;
  wire [63:0]        _GEN_28 = {v0_59, v0_58};
  wire [63:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi = _GEN_28;
  wire [63:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi = _GEN_28;
  wire [63:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi = _GEN_28;
  wire [127:0]       loadUnit_maskInput_lo_lo_hi_hi_hi_lo = {loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo};
  wire [63:0]        _GEN_29 = {v0_61, v0_60};
  wire [63:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo = _GEN_29;
  wire [63:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo = _GEN_29;
  wire [63:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo = _GEN_29;
  wire [63:0]        _GEN_30 = {v0_63, v0_62};
  wire [63:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi = _GEN_30;
  wire [63:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi = _GEN_30;
  wire [63:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi = _GEN_30;
  wire [127:0]       loadUnit_maskInput_lo_lo_hi_hi_hi_hi = {loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]       loadUnit_maskInput_lo_lo_hi_hi_hi = {loadUnit_maskInput_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_lo};
  wire [511:0]       loadUnit_maskInput_lo_lo_hi_hi = {loadUnit_maskInput_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_lo};
  wire [1023:0]      loadUnit_maskInput_lo_lo_hi = {loadUnit_maskInput_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo};
  wire [2047:0]      loadUnit_maskInput_lo_lo = {loadUnit_maskInput_lo_lo_hi, loadUnit_maskInput_lo_lo_lo};
  wire [63:0]        _GEN_31 = {v0_65, v0_64};
  wire [63:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo = _GEN_31;
  wire [63:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo = _GEN_31;
  wire [63:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo = _GEN_31;
  wire [63:0]        _GEN_32 = {v0_67, v0_66};
  wire [63:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi = _GEN_32;
  wire [63:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi = _GEN_32;
  wire [63:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi = _GEN_32;
  wire [127:0]       loadUnit_maskInput_lo_hi_lo_lo_lo_lo = {loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo};
  wire [63:0]        _GEN_33 = {v0_69, v0_68};
  wire [63:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo = _GEN_33;
  wire [63:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo = _GEN_33;
  wire [63:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo = _GEN_33;
  wire [63:0]        _GEN_34 = {v0_71, v0_70};
  wire [63:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi = _GEN_34;
  wire [63:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi = _GEN_34;
  wire [63:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi = _GEN_34;
  wire [127:0]       loadUnit_maskInput_lo_hi_lo_lo_lo_hi = {loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]       loadUnit_maskInput_lo_hi_lo_lo_lo = {loadUnit_maskInput_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_lo};
  wire [63:0]        _GEN_35 = {v0_73, v0_72};
  wire [63:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo = _GEN_35;
  wire [63:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo = _GEN_35;
  wire [63:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo = _GEN_35;
  wire [63:0]        _GEN_36 = {v0_75, v0_74};
  wire [63:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi = _GEN_36;
  wire [63:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi = _GEN_36;
  wire [63:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi = _GEN_36;
  wire [127:0]       loadUnit_maskInput_lo_hi_lo_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo};
  wire [63:0]        _GEN_37 = {v0_77, v0_76};
  wire [63:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo = _GEN_37;
  wire [63:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo = _GEN_37;
  wire [63:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo = _GEN_37;
  wire [63:0]        _GEN_38 = {v0_79, v0_78};
  wire [63:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi = _GEN_38;
  wire [63:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi = _GEN_38;
  wire [63:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi = _GEN_38;
  wire [127:0]       loadUnit_maskInput_lo_hi_lo_lo_hi_hi = {loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]       loadUnit_maskInput_lo_hi_lo_lo_hi = {loadUnit_maskInput_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_lo};
  wire [511:0]       loadUnit_maskInput_lo_hi_lo_lo = {loadUnit_maskInput_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_lo};
  wire [63:0]        _GEN_39 = {v0_81, v0_80};
  wire [63:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo = _GEN_39;
  wire [63:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo = _GEN_39;
  wire [63:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo = _GEN_39;
  wire [63:0]        _GEN_40 = {v0_83, v0_82};
  wire [63:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi = _GEN_40;
  wire [63:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi = _GEN_40;
  wire [63:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi = _GEN_40;
  wire [127:0]       loadUnit_maskInput_lo_hi_lo_hi_lo_lo = {loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo};
  wire [63:0]        _GEN_41 = {v0_85, v0_84};
  wire [63:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo = _GEN_41;
  wire [63:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo = _GEN_41;
  wire [63:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo = _GEN_41;
  wire [63:0]        _GEN_42 = {v0_87, v0_86};
  wire [63:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi = _GEN_42;
  wire [63:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi = _GEN_42;
  wire [63:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi = _GEN_42;
  wire [127:0]       loadUnit_maskInput_lo_hi_lo_hi_lo_hi = {loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]       loadUnit_maskInput_lo_hi_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_lo};
  wire [63:0]        _GEN_43 = {v0_89, v0_88};
  wire [63:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo = _GEN_43;
  wire [63:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo = _GEN_43;
  wire [63:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo = _GEN_43;
  wire [63:0]        _GEN_44 = {v0_91, v0_90};
  wire [63:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi = _GEN_44;
  wire [63:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi = _GEN_44;
  wire [63:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi = _GEN_44;
  wire [127:0]       loadUnit_maskInput_lo_hi_lo_hi_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo};
  wire [63:0]        _GEN_45 = {v0_93, v0_92};
  wire [63:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo = _GEN_45;
  wire [63:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo = _GEN_45;
  wire [63:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo = _GEN_45;
  wire [63:0]        _GEN_46 = {v0_95, v0_94};
  wire [63:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi = _GEN_46;
  wire [63:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi = _GEN_46;
  wire [63:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi = _GEN_46;
  wire [127:0]       loadUnit_maskInput_lo_hi_lo_hi_hi_hi = {loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]       loadUnit_maskInput_lo_hi_lo_hi_hi = {loadUnit_maskInput_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_lo};
  wire [511:0]       loadUnit_maskInput_lo_hi_lo_hi = {loadUnit_maskInput_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_lo};
  wire [1023:0]      loadUnit_maskInput_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_lo};
  wire [63:0]        _GEN_47 = {v0_97, v0_96};
  wire [63:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo = _GEN_47;
  wire [63:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo = _GEN_47;
  wire [63:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo = _GEN_47;
  wire [63:0]        _GEN_48 = {v0_99, v0_98};
  wire [63:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi = _GEN_48;
  wire [63:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi = _GEN_48;
  wire [63:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi = _GEN_48;
  wire [127:0]       loadUnit_maskInput_lo_hi_hi_lo_lo_lo = {loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo};
  wire [63:0]        _GEN_49 = {v0_101, v0_100};
  wire [63:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo = _GEN_49;
  wire [63:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo = _GEN_49;
  wire [63:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo = _GEN_49;
  wire [63:0]        _GEN_50 = {v0_103, v0_102};
  wire [63:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi = _GEN_50;
  wire [63:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi = _GEN_50;
  wire [63:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi = _GEN_50;
  wire [127:0]       loadUnit_maskInput_lo_hi_hi_lo_lo_hi = {loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]       loadUnit_maskInput_lo_hi_hi_lo_lo = {loadUnit_maskInput_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_lo};
  wire [63:0]        _GEN_51 = {v0_105, v0_104};
  wire [63:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo = _GEN_51;
  wire [63:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo = _GEN_51;
  wire [63:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo = _GEN_51;
  wire [63:0]        _GEN_52 = {v0_107, v0_106};
  wire [63:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi = _GEN_52;
  wire [63:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi = _GEN_52;
  wire [63:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi = _GEN_52;
  wire [127:0]       loadUnit_maskInput_lo_hi_hi_lo_hi_lo = {loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo};
  wire [63:0]        _GEN_53 = {v0_109, v0_108};
  wire [63:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo = _GEN_53;
  wire [63:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo = _GEN_53;
  wire [63:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo = _GEN_53;
  wire [63:0]        _GEN_54 = {v0_111, v0_110};
  wire [63:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi = _GEN_54;
  wire [63:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi = _GEN_54;
  wire [63:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi = _GEN_54;
  wire [127:0]       loadUnit_maskInput_lo_hi_hi_lo_hi_hi = {loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]       loadUnit_maskInput_lo_hi_hi_lo_hi = {loadUnit_maskInput_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_lo};
  wire [511:0]       loadUnit_maskInput_lo_hi_hi_lo = {loadUnit_maskInput_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_lo};
  wire [63:0]        _GEN_55 = {v0_113, v0_112};
  wire [63:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo = _GEN_55;
  wire [63:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo = _GEN_55;
  wire [63:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo = _GEN_55;
  wire [63:0]        _GEN_56 = {v0_115, v0_114};
  wire [63:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi = _GEN_56;
  wire [63:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi = _GEN_56;
  wire [63:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi = _GEN_56;
  wire [127:0]       loadUnit_maskInput_lo_hi_hi_hi_lo_lo = {loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo};
  wire [63:0]        _GEN_57 = {v0_117, v0_116};
  wire [63:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo = _GEN_57;
  wire [63:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo = _GEN_57;
  wire [63:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo = _GEN_57;
  wire [63:0]        _GEN_58 = {v0_119, v0_118};
  wire [63:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi = _GEN_58;
  wire [63:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi = _GEN_58;
  wire [63:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi = _GEN_58;
  wire [127:0]       loadUnit_maskInput_lo_hi_hi_hi_lo_hi = {loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]       loadUnit_maskInput_lo_hi_hi_hi_lo = {loadUnit_maskInput_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_lo};
  wire [63:0]        _GEN_59 = {v0_121, v0_120};
  wire [63:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo = _GEN_59;
  wire [63:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo = _GEN_59;
  wire [63:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo = _GEN_59;
  wire [63:0]        _GEN_60 = {v0_123, v0_122};
  wire [63:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi = _GEN_60;
  wire [63:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi = _GEN_60;
  wire [63:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi = _GEN_60;
  wire [127:0]       loadUnit_maskInput_lo_hi_hi_hi_hi_lo = {loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo};
  wire [63:0]        _GEN_61 = {v0_125, v0_124};
  wire [63:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo = _GEN_61;
  wire [63:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo = _GEN_61;
  wire [63:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo = _GEN_61;
  wire [63:0]        _GEN_62 = {v0_127, v0_126};
  wire [63:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi = _GEN_62;
  wire [63:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi = _GEN_62;
  wire [63:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi = _GEN_62;
  wire [127:0]       loadUnit_maskInput_lo_hi_hi_hi_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]       loadUnit_maskInput_lo_hi_hi_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_lo};
  wire [511:0]       loadUnit_maskInput_lo_hi_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_lo};
  wire [1023:0]      loadUnit_maskInput_lo_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_lo};
  wire [2047:0]      loadUnit_maskInput_lo_hi = {loadUnit_maskInput_lo_hi_hi, loadUnit_maskInput_lo_hi_lo};
  wire [4095:0]      loadUnit_maskInput_lo = {loadUnit_maskInput_lo_hi, loadUnit_maskInput_lo_lo};
  wire [63:0]        _GEN_63 = {v0_129, v0_128};
  wire [63:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo = _GEN_63;
  wire [63:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo = _GEN_63;
  wire [63:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo = _GEN_63;
  wire [63:0]        _GEN_64 = {v0_131, v0_130};
  wire [63:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi = _GEN_64;
  wire [63:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi = _GEN_64;
  wire [63:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi = _GEN_64;
  wire [127:0]       loadUnit_maskInput_hi_lo_lo_lo_lo_lo = {loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo};
  wire [63:0]        _GEN_65 = {v0_133, v0_132};
  wire [63:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo = _GEN_65;
  wire [63:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo = _GEN_65;
  wire [63:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo = _GEN_65;
  wire [63:0]        _GEN_66 = {v0_135, v0_134};
  wire [63:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi = _GEN_66;
  wire [63:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi = _GEN_66;
  wire [63:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi = _GEN_66;
  wire [127:0]       loadUnit_maskInput_hi_lo_lo_lo_lo_hi = {loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]       loadUnit_maskInput_hi_lo_lo_lo_lo = {loadUnit_maskInput_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_lo};
  wire [63:0]        _GEN_67 = {v0_137, v0_136};
  wire [63:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo = _GEN_67;
  wire [63:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo = _GEN_67;
  wire [63:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo = _GEN_67;
  wire [63:0]        _GEN_68 = {v0_139, v0_138};
  wire [63:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi = _GEN_68;
  wire [63:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi = _GEN_68;
  wire [63:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi = _GEN_68;
  wire [127:0]       loadUnit_maskInput_hi_lo_lo_lo_hi_lo = {loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo};
  wire [63:0]        _GEN_69 = {v0_141, v0_140};
  wire [63:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo = _GEN_69;
  wire [63:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo = _GEN_69;
  wire [63:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo = _GEN_69;
  wire [63:0]        _GEN_70 = {v0_143, v0_142};
  wire [63:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi = _GEN_70;
  wire [63:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi = _GEN_70;
  wire [63:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi = _GEN_70;
  wire [127:0]       loadUnit_maskInput_hi_lo_lo_lo_hi_hi = {loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]       loadUnit_maskInput_hi_lo_lo_lo_hi = {loadUnit_maskInput_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_lo};
  wire [511:0]       loadUnit_maskInput_hi_lo_lo_lo = {loadUnit_maskInput_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_lo};
  wire [63:0]        _GEN_71 = {v0_145, v0_144};
  wire [63:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo = _GEN_71;
  wire [63:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo = _GEN_71;
  wire [63:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo = _GEN_71;
  wire [63:0]        _GEN_72 = {v0_147, v0_146};
  wire [63:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi = _GEN_72;
  wire [63:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi = _GEN_72;
  wire [63:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi = _GEN_72;
  wire [127:0]       loadUnit_maskInput_hi_lo_lo_hi_lo_lo = {loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo};
  wire [63:0]        _GEN_73 = {v0_149, v0_148};
  wire [63:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo = _GEN_73;
  wire [63:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo = _GEN_73;
  wire [63:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo = _GEN_73;
  wire [63:0]        _GEN_74 = {v0_151, v0_150};
  wire [63:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi = _GEN_74;
  wire [63:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi = _GEN_74;
  wire [63:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi = _GEN_74;
  wire [127:0]       loadUnit_maskInput_hi_lo_lo_hi_lo_hi = {loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]       loadUnit_maskInput_hi_lo_lo_hi_lo = {loadUnit_maskInput_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_lo};
  wire [63:0]        _GEN_75 = {v0_153, v0_152};
  wire [63:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo = _GEN_75;
  wire [63:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo = _GEN_75;
  wire [63:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo = _GEN_75;
  wire [63:0]        _GEN_76 = {v0_155, v0_154};
  wire [63:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi = _GEN_76;
  wire [63:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi = _GEN_76;
  wire [63:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi = _GEN_76;
  wire [127:0]       loadUnit_maskInput_hi_lo_lo_hi_hi_lo = {loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo};
  wire [63:0]        _GEN_77 = {v0_157, v0_156};
  wire [63:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo = _GEN_77;
  wire [63:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo = _GEN_77;
  wire [63:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo = _GEN_77;
  wire [63:0]        _GEN_78 = {v0_159, v0_158};
  wire [63:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi = _GEN_78;
  wire [63:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi = _GEN_78;
  wire [63:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi = _GEN_78;
  wire [127:0]       loadUnit_maskInput_hi_lo_lo_hi_hi_hi = {loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]       loadUnit_maskInput_hi_lo_lo_hi_hi = {loadUnit_maskInput_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_lo};
  wire [511:0]       loadUnit_maskInput_hi_lo_lo_hi = {loadUnit_maskInput_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_lo};
  wire [1023:0]      loadUnit_maskInput_hi_lo_lo = {loadUnit_maskInput_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo};
  wire [63:0]        _GEN_79 = {v0_161, v0_160};
  wire [63:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo = _GEN_79;
  wire [63:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo = _GEN_79;
  wire [63:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo = _GEN_79;
  wire [63:0]        _GEN_80 = {v0_163, v0_162};
  wire [63:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi = _GEN_80;
  wire [63:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi = _GEN_80;
  wire [63:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi = _GEN_80;
  wire [127:0]       loadUnit_maskInput_hi_lo_hi_lo_lo_lo = {loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo};
  wire [63:0]        _GEN_81 = {v0_165, v0_164};
  wire [63:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo = _GEN_81;
  wire [63:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo = _GEN_81;
  wire [63:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo = _GEN_81;
  wire [63:0]        _GEN_82 = {v0_167, v0_166};
  wire [63:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi = _GEN_82;
  wire [63:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi = _GEN_82;
  wire [63:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi = _GEN_82;
  wire [127:0]       loadUnit_maskInput_hi_lo_hi_lo_lo_hi = {loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]       loadUnit_maskInput_hi_lo_hi_lo_lo = {loadUnit_maskInput_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_lo};
  wire [63:0]        _GEN_83 = {v0_169, v0_168};
  wire [63:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo = _GEN_83;
  wire [63:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo = _GEN_83;
  wire [63:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo = _GEN_83;
  wire [63:0]        _GEN_84 = {v0_171, v0_170};
  wire [63:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi = _GEN_84;
  wire [63:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi = _GEN_84;
  wire [63:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi = _GEN_84;
  wire [127:0]       loadUnit_maskInput_hi_lo_hi_lo_hi_lo = {loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo};
  wire [63:0]        _GEN_85 = {v0_173, v0_172};
  wire [63:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo = _GEN_85;
  wire [63:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo = _GEN_85;
  wire [63:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo = _GEN_85;
  wire [63:0]        _GEN_86 = {v0_175, v0_174};
  wire [63:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi = _GEN_86;
  wire [63:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi = _GEN_86;
  wire [63:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi = _GEN_86;
  wire [127:0]       loadUnit_maskInput_hi_lo_hi_lo_hi_hi = {loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]       loadUnit_maskInput_hi_lo_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_lo};
  wire [511:0]       loadUnit_maskInput_hi_lo_hi_lo = {loadUnit_maskInput_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_lo};
  wire [63:0]        _GEN_87 = {v0_177, v0_176};
  wire [63:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo = _GEN_87;
  wire [63:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo = _GEN_87;
  wire [63:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo = _GEN_87;
  wire [63:0]        _GEN_88 = {v0_179, v0_178};
  wire [63:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi = _GEN_88;
  wire [63:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi = _GEN_88;
  wire [63:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi = _GEN_88;
  wire [127:0]       loadUnit_maskInput_hi_lo_hi_hi_lo_lo = {loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo};
  wire [63:0]        _GEN_89 = {v0_181, v0_180};
  wire [63:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo = _GEN_89;
  wire [63:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo = _GEN_89;
  wire [63:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo = _GEN_89;
  wire [63:0]        _GEN_90 = {v0_183, v0_182};
  wire [63:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi = _GEN_90;
  wire [63:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi = _GEN_90;
  wire [63:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi = _GEN_90;
  wire [127:0]       loadUnit_maskInput_hi_lo_hi_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]       loadUnit_maskInput_hi_lo_hi_hi_lo = {loadUnit_maskInput_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_lo};
  wire [63:0]        _GEN_91 = {v0_185, v0_184};
  wire [63:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo = _GEN_91;
  wire [63:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo = _GEN_91;
  wire [63:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo = _GEN_91;
  wire [63:0]        _GEN_92 = {v0_187, v0_186};
  wire [63:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi = _GEN_92;
  wire [63:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi = _GEN_92;
  wire [63:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi = _GEN_92;
  wire [127:0]       loadUnit_maskInput_hi_lo_hi_hi_hi_lo = {loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo};
  wire [63:0]        _GEN_93 = {v0_189, v0_188};
  wire [63:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo = _GEN_93;
  wire [63:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo = _GEN_93;
  wire [63:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo = _GEN_93;
  wire [63:0]        _GEN_94 = {v0_191, v0_190};
  wire [63:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi = _GEN_94;
  wire [63:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi = _GEN_94;
  wire [63:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi = _GEN_94;
  wire [127:0]       loadUnit_maskInput_hi_lo_hi_hi_hi_hi = {loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]       loadUnit_maskInput_hi_lo_hi_hi_hi = {loadUnit_maskInput_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_lo};
  wire [511:0]       loadUnit_maskInput_hi_lo_hi_hi = {loadUnit_maskInput_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_lo};
  wire [1023:0]      loadUnit_maskInput_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo};
  wire [2047:0]      loadUnit_maskInput_hi_lo = {loadUnit_maskInput_hi_lo_hi, loadUnit_maskInput_hi_lo_lo};
  wire [63:0]        _GEN_95 = {v0_193, v0_192};
  wire [63:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo = _GEN_95;
  wire [63:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo = _GEN_95;
  wire [63:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo = _GEN_95;
  wire [63:0]        _GEN_96 = {v0_195, v0_194};
  wire [63:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi = _GEN_96;
  wire [63:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi = _GEN_96;
  wire [63:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi = _GEN_96;
  wire [127:0]       loadUnit_maskInput_hi_hi_lo_lo_lo_lo = {loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo};
  wire [63:0]        _GEN_97 = {v0_197, v0_196};
  wire [63:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo = _GEN_97;
  wire [63:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo = _GEN_97;
  wire [63:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo = _GEN_97;
  wire [63:0]        _GEN_98 = {v0_199, v0_198};
  wire [63:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi = _GEN_98;
  wire [63:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi = _GEN_98;
  wire [63:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi = _GEN_98;
  wire [127:0]       loadUnit_maskInput_hi_hi_lo_lo_lo_hi = {loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]       loadUnit_maskInput_hi_hi_lo_lo_lo = {loadUnit_maskInput_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_lo};
  wire [63:0]        _GEN_99 = {v0_201, v0_200};
  wire [63:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo = _GEN_99;
  wire [63:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo = _GEN_99;
  wire [63:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo = _GEN_99;
  wire [63:0]        _GEN_100 = {v0_203, v0_202};
  wire [63:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi = _GEN_100;
  wire [63:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi = _GEN_100;
  wire [63:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi = _GEN_100;
  wire [127:0]       loadUnit_maskInput_hi_hi_lo_lo_hi_lo = {loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo};
  wire [63:0]        _GEN_101 = {v0_205, v0_204};
  wire [63:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo = _GEN_101;
  wire [63:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo = _GEN_101;
  wire [63:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo = _GEN_101;
  wire [63:0]        _GEN_102 = {v0_207, v0_206};
  wire [63:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi = _GEN_102;
  wire [63:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi = _GEN_102;
  wire [63:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi = _GEN_102;
  wire [127:0]       loadUnit_maskInput_hi_hi_lo_lo_hi_hi = {loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]       loadUnit_maskInput_hi_hi_lo_lo_hi = {loadUnit_maskInput_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_lo};
  wire [511:0]       loadUnit_maskInput_hi_hi_lo_lo = {loadUnit_maskInput_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_lo};
  wire [63:0]        _GEN_103 = {v0_209, v0_208};
  wire [63:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo = _GEN_103;
  wire [63:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo = _GEN_103;
  wire [63:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo = _GEN_103;
  wire [63:0]        _GEN_104 = {v0_211, v0_210};
  wire [63:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi = _GEN_104;
  wire [63:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi = _GEN_104;
  wire [63:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi = _GEN_104;
  wire [127:0]       loadUnit_maskInput_hi_hi_lo_hi_lo_lo = {loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo};
  wire [63:0]        _GEN_105 = {v0_213, v0_212};
  wire [63:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo = _GEN_105;
  wire [63:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo = _GEN_105;
  wire [63:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo = _GEN_105;
  wire [63:0]        _GEN_106 = {v0_215, v0_214};
  wire [63:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi = _GEN_106;
  wire [63:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi = _GEN_106;
  wire [63:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi = _GEN_106;
  wire [127:0]       loadUnit_maskInput_hi_hi_lo_hi_lo_hi = {loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]       loadUnit_maskInput_hi_hi_lo_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_lo};
  wire [63:0]        _GEN_107 = {v0_217, v0_216};
  wire [63:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo = _GEN_107;
  wire [63:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo = _GEN_107;
  wire [63:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo = _GEN_107;
  wire [63:0]        _GEN_108 = {v0_219, v0_218};
  wire [63:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi = _GEN_108;
  wire [63:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi = _GEN_108;
  wire [63:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi = _GEN_108;
  wire [127:0]       loadUnit_maskInput_hi_hi_lo_hi_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo};
  wire [63:0]        _GEN_109 = {v0_221, v0_220};
  wire [63:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo = _GEN_109;
  wire [63:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo = _GEN_109;
  wire [63:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo = _GEN_109;
  wire [63:0]        _GEN_110 = {v0_223, v0_222};
  wire [63:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi = _GEN_110;
  wire [63:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi = _GEN_110;
  wire [63:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi = _GEN_110;
  wire [127:0]       loadUnit_maskInput_hi_hi_lo_hi_hi_hi = {loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]       loadUnit_maskInput_hi_hi_lo_hi_hi = {loadUnit_maskInput_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_lo};
  wire [511:0]       loadUnit_maskInput_hi_hi_lo_hi = {loadUnit_maskInput_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_lo};
  wire [1023:0]      loadUnit_maskInput_hi_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_lo};
  wire [63:0]        _GEN_111 = {v0_225, v0_224};
  wire [63:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo = _GEN_111;
  wire [63:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo = _GEN_111;
  wire [63:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo = _GEN_111;
  wire [63:0]        _GEN_112 = {v0_227, v0_226};
  wire [63:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi = _GEN_112;
  wire [63:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi = _GEN_112;
  wire [63:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi = _GEN_112;
  wire [127:0]       loadUnit_maskInput_hi_hi_hi_lo_lo_lo = {loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo};
  wire [63:0]        _GEN_113 = {v0_229, v0_228};
  wire [63:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo = _GEN_113;
  wire [63:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo = _GEN_113;
  wire [63:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo = _GEN_113;
  wire [63:0]        _GEN_114 = {v0_231, v0_230};
  wire [63:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi = _GEN_114;
  wire [63:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi = _GEN_114;
  wire [63:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi = _GEN_114;
  wire [127:0]       loadUnit_maskInput_hi_hi_hi_lo_lo_hi = {loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]       loadUnit_maskInput_hi_hi_hi_lo_lo = {loadUnit_maskInput_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_lo};
  wire [63:0]        _GEN_115 = {v0_233, v0_232};
  wire [63:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo = _GEN_115;
  wire [63:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo = _GEN_115;
  wire [63:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo = _GEN_115;
  wire [63:0]        _GEN_116 = {v0_235, v0_234};
  wire [63:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi = _GEN_116;
  wire [63:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi = _GEN_116;
  wire [63:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi = _GEN_116;
  wire [127:0]       loadUnit_maskInput_hi_hi_hi_lo_hi_lo = {loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo};
  wire [63:0]        _GEN_117 = {v0_237, v0_236};
  wire [63:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo = _GEN_117;
  wire [63:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo = _GEN_117;
  wire [63:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo = _GEN_117;
  wire [63:0]        _GEN_118 = {v0_239, v0_238};
  wire [63:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi = _GEN_118;
  wire [63:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi = _GEN_118;
  wire [63:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi = _GEN_118;
  wire [127:0]       loadUnit_maskInput_hi_hi_hi_lo_hi_hi = {loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]       loadUnit_maskInput_hi_hi_hi_lo_hi = {loadUnit_maskInput_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_lo};
  wire [511:0]       loadUnit_maskInput_hi_hi_hi_lo = {loadUnit_maskInput_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_lo};
  wire [63:0]        _GEN_119 = {v0_241, v0_240};
  wire [63:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo = _GEN_119;
  wire [63:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo = _GEN_119;
  wire [63:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo = _GEN_119;
  wire [63:0]        _GEN_120 = {v0_243, v0_242};
  wire [63:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi = _GEN_120;
  wire [63:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi = _GEN_120;
  wire [63:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi = _GEN_120;
  wire [127:0]       loadUnit_maskInput_hi_hi_hi_hi_lo_lo = {loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo};
  wire [63:0]        _GEN_121 = {v0_245, v0_244};
  wire [63:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo = _GEN_121;
  wire [63:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo = _GEN_121;
  wire [63:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo = _GEN_121;
  wire [63:0]        _GEN_122 = {v0_247, v0_246};
  wire [63:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi = _GEN_122;
  wire [63:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi = _GEN_122;
  wire [63:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi = _GEN_122;
  wire [127:0]       loadUnit_maskInput_hi_hi_hi_hi_lo_hi = {loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]       loadUnit_maskInput_hi_hi_hi_hi_lo = {loadUnit_maskInput_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_lo};
  wire [63:0]        _GEN_123 = {v0_249, v0_248};
  wire [63:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo = _GEN_123;
  wire [63:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo = _GEN_123;
  wire [63:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo = _GEN_123;
  wire [63:0]        _GEN_124 = {v0_251, v0_250};
  wire [63:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi = _GEN_124;
  wire [63:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi = _GEN_124;
  wire [63:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi = _GEN_124;
  wire [127:0]       loadUnit_maskInput_hi_hi_hi_hi_hi_lo = {loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo};
  wire [63:0]        _GEN_125 = {v0_253, v0_252};
  wire [63:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo = _GEN_125;
  wire [63:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo = _GEN_125;
  wire [63:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo = _GEN_125;
  wire [63:0]        _GEN_126 = {v0_255, v0_254};
  wire [63:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi = _GEN_126;
  wire [63:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi = _GEN_126;
  wire [63:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi = _GEN_126;
  wire [127:0]       loadUnit_maskInput_hi_hi_hi_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]       loadUnit_maskInput_hi_hi_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_lo};
  wire [511:0]       loadUnit_maskInput_hi_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_lo};
  wire [1023:0]      loadUnit_maskInput_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_lo};
  wire [2047:0]      loadUnit_maskInput_hi_hi = {loadUnit_maskInput_hi_hi_hi, loadUnit_maskInput_hi_hi_lo};
  wire [4095:0]      loadUnit_maskInput_hi = {loadUnit_maskInput_hi_hi, loadUnit_maskInput_hi_lo};
  wire [511:0][15:0] _GEN_127 =
    {{loadUnit_maskInput_hi[4095:4080]},
     {loadUnit_maskInput_hi[4079:4064]},
     {loadUnit_maskInput_hi[4063:4048]},
     {loadUnit_maskInput_hi[4047:4032]},
     {loadUnit_maskInput_hi[4031:4016]},
     {loadUnit_maskInput_hi[4015:4000]},
     {loadUnit_maskInput_hi[3999:3984]},
     {loadUnit_maskInput_hi[3983:3968]},
     {loadUnit_maskInput_hi[3967:3952]},
     {loadUnit_maskInput_hi[3951:3936]},
     {loadUnit_maskInput_hi[3935:3920]},
     {loadUnit_maskInput_hi[3919:3904]},
     {loadUnit_maskInput_hi[3903:3888]},
     {loadUnit_maskInput_hi[3887:3872]},
     {loadUnit_maskInput_hi[3871:3856]},
     {loadUnit_maskInput_hi[3855:3840]},
     {loadUnit_maskInput_hi[3839:3824]},
     {loadUnit_maskInput_hi[3823:3808]},
     {loadUnit_maskInput_hi[3807:3792]},
     {loadUnit_maskInput_hi[3791:3776]},
     {loadUnit_maskInput_hi[3775:3760]},
     {loadUnit_maskInput_hi[3759:3744]},
     {loadUnit_maskInput_hi[3743:3728]},
     {loadUnit_maskInput_hi[3727:3712]},
     {loadUnit_maskInput_hi[3711:3696]},
     {loadUnit_maskInput_hi[3695:3680]},
     {loadUnit_maskInput_hi[3679:3664]},
     {loadUnit_maskInput_hi[3663:3648]},
     {loadUnit_maskInput_hi[3647:3632]},
     {loadUnit_maskInput_hi[3631:3616]},
     {loadUnit_maskInput_hi[3615:3600]},
     {loadUnit_maskInput_hi[3599:3584]},
     {loadUnit_maskInput_hi[3583:3568]},
     {loadUnit_maskInput_hi[3567:3552]},
     {loadUnit_maskInput_hi[3551:3536]},
     {loadUnit_maskInput_hi[3535:3520]},
     {loadUnit_maskInput_hi[3519:3504]},
     {loadUnit_maskInput_hi[3503:3488]},
     {loadUnit_maskInput_hi[3487:3472]},
     {loadUnit_maskInput_hi[3471:3456]},
     {loadUnit_maskInput_hi[3455:3440]},
     {loadUnit_maskInput_hi[3439:3424]},
     {loadUnit_maskInput_hi[3423:3408]},
     {loadUnit_maskInput_hi[3407:3392]},
     {loadUnit_maskInput_hi[3391:3376]},
     {loadUnit_maskInput_hi[3375:3360]},
     {loadUnit_maskInput_hi[3359:3344]},
     {loadUnit_maskInput_hi[3343:3328]},
     {loadUnit_maskInput_hi[3327:3312]},
     {loadUnit_maskInput_hi[3311:3296]},
     {loadUnit_maskInput_hi[3295:3280]},
     {loadUnit_maskInput_hi[3279:3264]},
     {loadUnit_maskInput_hi[3263:3248]},
     {loadUnit_maskInput_hi[3247:3232]},
     {loadUnit_maskInput_hi[3231:3216]},
     {loadUnit_maskInput_hi[3215:3200]},
     {loadUnit_maskInput_hi[3199:3184]},
     {loadUnit_maskInput_hi[3183:3168]},
     {loadUnit_maskInput_hi[3167:3152]},
     {loadUnit_maskInput_hi[3151:3136]},
     {loadUnit_maskInput_hi[3135:3120]},
     {loadUnit_maskInput_hi[3119:3104]},
     {loadUnit_maskInput_hi[3103:3088]},
     {loadUnit_maskInput_hi[3087:3072]},
     {loadUnit_maskInput_hi[3071:3056]},
     {loadUnit_maskInput_hi[3055:3040]},
     {loadUnit_maskInput_hi[3039:3024]},
     {loadUnit_maskInput_hi[3023:3008]},
     {loadUnit_maskInput_hi[3007:2992]},
     {loadUnit_maskInput_hi[2991:2976]},
     {loadUnit_maskInput_hi[2975:2960]},
     {loadUnit_maskInput_hi[2959:2944]},
     {loadUnit_maskInput_hi[2943:2928]},
     {loadUnit_maskInput_hi[2927:2912]},
     {loadUnit_maskInput_hi[2911:2896]},
     {loadUnit_maskInput_hi[2895:2880]},
     {loadUnit_maskInput_hi[2879:2864]},
     {loadUnit_maskInput_hi[2863:2848]},
     {loadUnit_maskInput_hi[2847:2832]},
     {loadUnit_maskInput_hi[2831:2816]},
     {loadUnit_maskInput_hi[2815:2800]},
     {loadUnit_maskInput_hi[2799:2784]},
     {loadUnit_maskInput_hi[2783:2768]},
     {loadUnit_maskInput_hi[2767:2752]},
     {loadUnit_maskInput_hi[2751:2736]},
     {loadUnit_maskInput_hi[2735:2720]},
     {loadUnit_maskInput_hi[2719:2704]},
     {loadUnit_maskInput_hi[2703:2688]},
     {loadUnit_maskInput_hi[2687:2672]},
     {loadUnit_maskInput_hi[2671:2656]},
     {loadUnit_maskInput_hi[2655:2640]},
     {loadUnit_maskInput_hi[2639:2624]},
     {loadUnit_maskInput_hi[2623:2608]},
     {loadUnit_maskInput_hi[2607:2592]},
     {loadUnit_maskInput_hi[2591:2576]},
     {loadUnit_maskInput_hi[2575:2560]},
     {loadUnit_maskInput_hi[2559:2544]},
     {loadUnit_maskInput_hi[2543:2528]},
     {loadUnit_maskInput_hi[2527:2512]},
     {loadUnit_maskInput_hi[2511:2496]},
     {loadUnit_maskInput_hi[2495:2480]},
     {loadUnit_maskInput_hi[2479:2464]},
     {loadUnit_maskInput_hi[2463:2448]},
     {loadUnit_maskInput_hi[2447:2432]},
     {loadUnit_maskInput_hi[2431:2416]},
     {loadUnit_maskInput_hi[2415:2400]},
     {loadUnit_maskInput_hi[2399:2384]},
     {loadUnit_maskInput_hi[2383:2368]},
     {loadUnit_maskInput_hi[2367:2352]},
     {loadUnit_maskInput_hi[2351:2336]},
     {loadUnit_maskInput_hi[2335:2320]},
     {loadUnit_maskInput_hi[2319:2304]},
     {loadUnit_maskInput_hi[2303:2288]},
     {loadUnit_maskInput_hi[2287:2272]},
     {loadUnit_maskInput_hi[2271:2256]},
     {loadUnit_maskInput_hi[2255:2240]},
     {loadUnit_maskInput_hi[2239:2224]},
     {loadUnit_maskInput_hi[2223:2208]},
     {loadUnit_maskInput_hi[2207:2192]},
     {loadUnit_maskInput_hi[2191:2176]},
     {loadUnit_maskInput_hi[2175:2160]},
     {loadUnit_maskInput_hi[2159:2144]},
     {loadUnit_maskInput_hi[2143:2128]},
     {loadUnit_maskInput_hi[2127:2112]},
     {loadUnit_maskInput_hi[2111:2096]},
     {loadUnit_maskInput_hi[2095:2080]},
     {loadUnit_maskInput_hi[2079:2064]},
     {loadUnit_maskInput_hi[2063:2048]},
     {loadUnit_maskInput_hi[2047:2032]},
     {loadUnit_maskInput_hi[2031:2016]},
     {loadUnit_maskInput_hi[2015:2000]},
     {loadUnit_maskInput_hi[1999:1984]},
     {loadUnit_maskInput_hi[1983:1968]},
     {loadUnit_maskInput_hi[1967:1952]},
     {loadUnit_maskInput_hi[1951:1936]},
     {loadUnit_maskInput_hi[1935:1920]},
     {loadUnit_maskInput_hi[1919:1904]},
     {loadUnit_maskInput_hi[1903:1888]},
     {loadUnit_maskInput_hi[1887:1872]},
     {loadUnit_maskInput_hi[1871:1856]},
     {loadUnit_maskInput_hi[1855:1840]},
     {loadUnit_maskInput_hi[1839:1824]},
     {loadUnit_maskInput_hi[1823:1808]},
     {loadUnit_maskInput_hi[1807:1792]},
     {loadUnit_maskInput_hi[1791:1776]},
     {loadUnit_maskInput_hi[1775:1760]},
     {loadUnit_maskInput_hi[1759:1744]},
     {loadUnit_maskInput_hi[1743:1728]},
     {loadUnit_maskInput_hi[1727:1712]},
     {loadUnit_maskInput_hi[1711:1696]},
     {loadUnit_maskInput_hi[1695:1680]},
     {loadUnit_maskInput_hi[1679:1664]},
     {loadUnit_maskInput_hi[1663:1648]},
     {loadUnit_maskInput_hi[1647:1632]},
     {loadUnit_maskInput_hi[1631:1616]},
     {loadUnit_maskInput_hi[1615:1600]},
     {loadUnit_maskInput_hi[1599:1584]},
     {loadUnit_maskInput_hi[1583:1568]},
     {loadUnit_maskInput_hi[1567:1552]},
     {loadUnit_maskInput_hi[1551:1536]},
     {loadUnit_maskInput_hi[1535:1520]},
     {loadUnit_maskInput_hi[1519:1504]},
     {loadUnit_maskInput_hi[1503:1488]},
     {loadUnit_maskInput_hi[1487:1472]},
     {loadUnit_maskInput_hi[1471:1456]},
     {loadUnit_maskInput_hi[1455:1440]},
     {loadUnit_maskInput_hi[1439:1424]},
     {loadUnit_maskInput_hi[1423:1408]},
     {loadUnit_maskInput_hi[1407:1392]},
     {loadUnit_maskInput_hi[1391:1376]},
     {loadUnit_maskInput_hi[1375:1360]},
     {loadUnit_maskInput_hi[1359:1344]},
     {loadUnit_maskInput_hi[1343:1328]},
     {loadUnit_maskInput_hi[1327:1312]},
     {loadUnit_maskInput_hi[1311:1296]},
     {loadUnit_maskInput_hi[1295:1280]},
     {loadUnit_maskInput_hi[1279:1264]},
     {loadUnit_maskInput_hi[1263:1248]},
     {loadUnit_maskInput_hi[1247:1232]},
     {loadUnit_maskInput_hi[1231:1216]},
     {loadUnit_maskInput_hi[1215:1200]},
     {loadUnit_maskInput_hi[1199:1184]},
     {loadUnit_maskInput_hi[1183:1168]},
     {loadUnit_maskInput_hi[1167:1152]},
     {loadUnit_maskInput_hi[1151:1136]},
     {loadUnit_maskInput_hi[1135:1120]},
     {loadUnit_maskInput_hi[1119:1104]},
     {loadUnit_maskInput_hi[1103:1088]},
     {loadUnit_maskInput_hi[1087:1072]},
     {loadUnit_maskInput_hi[1071:1056]},
     {loadUnit_maskInput_hi[1055:1040]},
     {loadUnit_maskInput_hi[1039:1024]},
     {loadUnit_maskInput_hi[1023:1008]},
     {loadUnit_maskInput_hi[1007:992]},
     {loadUnit_maskInput_hi[991:976]},
     {loadUnit_maskInput_hi[975:960]},
     {loadUnit_maskInput_hi[959:944]},
     {loadUnit_maskInput_hi[943:928]},
     {loadUnit_maskInput_hi[927:912]},
     {loadUnit_maskInput_hi[911:896]},
     {loadUnit_maskInput_hi[895:880]},
     {loadUnit_maskInput_hi[879:864]},
     {loadUnit_maskInput_hi[863:848]},
     {loadUnit_maskInput_hi[847:832]},
     {loadUnit_maskInput_hi[831:816]},
     {loadUnit_maskInput_hi[815:800]},
     {loadUnit_maskInput_hi[799:784]},
     {loadUnit_maskInput_hi[783:768]},
     {loadUnit_maskInput_hi[767:752]},
     {loadUnit_maskInput_hi[751:736]},
     {loadUnit_maskInput_hi[735:720]},
     {loadUnit_maskInput_hi[719:704]},
     {loadUnit_maskInput_hi[703:688]},
     {loadUnit_maskInput_hi[687:672]},
     {loadUnit_maskInput_hi[671:656]},
     {loadUnit_maskInput_hi[655:640]},
     {loadUnit_maskInput_hi[639:624]},
     {loadUnit_maskInput_hi[623:608]},
     {loadUnit_maskInput_hi[607:592]},
     {loadUnit_maskInput_hi[591:576]},
     {loadUnit_maskInput_hi[575:560]},
     {loadUnit_maskInput_hi[559:544]},
     {loadUnit_maskInput_hi[543:528]},
     {loadUnit_maskInput_hi[527:512]},
     {loadUnit_maskInput_hi[511:496]},
     {loadUnit_maskInput_hi[495:480]},
     {loadUnit_maskInput_hi[479:464]},
     {loadUnit_maskInput_hi[463:448]},
     {loadUnit_maskInput_hi[447:432]},
     {loadUnit_maskInput_hi[431:416]},
     {loadUnit_maskInput_hi[415:400]},
     {loadUnit_maskInput_hi[399:384]},
     {loadUnit_maskInput_hi[383:368]},
     {loadUnit_maskInput_hi[367:352]},
     {loadUnit_maskInput_hi[351:336]},
     {loadUnit_maskInput_hi[335:320]},
     {loadUnit_maskInput_hi[319:304]},
     {loadUnit_maskInput_hi[303:288]},
     {loadUnit_maskInput_hi[287:272]},
     {loadUnit_maskInput_hi[271:256]},
     {loadUnit_maskInput_hi[255:240]},
     {loadUnit_maskInput_hi[239:224]},
     {loadUnit_maskInput_hi[223:208]},
     {loadUnit_maskInput_hi[207:192]},
     {loadUnit_maskInput_hi[191:176]},
     {loadUnit_maskInput_hi[175:160]},
     {loadUnit_maskInput_hi[159:144]},
     {loadUnit_maskInput_hi[143:128]},
     {loadUnit_maskInput_hi[127:112]},
     {loadUnit_maskInput_hi[111:96]},
     {loadUnit_maskInput_hi[95:80]},
     {loadUnit_maskInput_hi[79:64]},
     {loadUnit_maskInput_hi[63:48]},
     {loadUnit_maskInput_hi[47:32]},
     {loadUnit_maskInput_hi[31:16]},
     {loadUnit_maskInput_hi[15:0]},
     {loadUnit_maskInput_lo[4095:4080]},
     {loadUnit_maskInput_lo[4079:4064]},
     {loadUnit_maskInput_lo[4063:4048]},
     {loadUnit_maskInput_lo[4047:4032]},
     {loadUnit_maskInput_lo[4031:4016]},
     {loadUnit_maskInput_lo[4015:4000]},
     {loadUnit_maskInput_lo[3999:3984]},
     {loadUnit_maskInput_lo[3983:3968]},
     {loadUnit_maskInput_lo[3967:3952]},
     {loadUnit_maskInput_lo[3951:3936]},
     {loadUnit_maskInput_lo[3935:3920]},
     {loadUnit_maskInput_lo[3919:3904]},
     {loadUnit_maskInput_lo[3903:3888]},
     {loadUnit_maskInput_lo[3887:3872]},
     {loadUnit_maskInput_lo[3871:3856]},
     {loadUnit_maskInput_lo[3855:3840]},
     {loadUnit_maskInput_lo[3839:3824]},
     {loadUnit_maskInput_lo[3823:3808]},
     {loadUnit_maskInput_lo[3807:3792]},
     {loadUnit_maskInput_lo[3791:3776]},
     {loadUnit_maskInput_lo[3775:3760]},
     {loadUnit_maskInput_lo[3759:3744]},
     {loadUnit_maskInput_lo[3743:3728]},
     {loadUnit_maskInput_lo[3727:3712]},
     {loadUnit_maskInput_lo[3711:3696]},
     {loadUnit_maskInput_lo[3695:3680]},
     {loadUnit_maskInput_lo[3679:3664]},
     {loadUnit_maskInput_lo[3663:3648]},
     {loadUnit_maskInput_lo[3647:3632]},
     {loadUnit_maskInput_lo[3631:3616]},
     {loadUnit_maskInput_lo[3615:3600]},
     {loadUnit_maskInput_lo[3599:3584]},
     {loadUnit_maskInput_lo[3583:3568]},
     {loadUnit_maskInput_lo[3567:3552]},
     {loadUnit_maskInput_lo[3551:3536]},
     {loadUnit_maskInput_lo[3535:3520]},
     {loadUnit_maskInput_lo[3519:3504]},
     {loadUnit_maskInput_lo[3503:3488]},
     {loadUnit_maskInput_lo[3487:3472]},
     {loadUnit_maskInput_lo[3471:3456]},
     {loadUnit_maskInput_lo[3455:3440]},
     {loadUnit_maskInput_lo[3439:3424]},
     {loadUnit_maskInput_lo[3423:3408]},
     {loadUnit_maskInput_lo[3407:3392]},
     {loadUnit_maskInput_lo[3391:3376]},
     {loadUnit_maskInput_lo[3375:3360]},
     {loadUnit_maskInput_lo[3359:3344]},
     {loadUnit_maskInput_lo[3343:3328]},
     {loadUnit_maskInput_lo[3327:3312]},
     {loadUnit_maskInput_lo[3311:3296]},
     {loadUnit_maskInput_lo[3295:3280]},
     {loadUnit_maskInput_lo[3279:3264]},
     {loadUnit_maskInput_lo[3263:3248]},
     {loadUnit_maskInput_lo[3247:3232]},
     {loadUnit_maskInput_lo[3231:3216]},
     {loadUnit_maskInput_lo[3215:3200]},
     {loadUnit_maskInput_lo[3199:3184]},
     {loadUnit_maskInput_lo[3183:3168]},
     {loadUnit_maskInput_lo[3167:3152]},
     {loadUnit_maskInput_lo[3151:3136]},
     {loadUnit_maskInput_lo[3135:3120]},
     {loadUnit_maskInput_lo[3119:3104]},
     {loadUnit_maskInput_lo[3103:3088]},
     {loadUnit_maskInput_lo[3087:3072]},
     {loadUnit_maskInput_lo[3071:3056]},
     {loadUnit_maskInput_lo[3055:3040]},
     {loadUnit_maskInput_lo[3039:3024]},
     {loadUnit_maskInput_lo[3023:3008]},
     {loadUnit_maskInput_lo[3007:2992]},
     {loadUnit_maskInput_lo[2991:2976]},
     {loadUnit_maskInput_lo[2975:2960]},
     {loadUnit_maskInput_lo[2959:2944]},
     {loadUnit_maskInput_lo[2943:2928]},
     {loadUnit_maskInput_lo[2927:2912]},
     {loadUnit_maskInput_lo[2911:2896]},
     {loadUnit_maskInput_lo[2895:2880]},
     {loadUnit_maskInput_lo[2879:2864]},
     {loadUnit_maskInput_lo[2863:2848]},
     {loadUnit_maskInput_lo[2847:2832]},
     {loadUnit_maskInput_lo[2831:2816]},
     {loadUnit_maskInput_lo[2815:2800]},
     {loadUnit_maskInput_lo[2799:2784]},
     {loadUnit_maskInput_lo[2783:2768]},
     {loadUnit_maskInput_lo[2767:2752]},
     {loadUnit_maskInput_lo[2751:2736]},
     {loadUnit_maskInput_lo[2735:2720]},
     {loadUnit_maskInput_lo[2719:2704]},
     {loadUnit_maskInput_lo[2703:2688]},
     {loadUnit_maskInput_lo[2687:2672]},
     {loadUnit_maskInput_lo[2671:2656]},
     {loadUnit_maskInput_lo[2655:2640]},
     {loadUnit_maskInput_lo[2639:2624]},
     {loadUnit_maskInput_lo[2623:2608]},
     {loadUnit_maskInput_lo[2607:2592]},
     {loadUnit_maskInput_lo[2591:2576]},
     {loadUnit_maskInput_lo[2575:2560]},
     {loadUnit_maskInput_lo[2559:2544]},
     {loadUnit_maskInput_lo[2543:2528]},
     {loadUnit_maskInput_lo[2527:2512]},
     {loadUnit_maskInput_lo[2511:2496]},
     {loadUnit_maskInput_lo[2495:2480]},
     {loadUnit_maskInput_lo[2479:2464]},
     {loadUnit_maskInput_lo[2463:2448]},
     {loadUnit_maskInput_lo[2447:2432]},
     {loadUnit_maskInput_lo[2431:2416]},
     {loadUnit_maskInput_lo[2415:2400]},
     {loadUnit_maskInput_lo[2399:2384]},
     {loadUnit_maskInput_lo[2383:2368]},
     {loadUnit_maskInput_lo[2367:2352]},
     {loadUnit_maskInput_lo[2351:2336]},
     {loadUnit_maskInput_lo[2335:2320]},
     {loadUnit_maskInput_lo[2319:2304]},
     {loadUnit_maskInput_lo[2303:2288]},
     {loadUnit_maskInput_lo[2287:2272]},
     {loadUnit_maskInput_lo[2271:2256]},
     {loadUnit_maskInput_lo[2255:2240]},
     {loadUnit_maskInput_lo[2239:2224]},
     {loadUnit_maskInput_lo[2223:2208]},
     {loadUnit_maskInput_lo[2207:2192]},
     {loadUnit_maskInput_lo[2191:2176]},
     {loadUnit_maskInput_lo[2175:2160]},
     {loadUnit_maskInput_lo[2159:2144]},
     {loadUnit_maskInput_lo[2143:2128]},
     {loadUnit_maskInput_lo[2127:2112]},
     {loadUnit_maskInput_lo[2111:2096]},
     {loadUnit_maskInput_lo[2095:2080]},
     {loadUnit_maskInput_lo[2079:2064]},
     {loadUnit_maskInput_lo[2063:2048]},
     {loadUnit_maskInput_lo[2047:2032]},
     {loadUnit_maskInput_lo[2031:2016]},
     {loadUnit_maskInput_lo[2015:2000]},
     {loadUnit_maskInput_lo[1999:1984]},
     {loadUnit_maskInput_lo[1983:1968]},
     {loadUnit_maskInput_lo[1967:1952]},
     {loadUnit_maskInput_lo[1951:1936]},
     {loadUnit_maskInput_lo[1935:1920]},
     {loadUnit_maskInput_lo[1919:1904]},
     {loadUnit_maskInput_lo[1903:1888]},
     {loadUnit_maskInput_lo[1887:1872]},
     {loadUnit_maskInput_lo[1871:1856]},
     {loadUnit_maskInput_lo[1855:1840]},
     {loadUnit_maskInput_lo[1839:1824]},
     {loadUnit_maskInput_lo[1823:1808]},
     {loadUnit_maskInput_lo[1807:1792]},
     {loadUnit_maskInput_lo[1791:1776]},
     {loadUnit_maskInput_lo[1775:1760]},
     {loadUnit_maskInput_lo[1759:1744]},
     {loadUnit_maskInput_lo[1743:1728]},
     {loadUnit_maskInput_lo[1727:1712]},
     {loadUnit_maskInput_lo[1711:1696]},
     {loadUnit_maskInput_lo[1695:1680]},
     {loadUnit_maskInput_lo[1679:1664]},
     {loadUnit_maskInput_lo[1663:1648]},
     {loadUnit_maskInput_lo[1647:1632]},
     {loadUnit_maskInput_lo[1631:1616]},
     {loadUnit_maskInput_lo[1615:1600]},
     {loadUnit_maskInput_lo[1599:1584]},
     {loadUnit_maskInput_lo[1583:1568]},
     {loadUnit_maskInput_lo[1567:1552]},
     {loadUnit_maskInput_lo[1551:1536]},
     {loadUnit_maskInput_lo[1535:1520]},
     {loadUnit_maskInput_lo[1519:1504]},
     {loadUnit_maskInput_lo[1503:1488]},
     {loadUnit_maskInput_lo[1487:1472]},
     {loadUnit_maskInput_lo[1471:1456]},
     {loadUnit_maskInput_lo[1455:1440]},
     {loadUnit_maskInput_lo[1439:1424]},
     {loadUnit_maskInput_lo[1423:1408]},
     {loadUnit_maskInput_lo[1407:1392]},
     {loadUnit_maskInput_lo[1391:1376]},
     {loadUnit_maskInput_lo[1375:1360]},
     {loadUnit_maskInput_lo[1359:1344]},
     {loadUnit_maskInput_lo[1343:1328]},
     {loadUnit_maskInput_lo[1327:1312]},
     {loadUnit_maskInput_lo[1311:1296]},
     {loadUnit_maskInput_lo[1295:1280]},
     {loadUnit_maskInput_lo[1279:1264]},
     {loadUnit_maskInput_lo[1263:1248]},
     {loadUnit_maskInput_lo[1247:1232]},
     {loadUnit_maskInput_lo[1231:1216]},
     {loadUnit_maskInput_lo[1215:1200]},
     {loadUnit_maskInput_lo[1199:1184]},
     {loadUnit_maskInput_lo[1183:1168]},
     {loadUnit_maskInput_lo[1167:1152]},
     {loadUnit_maskInput_lo[1151:1136]},
     {loadUnit_maskInput_lo[1135:1120]},
     {loadUnit_maskInput_lo[1119:1104]},
     {loadUnit_maskInput_lo[1103:1088]},
     {loadUnit_maskInput_lo[1087:1072]},
     {loadUnit_maskInput_lo[1071:1056]},
     {loadUnit_maskInput_lo[1055:1040]},
     {loadUnit_maskInput_lo[1039:1024]},
     {loadUnit_maskInput_lo[1023:1008]},
     {loadUnit_maskInput_lo[1007:992]},
     {loadUnit_maskInput_lo[991:976]},
     {loadUnit_maskInput_lo[975:960]},
     {loadUnit_maskInput_lo[959:944]},
     {loadUnit_maskInput_lo[943:928]},
     {loadUnit_maskInput_lo[927:912]},
     {loadUnit_maskInput_lo[911:896]},
     {loadUnit_maskInput_lo[895:880]},
     {loadUnit_maskInput_lo[879:864]},
     {loadUnit_maskInput_lo[863:848]},
     {loadUnit_maskInput_lo[847:832]},
     {loadUnit_maskInput_lo[831:816]},
     {loadUnit_maskInput_lo[815:800]},
     {loadUnit_maskInput_lo[799:784]},
     {loadUnit_maskInput_lo[783:768]},
     {loadUnit_maskInput_lo[767:752]},
     {loadUnit_maskInput_lo[751:736]},
     {loadUnit_maskInput_lo[735:720]},
     {loadUnit_maskInput_lo[719:704]},
     {loadUnit_maskInput_lo[703:688]},
     {loadUnit_maskInput_lo[687:672]},
     {loadUnit_maskInput_lo[671:656]},
     {loadUnit_maskInput_lo[655:640]},
     {loadUnit_maskInput_lo[639:624]},
     {loadUnit_maskInput_lo[623:608]},
     {loadUnit_maskInput_lo[607:592]},
     {loadUnit_maskInput_lo[591:576]},
     {loadUnit_maskInput_lo[575:560]},
     {loadUnit_maskInput_lo[559:544]},
     {loadUnit_maskInput_lo[543:528]},
     {loadUnit_maskInput_lo[527:512]},
     {loadUnit_maskInput_lo[511:496]},
     {loadUnit_maskInput_lo[495:480]},
     {loadUnit_maskInput_lo[479:464]},
     {loadUnit_maskInput_lo[463:448]},
     {loadUnit_maskInput_lo[447:432]},
     {loadUnit_maskInput_lo[431:416]},
     {loadUnit_maskInput_lo[415:400]},
     {loadUnit_maskInput_lo[399:384]},
     {loadUnit_maskInput_lo[383:368]},
     {loadUnit_maskInput_lo[367:352]},
     {loadUnit_maskInput_lo[351:336]},
     {loadUnit_maskInput_lo[335:320]},
     {loadUnit_maskInput_lo[319:304]},
     {loadUnit_maskInput_lo[303:288]},
     {loadUnit_maskInput_lo[287:272]},
     {loadUnit_maskInput_lo[271:256]},
     {loadUnit_maskInput_lo[255:240]},
     {loadUnit_maskInput_lo[239:224]},
     {loadUnit_maskInput_lo[223:208]},
     {loadUnit_maskInput_lo[207:192]},
     {loadUnit_maskInput_lo[191:176]},
     {loadUnit_maskInput_lo[175:160]},
     {loadUnit_maskInput_lo[159:144]},
     {loadUnit_maskInput_lo[143:128]},
     {loadUnit_maskInput_lo[127:112]},
     {loadUnit_maskInput_lo[111:96]},
     {loadUnit_maskInput_lo[95:80]},
     {loadUnit_maskInput_lo[79:64]},
     {loadUnit_maskInput_lo[63:48]},
     {loadUnit_maskInput_lo[47:32]},
     {loadUnit_maskInput_lo[31:16]},
     {loadUnit_maskInput_lo[15:0]}};
  wire [8:0]         maskSelect_1 = _storeUnit_maskSelect_valid ? _storeUnit_maskSelect_bits : 9'h0;
  wire [127:0]       storeUnit_maskInput_lo_lo_lo_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_lo_lo_lo_lo_hi = {storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]       storeUnit_maskInput_lo_lo_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_lo_lo_lo_hi_lo = {storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_lo_lo_lo_hi_hi = {storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]       storeUnit_maskInput_lo_lo_lo_lo_hi = {storeUnit_maskInput_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_lo};
  wire [511:0]       storeUnit_maskInput_lo_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_lo_lo_hi_lo_lo = {storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_lo_lo_hi_lo_hi = {storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]       storeUnit_maskInput_lo_lo_lo_hi_lo = {storeUnit_maskInput_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_lo_lo_hi_hi_lo = {storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_lo_lo_hi_hi_hi = {storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]       storeUnit_maskInput_lo_lo_lo_hi_hi = {storeUnit_maskInput_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_lo};
  wire [511:0]       storeUnit_maskInput_lo_lo_lo_hi = {storeUnit_maskInput_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_lo};
  wire [1023:0]      storeUnit_maskInput_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_lo_hi_lo_lo_lo = {storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_lo_hi_lo_lo_hi = {storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]       storeUnit_maskInput_lo_lo_hi_lo_lo = {storeUnit_maskInput_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_lo_hi_lo_hi_lo = {storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_lo_hi_lo_hi_hi = {storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]       storeUnit_maskInput_lo_lo_hi_lo_hi = {storeUnit_maskInput_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_lo};
  wire [511:0]       storeUnit_maskInput_lo_lo_hi_lo = {storeUnit_maskInput_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_lo_hi_hi_lo_lo = {storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_lo_hi_hi_lo_hi = {storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]       storeUnit_maskInput_lo_lo_hi_hi_lo = {storeUnit_maskInput_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_lo_hi_hi_hi_lo = {storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_lo_hi_hi_hi_hi = {storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]       storeUnit_maskInput_lo_lo_hi_hi_hi = {storeUnit_maskInput_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_lo};
  wire [511:0]       storeUnit_maskInput_lo_lo_hi_hi = {storeUnit_maskInput_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_lo};
  wire [1023:0]      storeUnit_maskInput_lo_lo_hi = {storeUnit_maskInput_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo};
  wire [2047:0]      storeUnit_maskInput_lo_lo = {storeUnit_maskInput_lo_lo_hi, storeUnit_maskInput_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_hi_lo_lo_lo_lo = {storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_hi_lo_lo_lo_hi = {storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]       storeUnit_maskInput_lo_hi_lo_lo_lo = {storeUnit_maskInput_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_hi_lo_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_hi_lo_lo_hi_hi = {storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]       storeUnit_maskInput_lo_hi_lo_lo_hi = {storeUnit_maskInput_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_lo};
  wire [511:0]       storeUnit_maskInput_lo_hi_lo_lo = {storeUnit_maskInput_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_hi_lo_hi_lo_lo = {storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_hi_lo_hi_lo_hi = {storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]       storeUnit_maskInput_lo_hi_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_hi_lo_hi_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_hi_lo_hi_hi_hi = {storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]       storeUnit_maskInput_lo_hi_lo_hi_hi = {storeUnit_maskInput_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_lo};
  wire [511:0]       storeUnit_maskInput_lo_hi_lo_hi = {storeUnit_maskInput_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_lo};
  wire [1023:0]      storeUnit_maskInput_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_hi_hi_lo_lo_lo = {storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_hi_hi_lo_lo_hi = {storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]       storeUnit_maskInput_lo_hi_hi_lo_lo = {storeUnit_maskInput_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_hi_hi_lo_hi_lo = {storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_hi_hi_lo_hi_hi = {storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]       storeUnit_maskInput_lo_hi_hi_lo_hi = {storeUnit_maskInput_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_lo};
  wire [511:0]       storeUnit_maskInput_lo_hi_hi_lo = {storeUnit_maskInput_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_hi_hi_hi_lo_lo = {storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_hi_hi_hi_lo_hi = {storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]       storeUnit_maskInput_lo_hi_hi_hi_lo = {storeUnit_maskInput_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_hi_hi_hi_hi_lo = {storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_lo_hi_hi_hi_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]       storeUnit_maskInput_lo_hi_hi_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_lo};
  wire [511:0]       storeUnit_maskInput_lo_hi_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_lo};
  wire [1023:0]      storeUnit_maskInput_lo_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_lo};
  wire [2047:0]      storeUnit_maskInput_lo_hi = {storeUnit_maskInput_lo_hi_hi, storeUnit_maskInput_lo_hi_lo};
  wire [4095:0]      storeUnit_maskInput_lo = {storeUnit_maskInput_lo_hi, storeUnit_maskInput_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_lo_lo_lo_lo_lo = {storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_lo_lo_lo_lo_hi = {storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]       storeUnit_maskInput_hi_lo_lo_lo_lo = {storeUnit_maskInput_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_lo_lo_lo_hi_lo = {storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_lo_lo_lo_hi_hi = {storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]       storeUnit_maskInput_hi_lo_lo_lo_hi = {storeUnit_maskInput_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_lo};
  wire [511:0]       storeUnit_maskInput_hi_lo_lo_lo = {storeUnit_maskInput_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_lo_lo_hi_lo_lo = {storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_lo_lo_hi_lo_hi = {storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]       storeUnit_maskInput_hi_lo_lo_hi_lo = {storeUnit_maskInput_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_lo_lo_hi_hi_lo = {storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_lo_lo_hi_hi_hi = {storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]       storeUnit_maskInput_hi_lo_lo_hi_hi = {storeUnit_maskInput_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_lo};
  wire [511:0]       storeUnit_maskInput_hi_lo_lo_hi = {storeUnit_maskInput_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_lo};
  wire [1023:0]      storeUnit_maskInput_hi_lo_lo = {storeUnit_maskInput_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_lo_hi_lo_lo_lo = {storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_lo_hi_lo_lo_hi = {storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]       storeUnit_maskInput_hi_lo_hi_lo_lo = {storeUnit_maskInput_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_lo_hi_lo_hi_lo = {storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_lo_hi_lo_hi_hi = {storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]       storeUnit_maskInput_hi_lo_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_lo};
  wire [511:0]       storeUnit_maskInput_hi_lo_hi_lo = {storeUnit_maskInput_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_lo_hi_hi_lo_lo = {storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_lo_hi_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]       storeUnit_maskInput_hi_lo_hi_hi_lo = {storeUnit_maskInput_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_lo_hi_hi_hi_lo = {storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_lo_hi_hi_hi_hi = {storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]       storeUnit_maskInput_hi_lo_hi_hi_hi = {storeUnit_maskInput_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_lo};
  wire [511:0]       storeUnit_maskInput_hi_lo_hi_hi = {storeUnit_maskInput_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_lo};
  wire [1023:0]      storeUnit_maskInput_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo};
  wire [2047:0]      storeUnit_maskInput_hi_lo = {storeUnit_maskInput_hi_lo_hi, storeUnit_maskInput_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_hi_lo_lo_lo_lo = {storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_hi_lo_lo_lo_hi = {storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]       storeUnit_maskInput_hi_hi_lo_lo_lo = {storeUnit_maskInput_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_hi_lo_lo_hi_lo = {storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_hi_lo_lo_hi_hi = {storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]       storeUnit_maskInput_hi_hi_lo_lo_hi = {storeUnit_maskInput_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_lo};
  wire [511:0]       storeUnit_maskInput_hi_hi_lo_lo = {storeUnit_maskInput_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_hi_lo_hi_lo_lo = {storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_hi_lo_hi_lo_hi = {storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]       storeUnit_maskInput_hi_hi_lo_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_hi_lo_hi_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_hi_lo_hi_hi_hi = {storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]       storeUnit_maskInput_hi_hi_lo_hi_hi = {storeUnit_maskInput_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_lo};
  wire [511:0]       storeUnit_maskInput_hi_hi_lo_hi = {storeUnit_maskInput_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_lo};
  wire [1023:0]      storeUnit_maskInput_hi_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_hi_hi_lo_lo_lo = {storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_hi_hi_lo_lo_hi = {storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]       storeUnit_maskInput_hi_hi_hi_lo_lo = {storeUnit_maskInput_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_hi_hi_lo_hi_lo = {storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_hi_hi_lo_hi_hi = {storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]       storeUnit_maskInput_hi_hi_hi_lo_hi = {storeUnit_maskInput_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_lo};
  wire [511:0]       storeUnit_maskInput_hi_hi_hi_lo = {storeUnit_maskInput_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_hi_hi_hi_lo_lo = {storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_hi_hi_hi_lo_hi = {storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]       storeUnit_maskInput_hi_hi_hi_hi_lo = {storeUnit_maskInput_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_hi_hi_hi_hi_lo = {storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]       storeUnit_maskInput_hi_hi_hi_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]       storeUnit_maskInput_hi_hi_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_lo};
  wire [511:0]       storeUnit_maskInput_hi_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_lo};
  wire [1023:0]      storeUnit_maskInput_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_lo};
  wire [2047:0]      storeUnit_maskInput_hi_hi = {storeUnit_maskInput_hi_hi_hi, storeUnit_maskInput_hi_hi_lo};
  wire [4095:0]      storeUnit_maskInput_hi = {storeUnit_maskInput_hi_hi, storeUnit_maskInput_hi_lo};
  wire [511:0][15:0] _GEN_128 =
    {{storeUnit_maskInput_hi[4095:4080]},
     {storeUnit_maskInput_hi[4079:4064]},
     {storeUnit_maskInput_hi[4063:4048]},
     {storeUnit_maskInput_hi[4047:4032]},
     {storeUnit_maskInput_hi[4031:4016]},
     {storeUnit_maskInput_hi[4015:4000]},
     {storeUnit_maskInput_hi[3999:3984]},
     {storeUnit_maskInput_hi[3983:3968]},
     {storeUnit_maskInput_hi[3967:3952]},
     {storeUnit_maskInput_hi[3951:3936]},
     {storeUnit_maskInput_hi[3935:3920]},
     {storeUnit_maskInput_hi[3919:3904]},
     {storeUnit_maskInput_hi[3903:3888]},
     {storeUnit_maskInput_hi[3887:3872]},
     {storeUnit_maskInput_hi[3871:3856]},
     {storeUnit_maskInput_hi[3855:3840]},
     {storeUnit_maskInput_hi[3839:3824]},
     {storeUnit_maskInput_hi[3823:3808]},
     {storeUnit_maskInput_hi[3807:3792]},
     {storeUnit_maskInput_hi[3791:3776]},
     {storeUnit_maskInput_hi[3775:3760]},
     {storeUnit_maskInput_hi[3759:3744]},
     {storeUnit_maskInput_hi[3743:3728]},
     {storeUnit_maskInput_hi[3727:3712]},
     {storeUnit_maskInput_hi[3711:3696]},
     {storeUnit_maskInput_hi[3695:3680]},
     {storeUnit_maskInput_hi[3679:3664]},
     {storeUnit_maskInput_hi[3663:3648]},
     {storeUnit_maskInput_hi[3647:3632]},
     {storeUnit_maskInput_hi[3631:3616]},
     {storeUnit_maskInput_hi[3615:3600]},
     {storeUnit_maskInput_hi[3599:3584]},
     {storeUnit_maskInput_hi[3583:3568]},
     {storeUnit_maskInput_hi[3567:3552]},
     {storeUnit_maskInput_hi[3551:3536]},
     {storeUnit_maskInput_hi[3535:3520]},
     {storeUnit_maskInput_hi[3519:3504]},
     {storeUnit_maskInput_hi[3503:3488]},
     {storeUnit_maskInput_hi[3487:3472]},
     {storeUnit_maskInput_hi[3471:3456]},
     {storeUnit_maskInput_hi[3455:3440]},
     {storeUnit_maskInput_hi[3439:3424]},
     {storeUnit_maskInput_hi[3423:3408]},
     {storeUnit_maskInput_hi[3407:3392]},
     {storeUnit_maskInput_hi[3391:3376]},
     {storeUnit_maskInput_hi[3375:3360]},
     {storeUnit_maskInput_hi[3359:3344]},
     {storeUnit_maskInput_hi[3343:3328]},
     {storeUnit_maskInput_hi[3327:3312]},
     {storeUnit_maskInput_hi[3311:3296]},
     {storeUnit_maskInput_hi[3295:3280]},
     {storeUnit_maskInput_hi[3279:3264]},
     {storeUnit_maskInput_hi[3263:3248]},
     {storeUnit_maskInput_hi[3247:3232]},
     {storeUnit_maskInput_hi[3231:3216]},
     {storeUnit_maskInput_hi[3215:3200]},
     {storeUnit_maskInput_hi[3199:3184]},
     {storeUnit_maskInput_hi[3183:3168]},
     {storeUnit_maskInput_hi[3167:3152]},
     {storeUnit_maskInput_hi[3151:3136]},
     {storeUnit_maskInput_hi[3135:3120]},
     {storeUnit_maskInput_hi[3119:3104]},
     {storeUnit_maskInput_hi[3103:3088]},
     {storeUnit_maskInput_hi[3087:3072]},
     {storeUnit_maskInput_hi[3071:3056]},
     {storeUnit_maskInput_hi[3055:3040]},
     {storeUnit_maskInput_hi[3039:3024]},
     {storeUnit_maskInput_hi[3023:3008]},
     {storeUnit_maskInput_hi[3007:2992]},
     {storeUnit_maskInput_hi[2991:2976]},
     {storeUnit_maskInput_hi[2975:2960]},
     {storeUnit_maskInput_hi[2959:2944]},
     {storeUnit_maskInput_hi[2943:2928]},
     {storeUnit_maskInput_hi[2927:2912]},
     {storeUnit_maskInput_hi[2911:2896]},
     {storeUnit_maskInput_hi[2895:2880]},
     {storeUnit_maskInput_hi[2879:2864]},
     {storeUnit_maskInput_hi[2863:2848]},
     {storeUnit_maskInput_hi[2847:2832]},
     {storeUnit_maskInput_hi[2831:2816]},
     {storeUnit_maskInput_hi[2815:2800]},
     {storeUnit_maskInput_hi[2799:2784]},
     {storeUnit_maskInput_hi[2783:2768]},
     {storeUnit_maskInput_hi[2767:2752]},
     {storeUnit_maskInput_hi[2751:2736]},
     {storeUnit_maskInput_hi[2735:2720]},
     {storeUnit_maskInput_hi[2719:2704]},
     {storeUnit_maskInput_hi[2703:2688]},
     {storeUnit_maskInput_hi[2687:2672]},
     {storeUnit_maskInput_hi[2671:2656]},
     {storeUnit_maskInput_hi[2655:2640]},
     {storeUnit_maskInput_hi[2639:2624]},
     {storeUnit_maskInput_hi[2623:2608]},
     {storeUnit_maskInput_hi[2607:2592]},
     {storeUnit_maskInput_hi[2591:2576]},
     {storeUnit_maskInput_hi[2575:2560]},
     {storeUnit_maskInput_hi[2559:2544]},
     {storeUnit_maskInput_hi[2543:2528]},
     {storeUnit_maskInput_hi[2527:2512]},
     {storeUnit_maskInput_hi[2511:2496]},
     {storeUnit_maskInput_hi[2495:2480]},
     {storeUnit_maskInput_hi[2479:2464]},
     {storeUnit_maskInput_hi[2463:2448]},
     {storeUnit_maskInput_hi[2447:2432]},
     {storeUnit_maskInput_hi[2431:2416]},
     {storeUnit_maskInput_hi[2415:2400]},
     {storeUnit_maskInput_hi[2399:2384]},
     {storeUnit_maskInput_hi[2383:2368]},
     {storeUnit_maskInput_hi[2367:2352]},
     {storeUnit_maskInput_hi[2351:2336]},
     {storeUnit_maskInput_hi[2335:2320]},
     {storeUnit_maskInput_hi[2319:2304]},
     {storeUnit_maskInput_hi[2303:2288]},
     {storeUnit_maskInput_hi[2287:2272]},
     {storeUnit_maskInput_hi[2271:2256]},
     {storeUnit_maskInput_hi[2255:2240]},
     {storeUnit_maskInput_hi[2239:2224]},
     {storeUnit_maskInput_hi[2223:2208]},
     {storeUnit_maskInput_hi[2207:2192]},
     {storeUnit_maskInput_hi[2191:2176]},
     {storeUnit_maskInput_hi[2175:2160]},
     {storeUnit_maskInput_hi[2159:2144]},
     {storeUnit_maskInput_hi[2143:2128]},
     {storeUnit_maskInput_hi[2127:2112]},
     {storeUnit_maskInput_hi[2111:2096]},
     {storeUnit_maskInput_hi[2095:2080]},
     {storeUnit_maskInput_hi[2079:2064]},
     {storeUnit_maskInput_hi[2063:2048]},
     {storeUnit_maskInput_hi[2047:2032]},
     {storeUnit_maskInput_hi[2031:2016]},
     {storeUnit_maskInput_hi[2015:2000]},
     {storeUnit_maskInput_hi[1999:1984]},
     {storeUnit_maskInput_hi[1983:1968]},
     {storeUnit_maskInput_hi[1967:1952]},
     {storeUnit_maskInput_hi[1951:1936]},
     {storeUnit_maskInput_hi[1935:1920]},
     {storeUnit_maskInput_hi[1919:1904]},
     {storeUnit_maskInput_hi[1903:1888]},
     {storeUnit_maskInput_hi[1887:1872]},
     {storeUnit_maskInput_hi[1871:1856]},
     {storeUnit_maskInput_hi[1855:1840]},
     {storeUnit_maskInput_hi[1839:1824]},
     {storeUnit_maskInput_hi[1823:1808]},
     {storeUnit_maskInput_hi[1807:1792]},
     {storeUnit_maskInput_hi[1791:1776]},
     {storeUnit_maskInput_hi[1775:1760]},
     {storeUnit_maskInput_hi[1759:1744]},
     {storeUnit_maskInput_hi[1743:1728]},
     {storeUnit_maskInput_hi[1727:1712]},
     {storeUnit_maskInput_hi[1711:1696]},
     {storeUnit_maskInput_hi[1695:1680]},
     {storeUnit_maskInput_hi[1679:1664]},
     {storeUnit_maskInput_hi[1663:1648]},
     {storeUnit_maskInput_hi[1647:1632]},
     {storeUnit_maskInput_hi[1631:1616]},
     {storeUnit_maskInput_hi[1615:1600]},
     {storeUnit_maskInput_hi[1599:1584]},
     {storeUnit_maskInput_hi[1583:1568]},
     {storeUnit_maskInput_hi[1567:1552]},
     {storeUnit_maskInput_hi[1551:1536]},
     {storeUnit_maskInput_hi[1535:1520]},
     {storeUnit_maskInput_hi[1519:1504]},
     {storeUnit_maskInput_hi[1503:1488]},
     {storeUnit_maskInput_hi[1487:1472]},
     {storeUnit_maskInput_hi[1471:1456]},
     {storeUnit_maskInput_hi[1455:1440]},
     {storeUnit_maskInput_hi[1439:1424]},
     {storeUnit_maskInput_hi[1423:1408]},
     {storeUnit_maskInput_hi[1407:1392]},
     {storeUnit_maskInput_hi[1391:1376]},
     {storeUnit_maskInput_hi[1375:1360]},
     {storeUnit_maskInput_hi[1359:1344]},
     {storeUnit_maskInput_hi[1343:1328]},
     {storeUnit_maskInput_hi[1327:1312]},
     {storeUnit_maskInput_hi[1311:1296]},
     {storeUnit_maskInput_hi[1295:1280]},
     {storeUnit_maskInput_hi[1279:1264]},
     {storeUnit_maskInput_hi[1263:1248]},
     {storeUnit_maskInput_hi[1247:1232]},
     {storeUnit_maskInput_hi[1231:1216]},
     {storeUnit_maskInput_hi[1215:1200]},
     {storeUnit_maskInput_hi[1199:1184]},
     {storeUnit_maskInput_hi[1183:1168]},
     {storeUnit_maskInput_hi[1167:1152]},
     {storeUnit_maskInput_hi[1151:1136]},
     {storeUnit_maskInput_hi[1135:1120]},
     {storeUnit_maskInput_hi[1119:1104]},
     {storeUnit_maskInput_hi[1103:1088]},
     {storeUnit_maskInput_hi[1087:1072]},
     {storeUnit_maskInput_hi[1071:1056]},
     {storeUnit_maskInput_hi[1055:1040]},
     {storeUnit_maskInput_hi[1039:1024]},
     {storeUnit_maskInput_hi[1023:1008]},
     {storeUnit_maskInput_hi[1007:992]},
     {storeUnit_maskInput_hi[991:976]},
     {storeUnit_maskInput_hi[975:960]},
     {storeUnit_maskInput_hi[959:944]},
     {storeUnit_maskInput_hi[943:928]},
     {storeUnit_maskInput_hi[927:912]},
     {storeUnit_maskInput_hi[911:896]},
     {storeUnit_maskInput_hi[895:880]},
     {storeUnit_maskInput_hi[879:864]},
     {storeUnit_maskInput_hi[863:848]},
     {storeUnit_maskInput_hi[847:832]},
     {storeUnit_maskInput_hi[831:816]},
     {storeUnit_maskInput_hi[815:800]},
     {storeUnit_maskInput_hi[799:784]},
     {storeUnit_maskInput_hi[783:768]},
     {storeUnit_maskInput_hi[767:752]},
     {storeUnit_maskInput_hi[751:736]},
     {storeUnit_maskInput_hi[735:720]},
     {storeUnit_maskInput_hi[719:704]},
     {storeUnit_maskInput_hi[703:688]},
     {storeUnit_maskInput_hi[687:672]},
     {storeUnit_maskInput_hi[671:656]},
     {storeUnit_maskInput_hi[655:640]},
     {storeUnit_maskInput_hi[639:624]},
     {storeUnit_maskInput_hi[623:608]},
     {storeUnit_maskInput_hi[607:592]},
     {storeUnit_maskInput_hi[591:576]},
     {storeUnit_maskInput_hi[575:560]},
     {storeUnit_maskInput_hi[559:544]},
     {storeUnit_maskInput_hi[543:528]},
     {storeUnit_maskInput_hi[527:512]},
     {storeUnit_maskInput_hi[511:496]},
     {storeUnit_maskInput_hi[495:480]},
     {storeUnit_maskInput_hi[479:464]},
     {storeUnit_maskInput_hi[463:448]},
     {storeUnit_maskInput_hi[447:432]},
     {storeUnit_maskInput_hi[431:416]},
     {storeUnit_maskInput_hi[415:400]},
     {storeUnit_maskInput_hi[399:384]},
     {storeUnit_maskInput_hi[383:368]},
     {storeUnit_maskInput_hi[367:352]},
     {storeUnit_maskInput_hi[351:336]},
     {storeUnit_maskInput_hi[335:320]},
     {storeUnit_maskInput_hi[319:304]},
     {storeUnit_maskInput_hi[303:288]},
     {storeUnit_maskInput_hi[287:272]},
     {storeUnit_maskInput_hi[271:256]},
     {storeUnit_maskInput_hi[255:240]},
     {storeUnit_maskInput_hi[239:224]},
     {storeUnit_maskInput_hi[223:208]},
     {storeUnit_maskInput_hi[207:192]},
     {storeUnit_maskInput_hi[191:176]},
     {storeUnit_maskInput_hi[175:160]},
     {storeUnit_maskInput_hi[159:144]},
     {storeUnit_maskInput_hi[143:128]},
     {storeUnit_maskInput_hi[127:112]},
     {storeUnit_maskInput_hi[111:96]},
     {storeUnit_maskInput_hi[95:80]},
     {storeUnit_maskInput_hi[79:64]},
     {storeUnit_maskInput_hi[63:48]},
     {storeUnit_maskInput_hi[47:32]},
     {storeUnit_maskInput_hi[31:16]},
     {storeUnit_maskInput_hi[15:0]},
     {storeUnit_maskInput_lo[4095:4080]},
     {storeUnit_maskInput_lo[4079:4064]},
     {storeUnit_maskInput_lo[4063:4048]},
     {storeUnit_maskInput_lo[4047:4032]},
     {storeUnit_maskInput_lo[4031:4016]},
     {storeUnit_maskInput_lo[4015:4000]},
     {storeUnit_maskInput_lo[3999:3984]},
     {storeUnit_maskInput_lo[3983:3968]},
     {storeUnit_maskInput_lo[3967:3952]},
     {storeUnit_maskInput_lo[3951:3936]},
     {storeUnit_maskInput_lo[3935:3920]},
     {storeUnit_maskInput_lo[3919:3904]},
     {storeUnit_maskInput_lo[3903:3888]},
     {storeUnit_maskInput_lo[3887:3872]},
     {storeUnit_maskInput_lo[3871:3856]},
     {storeUnit_maskInput_lo[3855:3840]},
     {storeUnit_maskInput_lo[3839:3824]},
     {storeUnit_maskInput_lo[3823:3808]},
     {storeUnit_maskInput_lo[3807:3792]},
     {storeUnit_maskInput_lo[3791:3776]},
     {storeUnit_maskInput_lo[3775:3760]},
     {storeUnit_maskInput_lo[3759:3744]},
     {storeUnit_maskInput_lo[3743:3728]},
     {storeUnit_maskInput_lo[3727:3712]},
     {storeUnit_maskInput_lo[3711:3696]},
     {storeUnit_maskInput_lo[3695:3680]},
     {storeUnit_maskInput_lo[3679:3664]},
     {storeUnit_maskInput_lo[3663:3648]},
     {storeUnit_maskInput_lo[3647:3632]},
     {storeUnit_maskInput_lo[3631:3616]},
     {storeUnit_maskInput_lo[3615:3600]},
     {storeUnit_maskInput_lo[3599:3584]},
     {storeUnit_maskInput_lo[3583:3568]},
     {storeUnit_maskInput_lo[3567:3552]},
     {storeUnit_maskInput_lo[3551:3536]},
     {storeUnit_maskInput_lo[3535:3520]},
     {storeUnit_maskInput_lo[3519:3504]},
     {storeUnit_maskInput_lo[3503:3488]},
     {storeUnit_maskInput_lo[3487:3472]},
     {storeUnit_maskInput_lo[3471:3456]},
     {storeUnit_maskInput_lo[3455:3440]},
     {storeUnit_maskInput_lo[3439:3424]},
     {storeUnit_maskInput_lo[3423:3408]},
     {storeUnit_maskInput_lo[3407:3392]},
     {storeUnit_maskInput_lo[3391:3376]},
     {storeUnit_maskInput_lo[3375:3360]},
     {storeUnit_maskInput_lo[3359:3344]},
     {storeUnit_maskInput_lo[3343:3328]},
     {storeUnit_maskInput_lo[3327:3312]},
     {storeUnit_maskInput_lo[3311:3296]},
     {storeUnit_maskInput_lo[3295:3280]},
     {storeUnit_maskInput_lo[3279:3264]},
     {storeUnit_maskInput_lo[3263:3248]},
     {storeUnit_maskInput_lo[3247:3232]},
     {storeUnit_maskInput_lo[3231:3216]},
     {storeUnit_maskInput_lo[3215:3200]},
     {storeUnit_maskInput_lo[3199:3184]},
     {storeUnit_maskInput_lo[3183:3168]},
     {storeUnit_maskInput_lo[3167:3152]},
     {storeUnit_maskInput_lo[3151:3136]},
     {storeUnit_maskInput_lo[3135:3120]},
     {storeUnit_maskInput_lo[3119:3104]},
     {storeUnit_maskInput_lo[3103:3088]},
     {storeUnit_maskInput_lo[3087:3072]},
     {storeUnit_maskInput_lo[3071:3056]},
     {storeUnit_maskInput_lo[3055:3040]},
     {storeUnit_maskInput_lo[3039:3024]},
     {storeUnit_maskInput_lo[3023:3008]},
     {storeUnit_maskInput_lo[3007:2992]},
     {storeUnit_maskInput_lo[2991:2976]},
     {storeUnit_maskInput_lo[2975:2960]},
     {storeUnit_maskInput_lo[2959:2944]},
     {storeUnit_maskInput_lo[2943:2928]},
     {storeUnit_maskInput_lo[2927:2912]},
     {storeUnit_maskInput_lo[2911:2896]},
     {storeUnit_maskInput_lo[2895:2880]},
     {storeUnit_maskInput_lo[2879:2864]},
     {storeUnit_maskInput_lo[2863:2848]},
     {storeUnit_maskInput_lo[2847:2832]},
     {storeUnit_maskInput_lo[2831:2816]},
     {storeUnit_maskInput_lo[2815:2800]},
     {storeUnit_maskInput_lo[2799:2784]},
     {storeUnit_maskInput_lo[2783:2768]},
     {storeUnit_maskInput_lo[2767:2752]},
     {storeUnit_maskInput_lo[2751:2736]},
     {storeUnit_maskInput_lo[2735:2720]},
     {storeUnit_maskInput_lo[2719:2704]},
     {storeUnit_maskInput_lo[2703:2688]},
     {storeUnit_maskInput_lo[2687:2672]},
     {storeUnit_maskInput_lo[2671:2656]},
     {storeUnit_maskInput_lo[2655:2640]},
     {storeUnit_maskInput_lo[2639:2624]},
     {storeUnit_maskInput_lo[2623:2608]},
     {storeUnit_maskInput_lo[2607:2592]},
     {storeUnit_maskInput_lo[2591:2576]},
     {storeUnit_maskInput_lo[2575:2560]},
     {storeUnit_maskInput_lo[2559:2544]},
     {storeUnit_maskInput_lo[2543:2528]},
     {storeUnit_maskInput_lo[2527:2512]},
     {storeUnit_maskInput_lo[2511:2496]},
     {storeUnit_maskInput_lo[2495:2480]},
     {storeUnit_maskInput_lo[2479:2464]},
     {storeUnit_maskInput_lo[2463:2448]},
     {storeUnit_maskInput_lo[2447:2432]},
     {storeUnit_maskInput_lo[2431:2416]},
     {storeUnit_maskInput_lo[2415:2400]},
     {storeUnit_maskInput_lo[2399:2384]},
     {storeUnit_maskInput_lo[2383:2368]},
     {storeUnit_maskInput_lo[2367:2352]},
     {storeUnit_maskInput_lo[2351:2336]},
     {storeUnit_maskInput_lo[2335:2320]},
     {storeUnit_maskInput_lo[2319:2304]},
     {storeUnit_maskInput_lo[2303:2288]},
     {storeUnit_maskInput_lo[2287:2272]},
     {storeUnit_maskInput_lo[2271:2256]},
     {storeUnit_maskInput_lo[2255:2240]},
     {storeUnit_maskInput_lo[2239:2224]},
     {storeUnit_maskInput_lo[2223:2208]},
     {storeUnit_maskInput_lo[2207:2192]},
     {storeUnit_maskInput_lo[2191:2176]},
     {storeUnit_maskInput_lo[2175:2160]},
     {storeUnit_maskInput_lo[2159:2144]},
     {storeUnit_maskInput_lo[2143:2128]},
     {storeUnit_maskInput_lo[2127:2112]},
     {storeUnit_maskInput_lo[2111:2096]},
     {storeUnit_maskInput_lo[2095:2080]},
     {storeUnit_maskInput_lo[2079:2064]},
     {storeUnit_maskInput_lo[2063:2048]},
     {storeUnit_maskInput_lo[2047:2032]},
     {storeUnit_maskInput_lo[2031:2016]},
     {storeUnit_maskInput_lo[2015:2000]},
     {storeUnit_maskInput_lo[1999:1984]},
     {storeUnit_maskInput_lo[1983:1968]},
     {storeUnit_maskInput_lo[1967:1952]},
     {storeUnit_maskInput_lo[1951:1936]},
     {storeUnit_maskInput_lo[1935:1920]},
     {storeUnit_maskInput_lo[1919:1904]},
     {storeUnit_maskInput_lo[1903:1888]},
     {storeUnit_maskInput_lo[1887:1872]},
     {storeUnit_maskInput_lo[1871:1856]},
     {storeUnit_maskInput_lo[1855:1840]},
     {storeUnit_maskInput_lo[1839:1824]},
     {storeUnit_maskInput_lo[1823:1808]},
     {storeUnit_maskInput_lo[1807:1792]},
     {storeUnit_maskInput_lo[1791:1776]},
     {storeUnit_maskInput_lo[1775:1760]},
     {storeUnit_maskInput_lo[1759:1744]},
     {storeUnit_maskInput_lo[1743:1728]},
     {storeUnit_maskInput_lo[1727:1712]},
     {storeUnit_maskInput_lo[1711:1696]},
     {storeUnit_maskInput_lo[1695:1680]},
     {storeUnit_maskInput_lo[1679:1664]},
     {storeUnit_maskInput_lo[1663:1648]},
     {storeUnit_maskInput_lo[1647:1632]},
     {storeUnit_maskInput_lo[1631:1616]},
     {storeUnit_maskInput_lo[1615:1600]},
     {storeUnit_maskInput_lo[1599:1584]},
     {storeUnit_maskInput_lo[1583:1568]},
     {storeUnit_maskInput_lo[1567:1552]},
     {storeUnit_maskInput_lo[1551:1536]},
     {storeUnit_maskInput_lo[1535:1520]},
     {storeUnit_maskInput_lo[1519:1504]},
     {storeUnit_maskInput_lo[1503:1488]},
     {storeUnit_maskInput_lo[1487:1472]},
     {storeUnit_maskInput_lo[1471:1456]},
     {storeUnit_maskInput_lo[1455:1440]},
     {storeUnit_maskInput_lo[1439:1424]},
     {storeUnit_maskInput_lo[1423:1408]},
     {storeUnit_maskInput_lo[1407:1392]},
     {storeUnit_maskInput_lo[1391:1376]},
     {storeUnit_maskInput_lo[1375:1360]},
     {storeUnit_maskInput_lo[1359:1344]},
     {storeUnit_maskInput_lo[1343:1328]},
     {storeUnit_maskInput_lo[1327:1312]},
     {storeUnit_maskInput_lo[1311:1296]},
     {storeUnit_maskInput_lo[1295:1280]},
     {storeUnit_maskInput_lo[1279:1264]},
     {storeUnit_maskInput_lo[1263:1248]},
     {storeUnit_maskInput_lo[1247:1232]},
     {storeUnit_maskInput_lo[1231:1216]},
     {storeUnit_maskInput_lo[1215:1200]},
     {storeUnit_maskInput_lo[1199:1184]},
     {storeUnit_maskInput_lo[1183:1168]},
     {storeUnit_maskInput_lo[1167:1152]},
     {storeUnit_maskInput_lo[1151:1136]},
     {storeUnit_maskInput_lo[1135:1120]},
     {storeUnit_maskInput_lo[1119:1104]},
     {storeUnit_maskInput_lo[1103:1088]},
     {storeUnit_maskInput_lo[1087:1072]},
     {storeUnit_maskInput_lo[1071:1056]},
     {storeUnit_maskInput_lo[1055:1040]},
     {storeUnit_maskInput_lo[1039:1024]},
     {storeUnit_maskInput_lo[1023:1008]},
     {storeUnit_maskInput_lo[1007:992]},
     {storeUnit_maskInput_lo[991:976]},
     {storeUnit_maskInput_lo[975:960]},
     {storeUnit_maskInput_lo[959:944]},
     {storeUnit_maskInput_lo[943:928]},
     {storeUnit_maskInput_lo[927:912]},
     {storeUnit_maskInput_lo[911:896]},
     {storeUnit_maskInput_lo[895:880]},
     {storeUnit_maskInput_lo[879:864]},
     {storeUnit_maskInput_lo[863:848]},
     {storeUnit_maskInput_lo[847:832]},
     {storeUnit_maskInput_lo[831:816]},
     {storeUnit_maskInput_lo[815:800]},
     {storeUnit_maskInput_lo[799:784]},
     {storeUnit_maskInput_lo[783:768]},
     {storeUnit_maskInput_lo[767:752]},
     {storeUnit_maskInput_lo[751:736]},
     {storeUnit_maskInput_lo[735:720]},
     {storeUnit_maskInput_lo[719:704]},
     {storeUnit_maskInput_lo[703:688]},
     {storeUnit_maskInput_lo[687:672]},
     {storeUnit_maskInput_lo[671:656]},
     {storeUnit_maskInput_lo[655:640]},
     {storeUnit_maskInput_lo[639:624]},
     {storeUnit_maskInput_lo[623:608]},
     {storeUnit_maskInput_lo[607:592]},
     {storeUnit_maskInput_lo[591:576]},
     {storeUnit_maskInput_lo[575:560]},
     {storeUnit_maskInput_lo[559:544]},
     {storeUnit_maskInput_lo[543:528]},
     {storeUnit_maskInput_lo[527:512]},
     {storeUnit_maskInput_lo[511:496]},
     {storeUnit_maskInput_lo[495:480]},
     {storeUnit_maskInput_lo[479:464]},
     {storeUnit_maskInput_lo[463:448]},
     {storeUnit_maskInput_lo[447:432]},
     {storeUnit_maskInput_lo[431:416]},
     {storeUnit_maskInput_lo[415:400]},
     {storeUnit_maskInput_lo[399:384]},
     {storeUnit_maskInput_lo[383:368]},
     {storeUnit_maskInput_lo[367:352]},
     {storeUnit_maskInput_lo[351:336]},
     {storeUnit_maskInput_lo[335:320]},
     {storeUnit_maskInput_lo[319:304]},
     {storeUnit_maskInput_lo[303:288]},
     {storeUnit_maskInput_lo[287:272]},
     {storeUnit_maskInput_lo[271:256]},
     {storeUnit_maskInput_lo[255:240]},
     {storeUnit_maskInput_lo[239:224]},
     {storeUnit_maskInput_lo[223:208]},
     {storeUnit_maskInput_lo[207:192]},
     {storeUnit_maskInput_lo[191:176]},
     {storeUnit_maskInput_lo[175:160]},
     {storeUnit_maskInput_lo[159:144]},
     {storeUnit_maskInput_lo[143:128]},
     {storeUnit_maskInput_lo[127:112]},
     {storeUnit_maskInput_lo[111:96]},
     {storeUnit_maskInput_lo[95:80]},
     {storeUnit_maskInput_lo[79:64]},
     {storeUnit_maskInput_lo[63:48]},
     {storeUnit_maskInput_lo[47:32]},
     {storeUnit_maskInput_lo[31:16]},
     {storeUnit_maskInput_lo[15:0]}};
  wire [8:0]         maskSelect_2 = _otherUnit_maskSelect_valid ? _otherUnit_maskSelect_bits : 9'h0;
  wire [127:0]       otherUnit_maskInput_lo_lo_lo_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_lo_lo_lo_lo_hi = {otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]       otherUnit_maskInput_lo_lo_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_lo_lo_lo_hi_lo = {otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_lo_lo_lo_hi_hi = {otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]       otherUnit_maskInput_lo_lo_lo_lo_hi = {otherUnit_maskInput_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_lo};
  wire [511:0]       otherUnit_maskInput_lo_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_lo_lo_hi_lo_lo = {otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_lo_lo_hi_lo_hi = {otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]       otherUnit_maskInput_lo_lo_lo_hi_lo = {otherUnit_maskInput_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_lo_lo_hi_hi_lo = {otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_lo_lo_hi_hi_hi = {otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]       otherUnit_maskInput_lo_lo_lo_hi_hi = {otherUnit_maskInput_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_lo};
  wire [511:0]       otherUnit_maskInput_lo_lo_lo_hi = {otherUnit_maskInput_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_lo};
  wire [1023:0]      otherUnit_maskInput_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_lo_hi_lo_lo_lo = {otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_lo_hi_lo_lo_hi = {otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]       otherUnit_maskInput_lo_lo_hi_lo_lo = {otherUnit_maskInput_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_lo_hi_lo_hi_lo = {otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_lo_hi_lo_hi_hi = {otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]       otherUnit_maskInput_lo_lo_hi_lo_hi = {otherUnit_maskInput_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_lo};
  wire [511:0]       otherUnit_maskInput_lo_lo_hi_lo = {otherUnit_maskInput_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_lo_hi_hi_lo_lo = {otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_lo_hi_hi_lo_hi = {otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]       otherUnit_maskInput_lo_lo_hi_hi_lo = {otherUnit_maskInput_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_lo_hi_hi_hi_lo = {otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_lo_hi_hi_hi_hi = {otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]       otherUnit_maskInput_lo_lo_hi_hi_hi = {otherUnit_maskInput_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_lo};
  wire [511:0]       otherUnit_maskInput_lo_lo_hi_hi = {otherUnit_maskInput_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_lo};
  wire [1023:0]      otherUnit_maskInput_lo_lo_hi = {otherUnit_maskInput_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo};
  wire [2047:0]      otherUnit_maskInput_lo_lo = {otherUnit_maskInput_lo_lo_hi, otherUnit_maskInput_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_hi_lo_lo_lo_lo = {otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_hi_lo_lo_lo_hi = {otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]       otherUnit_maskInput_lo_hi_lo_lo_lo = {otherUnit_maskInput_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_hi_lo_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_hi_lo_lo_hi_hi = {otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]       otherUnit_maskInput_lo_hi_lo_lo_hi = {otherUnit_maskInput_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_lo};
  wire [511:0]       otherUnit_maskInput_lo_hi_lo_lo = {otherUnit_maskInput_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_hi_lo_hi_lo_lo = {otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_hi_lo_hi_lo_hi = {otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]       otherUnit_maskInput_lo_hi_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_hi_lo_hi_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_hi_lo_hi_hi_hi = {otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]       otherUnit_maskInput_lo_hi_lo_hi_hi = {otherUnit_maskInput_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_lo};
  wire [511:0]       otherUnit_maskInput_lo_hi_lo_hi = {otherUnit_maskInput_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_lo};
  wire [1023:0]      otherUnit_maskInput_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_hi_hi_lo_lo_lo = {otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_hi_hi_lo_lo_hi = {otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]       otherUnit_maskInput_lo_hi_hi_lo_lo = {otherUnit_maskInput_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_hi_hi_lo_hi_lo = {otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_hi_hi_lo_hi_hi = {otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]       otherUnit_maskInput_lo_hi_hi_lo_hi = {otherUnit_maskInput_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_lo};
  wire [511:0]       otherUnit_maskInput_lo_hi_hi_lo = {otherUnit_maskInput_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_hi_hi_hi_lo_lo = {otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_hi_hi_hi_lo_hi = {otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]       otherUnit_maskInput_lo_hi_hi_hi_lo = {otherUnit_maskInput_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_hi_hi_hi_hi_lo = {otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_lo_hi_hi_hi_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]       otherUnit_maskInput_lo_hi_hi_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_lo};
  wire [511:0]       otherUnit_maskInput_lo_hi_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_lo};
  wire [1023:0]      otherUnit_maskInput_lo_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_lo};
  wire [2047:0]      otherUnit_maskInput_lo_hi = {otherUnit_maskInput_lo_hi_hi, otherUnit_maskInput_lo_hi_lo};
  wire [4095:0]      otherUnit_maskInput_lo = {otherUnit_maskInput_lo_hi, otherUnit_maskInput_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_lo_lo_lo_lo_lo = {otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_lo_lo_lo_lo_hi = {otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]       otherUnit_maskInput_hi_lo_lo_lo_lo = {otherUnit_maskInput_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_lo_lo_lo_hi_lo = {otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_lo_lo_lo_hi_hi = {otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]       otherUnit_maskInput_hi_lo_lo_lo_hi = {otherUnit_maskInput_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_lo};
  wire [511:0]       otherUnit_maskInput_hi_lo_lo_lo = {otherUnit_maskInput_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_lo_lo_hi_lo_lo = {otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_lo_lo_hi_lo_hi = {otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]       otherUnit_maskInput_hi_lo_lo_hi_lo = {otherUnit_maskInput_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_lo_lo_hi_hi_lo = {otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_lo_lo_hi_hi_hi = {otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]       otherUnit_maskInput_hi_lo_lo_hi_hi = {otherUnit_maskInput_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_lo};
  wire [511:0]       otherUnit_maskInput_hi_lo_lo_hi = {otherUnit_maskInput_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_lo};
  wire [1023:0]      otherUnit_maskInput_hi_lo_lo = {otherUnit_maskInput_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_lo_hi_lo_lo_lo = {otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_lo_hi_lo_lo_hi = {otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]       otherUnit_maskInput_hi_lo_hi_lo_lo = {otherUnit_maskInput_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_lo_hi_lo_hi_lo = {otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_lo_hi_lo_hi_hi = {otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]       otherUnit_maskInput_hi_lo_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_lo};
  wire [511:0]       otherUnit_maskInput_hi_lo_hi_lo = {otherUnit_maskInput_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_lo_hi_hi_lo_lo = {otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_lo_hi_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]       otherUnit_maskInput_hi_lo_hi_hi_lo = {otherUnit_maskInput_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_lo_hi_hi_hi_lo = {otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_lo_hi_hi_hi_hi = {otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]       otherUnit_maskInput_hi_lo_hi_hi_hi = {otherUnit_maskInput_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_lo};
  wire [511:0]       otherUnit_maskInput_hi_lo_hi_hi = {otherUnit_maskInput_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_lo};
  wire [1023:0]      otherUnit_maskInput_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo};
  wire [2047:0]      otherUnit_maskInput_hi_lo = {otherUnit_maskInput_hi_lo_hi, otherUnit_maskInput_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_hi_lo_lo_lo_lo = {otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_hi_lo_lo_lo_hi = {otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]       otherUnit_maskInput_hi_hi_lo_lo_lo = {otherUnit_maskInput_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_hi_lo_lo_hi_lo = {otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_hi_lo_lo_hi_hi = {otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]       otherUnit_maskInput_hi_hi_lo_lo_hi = {otherUnit_maskInput_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_lo};
  wire [511:0]       otherUnit_maskInput_hi_hi_lo_lo = {otherUnit_maskInput_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_hi_lo_hi_lo_lo = {otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_hi_lo_hi_lo_hi = {otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]       otherUnit_maskInput_hi_hi_lo_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_hi_lo_hi_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_hi_lo_hi_hi_hi = {otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]       otherUnit_maskInput_hi_hi_lo_hi_hi = {otherUnit_maskInput_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_lo};
  wire [511:0]       otherUnit_maskInput_hi_hi_lo_hi = {otherUnit_maskInput_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_lo};
  wire [1023:0]      otherUnit_maskInput_hi_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_hi_hi_lo_lo_lo = {otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_hi_hi_lo_lo_hi = {otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]       otherUnit_maskInput_hi_hi_hi_lo_lo = {otherUnit_maskInput_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_hi_hi_lo_hi_lo = {otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_hi_hi_lo_hi_hi = {otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]       otherUnit_maskInput_hi_hi_hi_lo_hi = {otherUnit_maskInput_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_lo};
  wire [511:0]       otherUnit_maskInput_hi_hi_hi_lo = {otherUnit_maskInput_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_hi_hi_hi_lo_lo = {otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_hi_hi_hi_lo_hi = {otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]       otherUnit_maskInput_hi_hi_hi_hi_lo = {otherUnit_maskInput_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_hi_hi_hi_hi_lo = {otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]       otherUnit_maskInput_hi_hi_hi_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]       otherUnit_maskInput_hi_hi_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_lo};
  wire [511:0]       otherUnit_maskInput_hi_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_lo};
  wire [1023:0]      otherUnit_maskInput_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_lo};
  wire [2047:0]      otherUnit_maskInput_hi_hi = {otherUnit_maskInput_hi_hi_hi, otherUnit_maskInput_hi_hi_lo};
  wire [4095:0]      otherUnit_maskInput_hi = {otherUnit_maskInput_hi_hi, otherUnit_maskInput_hi_lo};
  wire [511:0][15:0] _GEN_129 =
    {{otherUnit_maskInput_hi[4095:4080]},
     {otherUnit_maskInput_hi[4079:4064]},
     {otherUnit_maskInput_hi[4063:4048]},
     {otherUnit_maskInput_hi[4047:4032]},
     {otherUnit_maskInput_hi[4031:4016]},
     {otherUnit_maskInput_hi[4015:4000]},
     {otherUnit_maskInput_hi[3999:3984]},
     {otherUnit_maskInput_hi[3983:3968]},
     {otherUnit_maskInput_hi[3967:3952]},
     {otherUnit_maskInput_hi[3951:3936]},
     {otherUnit_maskInput_hi[3935:3920]},
     {otherUnit_maskInput_hi[3919:3904]},
     {otherUnit_maskInput_hi[3903:3888]},
     {otherUnit_maskInput_hi[3887:3872]},
     {otherUnit_maskInput_hi[3871:3856]},
     {otherUnit_maskInput_hi[3855:3840]},
     {otherUnit_maskInput_hi[3839:3824]},
     {otherUnit_maskInput_hi[3823:3808]},
     {otherUnit_maskInput_hi[3807:3792]},
     {otherUnit_maskInput_hi[3791:3776]},
     {otherUnit_maskInput_hi[3775:3760]},
     {otherUnit_maskInput_hi[3759:3744]},
     {otherUnit_maskInput_hi[3743:3728]},
     {otherUnit_maskInput_hi[3727:3712]},
     {otherUnit_maskInput_hi[3711:3696]},
     {otherUnit_maskInput_hi[3695:3680]},
     {otherUnit_maskInput_hi[3679:3664]},
     {otherUnit_maskInput_hi[3663:3648]},
     {otherUnit_maskInput_hi[3647:3632]},
     {otherUnit_maskInput_hi[3631:3616]},
     {otherUnit_maskInput_hi[3615:3600]},
     {otherUnit_maskInput_hi[3599:3584]},
     {otherUnit_maskInput_hi[3583:3568]},
     {otherUnit_maskInput_hi[3567:3552]},
     {otherUnit_maskInput_hi[3551:3536]},
     {otherUnit_maskInput_hi[3535:3520]},
     {otherUnit_maskInput_hi[3519:3504]},
     {otherUnit_maskInput_hi[3503:3488]},
     {otherUnit_maskInput_hi[3487:3472]},
     {otherUnit_maskInput_hi[3471:3456]},
     {otherUnit_maskInput_hi[3455:3440]},
     {otherUnit_maskInput_hi[3439:3424]},
     {otherUnit_maskInput_hi[3423:3408]},
     {otherUnit_maskInput_hi[3407:3392]},
     {otherUnit_maskInput_hi[3391:3376]},
     {otherUnit_maskInput_hi[3375:3360]},
     {otherUnit_maskInput_hi[3359:3344]},
     {otherUnit_maskInput_hi[3343:3328]},
     {otherUnit_maskInput_hi[3327:3312]},
     {otherUnit_maskInput_hi[3311:3296]},
     {otherUnit_maskInput_hi[3295:3280]},
     {otherUnit_maskInput_hi[3279:3264]},
     {otherUnit_maskInput_hi[3263:3248]},
     {otherUnit_maskInput_hi[3247:3232]},
     {otherUnit_maskInput_hi[3231:3216]},
     {otherUnit_maskInput_hi[3215:3200]},
     {otherUnit_maskInput_hi[3199:3184]},
     {otherUnit_maskInput_hi[3183:3168]},
     {otherUnit_maskInput_hi[3167:3152]},
     {otherUnit_maskInput_hi[3151:3136]},
     {otherUnit_maskInput_hi[3135:3120]},
     {otherUnit_maskInput_hi[3119:3104]},
     {otherUnit_maskInput_hi[3103:3088]},
     {otherUnit_maskInput_hi[3087:3072]},
     {otherUnit_maskInput_hi[3071:3056]},
     {otherUnit_maskInput_hi[3055:3040]},
     {otherUnit_maskInput_hi[3039:3024]},
     {otherUnit_maskInput_hi[3023:3008]},
     {otherUnit_maskInput_hi[3007:2992]},
     {otherUnit_maskInput_hi[2991:2976]},
     {otherUnit_maskInput_hi[2975:2960]},
     {otherUnit_maskInput_hi[2959:2944]},
     {otherUnit_maskInput_hi[2943:2928]},
     {otherUnit_maskInput_hi[2927:2912]},
     {otherUnit_maskInput_hi[2911:2896]},
     {otherUnit_maskInput_hi[2895:2880]},
     {otherUnit_maskInput_hi[2879:2864]},
     {otherUnit_maskInput_hi[2863:2848]},
     {otherUnit_maskInput_hi[2847:2832]},
     {otherUnit_maskInput_hi[2831:2816]},
     {otherUnit_maskInput_hi[2815:2800]},
     {otherUnit_maskInput_hi[2799:2784]},
     {otherUnit_maskInput_hi[2783:2768]},
     {otherUnit_maskInput_hi[2767:2752]},
     {otherUnit_maskInput_hi[2751:2736]},
     {otherUnit_maskInput_hi[2735:2720]},
     {otherUnit_maskInput_hi[2719:2704]},
     {otherUnit_maskInput_hi[2703:2688]},
     {otherUnit_maskInput_hi[2687:2672]},
     {otherUnit_maskInput_hi[2671:2656]},
     {otherUnit_maskInput_hi[2655:2640]},
     {otherUnit_maskInput_hi[2639:2624]},
     {otherUnit_maskInput_hi[2623:2608]},
     {otherUnit_maskInput_hi[2607:2592]},
     {otherUnit_maskInput_hi[2591:2576]},
     {otherUnit_maskInput_hi[2575:2560]},
     {otherUnit_maskInput_hi[2559:2544]},
     {otherUnit_maskInput_hi[2543:2528]},
     {otherUnit_maskInput_hi[2527:2512]},
     {otherUnit_maskInput_hi[2511:2496]},
     {otherUnit_maskInput_hi[2495:2480]},
     {otherUnit_maskInput_hi[2479:2464]},
     {otherUnit_maskInput_hi[2463:2448]},
     {otherUnit_maskInput_hi[2447:2432]},
     {otherUnit_maskInput_hi[2431:2416]},
     {otherUnit_maskInput_hi[2415:2400]},
     {otherUnit_maskInput_hi[2399:2384]},
     {otherUnit_maskInput_hi[2383:2368]},
     {otherUnit_maskInput_hi[2367:2352]},
     {otherUnit_maskInput_hi[2351:2336]},
     {otherUnit_maskInput_hi[2335:2320]},
     {otherUnit_maskInput_hi[2319:2304]},
     {otherUnit_maskInput_hi[2303:2288]},
     {otherUnit_maskInput_hi[2287:2272]},
     {otherUnit_maskInput_hi[2271:2256]},
     {otherUnit_maskInput_hi[2255:2240]},
     {otherUnit_maskInput_hi[2239:2224]},
     {otherUnit_maskInput_hi[2223:2208]},
     {otherUnit_maskInput_hi[2207:2192]},
     {otherUnit_maskInput_hi[2191:2176]},
     {otherUnit_maskInput_hi[2175:2160]},
     {otherUnit_maskInput_hi[2159:2144]},
     {otherUnit_maskInput_hi[2143:2128]},
     {otherUnit_maskInput_hi[2127:2112]},
     {otherUnit_maskInput_hi[2111:2096]},
     {otherUnit_maskInput_hi[2095:2080]},
     {otherUnit_maskInput_hi[2079:2064]},
     {otherUnit_maskInput_hi[2063:2048]},
     {otherUnit_maskInput_hi[2047:2032]},
     {otherUnit_maskInput_hi[2031:2016]},
     {otherUnit_maskInput_hi[2015:2000]},
     {otherUnit_maskInput_hi[1999:1984]},
     {otherUnit_maskInput_hi[1983:1968]},
     {otherUnit_maskInput_hi[1967:1952]},
     {otherUnit_maskInput_hi[1951:1936]},
     {otherUnit_maskInput_hi[1935:1920]},
     {otherUnit_maskInput_hi[1919:1904]},
     {otherUnit_maskInput_hi[1903:1888]},
     {otherUnit_maskInput_hi[1887:1872]},
     {otherUnit_maskInput_hi[1871:1856]},
     {otherUnit_maskInput_hi[1855:1840]},
     {otherUnit_maskInput_hi[1839:1824]},
     {otherUnit_maskInput_hi[1823:1808]},
     {otherUnit_maskInput_hi[1807:1792]},
     {otherUnit_maskInput_hi[1791:1776]},
     {otherUnit_maskInput_hi[1775:1760]},
     {otherUnit_maskInput_hi[1759:1744]},
     {otherUnit_maskInput_hi[1743:1728]},
     {otherUnit_maskInput_hi[1727:1712]},
     {otherUnit_maskInput_hi[1711:1696]},
     {otherUnit_maskInput_hi[1695:1680]},
     {otherUnit_maskInput_hi[1679:1664]},
     {otherUnit_maskInput_hi[1663:1648]},
     {otherUnit_maskInput_hi[1647:1632]},
     {otherUnit_maskInput_hi[1631:1616]},
     {otherUnit_maskInput_hi[1615:1600]},
     {otherUnit_maskInput_hi[1599:1584]},
     {otherUnit_maskInput_hi[1583:1568]},
     {otherUnit_maskInput_hi[1567:1552]},
     {otherUnit_maskInput_hi[1551:1536]},
     {otherUnit_maskInput_hi[1535:1520]},
     {otherUnit_maskInput_hi[1519:1504]},
     {otherUnit_maskInput_hi[1503:1488]},
     {otherUnit_maskInput_hi[1487:1472]},
     {otherUnit_maskInput_hi[1471:1456]},
     {otherUnit_maskInput_hi[1455:1440]},
     {otherUnit_maskInput_hi[1439:1424]},
     {otherUnit_maskInput_hi[1423:1408]},
     {otherUnit_maskInput_hi[1407:1392]},
     {otherUnit_maskInput_hi[1391:1376]},
     {otherUnit_maskInput_hi[1375:1360]},
     {otherUnit_maskInput_hi[1359:1344]},
     {otherUnit_maskInput_hi[1343:1328]},
     {otherUnit_maskInput_hi[1327:1312]},
     {otherUnit_maskInput_hi[1311:1296]},
     {otherUnit_maskInput_hi[1295:1280]},
     {otherUnit_maskInput_hi[1279:1264]},
     {otherUnit_maskInput_hi[1263:1248]},
     {otherUnit_maskInput_hi[1247:1232]},
     {otherUnit_maskInput_hi[1231:1216]},
     {otherUnit_maskInput_hi[1215:1200]},
     {otherUnit_maskInput_hi[1199:1184]},
     {otherUnit_maskInput_hi[1183:1168]},
     {otherUnit_maskInput_hi[1167:1152]},
     {otherUnit_maskInput_hi[1151:1136]},
     {otherUnit_maskInput_hi[1135:1120]},
     {otherUnit_maskInput_hi[1119:1104]},
     {otherUnit_maskInput_hi[1103:1088]},
     {otherUnit_maskInput_hi[1087:1072]},
     {otherUnit_maskInput_hi[1071:1056]},
     {otherUnit_maskInput_hi[1055:1040]},
     {otherUnit_maskInput_hi[1039:1024]},
     {otherUnit_maskInput_hi[1023:1008]},
     {otherUnit_maskInput_hi[1007:992]},
     {otherUnit_maskInput_hi[991:976]},
     {otherUnit_maskInput_hi[975:960]},
     {otherUnit_maskInput_hi[959:944]},
     {otherUnit_maskInput_hi[943:928]},
     {otherUnit_maskInput_hi[927:912]},
     {otherUnit_maskInput_hi[911:896]},
     {otherUnit_maskInput_hi[895:880]},
     {otherUnit_maskInput_hi[879:864]},
     {otherUnit_maskInput_hi[863:848]},
     {otherUnit_maskInput_hi[847:832]},
     {otherUnit_maskInput_hi[831:816]},
     {otherUnit_maskInput_hi[815:800]},
     {otherUnit_maskInput_hi[799:784]},
     {otherUnit_maskInput_hi[783:768]},
     {otherUnit_maskInput_hi[767:752]},
     {otherUnit_maskInput_hi[751:736]},
     {otherUnit_maskInput_hi[735:720]},
     {otherUnit_maskInput_hi[719:704]},
     {otherUnit_maskInput_hi[703:688]},
     {otherUnit_maskInput_hi[687:672]},
     {otherUnit_maskInput_hi[671:656]},
     {otherUnit_maskInput_hi[655:640]},
     {otherUnit_maskInput_hi[639:624]},
     {otherUnit_maskInput_hi[623:608]},
     {otherUnit_maskInput_hi[607:592]},
     {otherUnit_maskInput_hi[591:576]},
     {otherUnit_maskInput_hi[575:560]},
     {otherUnit_maskInput_hi[559:544]},
     {otherUnit_maskInput_hi[543:528]},
     {otherUnit_maskInput_hi[527:512]},
     {otherUnit_maskInput_hi[511:496]},
     {otherUnit_maskInput_hi[495:480]},
     {otherUnit_maskInput_hi[479:464]},
     {otherUnit_maskInput_hi[463:448]},
     {otherUnit_maskInput_hi[447:432]},
     {otherUnit_maskInput_hi[431:416]},
     {otherUnit_maskInput_hi[415:400]},
     {otherUnit_maskInput_hi[399:384]},
     {otherUnit_maskInput_hi[383:368]},
     {otherUnit_maskInput_hi[367:352]},
     {otherUnit_maskInput_hi[351:336]},
     {otherUnit_maskInput_hi[335:320]},
     {otherUnit_maskInput_hi[319:304]},
     {otherUnit_maskInput_hi[303:288]},
     {otherUnit_maskInput_hi[287:272]},
     {otherUnit_maskInput_hi[271:256]},
     {otherUnit_maskInput_hi[255:240]},
     {otherUnit_maskInput_hi[239:224]},
     {otherUnit_maskInput_hi[223:208]},
     {otherUnit_maskInput_hi[207:192]},
     {otherUnit_maskInput_hi[191:176]},
     {otherUnit_maskInput_hi[175:160]},
     {otherUnit_maskInput_hi[159:144]},
     {otherUnit_maskInput_hi[143:128]},
     {otherUnit_maskInput_hi[127:112]},
     {otherUnit_maskInput_hi[111:96]},
     {otherUnit_maskInput_hi[95:80]},
     {otherUnit_maskInput_hi[79:64]},
     {otherUnit_maskInput_hi[63:48]},
     {otherUnit_maskInput_hi[47:32]},
     {otherUnit_maskInput_hi[31:16]},
     {otherUnit_maskInput_hi[15:0]},
     {otherUnit_maskInput_lo[4095:4080]},
     {otherUnit_maskInput_lo[4079:4064]},
     {otherUnit_maskInput_lo[4063:4048]},
     {otherUnit_maskInput_lo[4047:4032]},
     {otherUnit_maskInput_lo[4031:4016]},
     {otherUnit_maskInput_lo[4015:4000]},
     {otherUnit_maskInput_lo[3999:3984]},
     {otherUnit_maskInput_lo[3983:3968]},
     {otherUnit_maskInput_lo[3967:3952]},
     {otherUnit_maskInput_lo[3951:3936]},
     {otherUnit_maskInput_lo[3935:3920]},
     {otherUnit_maskInput_lo[3919:3904]},
     {otherUnit_maskInput_lo[3903:3888]},
     {otherUnit_maskInput_lo[3887:3872]},
     {otherUnit_maskInput_lo[3871:3856]},
     {otherUnit_maskInput_lo[3855:3840]},
     {otherUnit_maskInput_lo[3839:3824]},
     {otherUnit_maskInput_lo[3823:3808]},
     {otherUnit_maskInput_lo[3807:3792]},
     {otherUnit_maskInput_lo[3791:3776]},
     {otherUnit_maskInput_lo[3775:3760]},
     {otherUnit_maskInput_lo[3759:3744]},
     {otherUnit_maskInput_lo[3743:3728]},
     {otherUnit_maskInput_lo[3727:3712]},
     {otherUnit_maskInput_lo[3711:3696]},
     {otherUnit_maskInput_lo[3695:3680]},
     {otherUnit_maskInput_lo[3679:3664]},
     {otherUnit_maskInput_lo[3663:3648]},
     {otherUnit_maskInput_lo[3647:3632]},
     {otherUnit_maskInput_lo[3631:3616]},
     {otherUnit_maskInput_lo[3615:3600]},
     {otherUnit_maskInput_lo[3599:3584]},
     {otherUnit_maskInput_lo[3583:3568]},
     {otherUnit_maskInput_lo[3567:3552]},
     {otherUnit_maskInput_lo[3551:3536]},
     {otherUnit_maskInput_lo[3535:3520]},
     {otherUnit_maskInput_lo[3519:3504]},
     {otherUnit_maskInput_lo[3503:3488]},
     {otherUnit_maskInput_lo[3487:3472]},
     {otherUnit_maskInput_lo[3471:3456]},
     {otherUnit_maskInput_lo[3455:3440]},
     {otherUnit_maskInput_lo[3439:3424]},
     {otherUnit_maskInput_lo[3423:3408]},
     {otherUnit_maskInput_lo[3407:3392]},
     {otherUnit_maskInput_lo[3391:3376]},
     {otherUnit_maskInput_lo[3375:3360]},
     {otherUnit_maskInput_lo[3359:3344]},
     {otherUnit_maskInput_lo[3343:3328]},
     {otherUnit_maskInput_lo[3327:3312]},
     {otherUnit_maskInput_lo[3311:3296]},
     {otherUnit_maskInput_lo[3295:3280]},
     {otherUnit_maskInput_lo[3279:3264]},
     {otherUnit_maskInput_lo[3263:3248]},
     {otherUnit_maskInput_lo[3247:3232]},
     {otherUnit_maskInput_lo[3231:3216]},
     {otherUnit_maskInput_lo[3215:3200]},
     {otherUnit_maskInput_lo[3199:3184]},
     {otherUnit_maskInput_lo[3183:3168]},
     {otherUnit_maskInput_lo[3167:3152]},
     {otherUnit_maskInput_lo[3151:3136]},
     {otherUnit_maskInput_lo[3135:3120]},
     {otherUnit_maskInput_lo[3119:3104]},
     {otherUnit_maskInput_lo[3103:3088]},
     {otherUnit_maskInput_lo[3087:3072]},
     {otherUnit_maskInput_lo[3071:3056]},
     {otherUnit_maskInput_lo[3055:3040]},
     {otherUnit_maskInput_lo[3039:3024]},
     {otherUnit_maskInput_lo[3023:3008]},
     {otherUnit_maskInput_lo[3007:2992]},
     {otherUnit_maskInput_lo[2991:2976]},
     {otherUnit_maskInput_lo[2975:2960]},
     {otherUnit_maskInput_lo[2959:2944]},
     {otherUnit_maskInput_lo[2943:2928]},
     {otherUnit_maskInput_lo[2927:2912]},
     {otherUnit_maskInput_lo[2911:2896]},
     {otherUnit_maskInput_lo[2895:2880]},
     {otherUnit_maskInput_lo[2879:2864]},
     {otherUnit_maskInput_lo[2863:2848]},
     {otherUnit_maskInput_lo[2847:2832]},
     {otherUnit_maskInput_lo[2831:2816]},
     {otherUnit_maskInput_lo[2815:2800]},
     {otherUnit_maskInput_lo[2799:2784]},
     {otherUnit_maskInput_lo[2783:2768]},
     {otherUnit_maskInput_lo[2767:2752]},
     {otherUnit_maskInput_lo[2751:2736]},
     {otherUnit_maskInput_lo[2735:2720]},
     {otherUnit_maskInput_lo[2719:2704]},
     {otherUnit_maskInput_lo[2703:2688]},
     {otherUnit_maskInput_lo[2687:2672]},
     {otherUnit_maskInput_lo[2671:2656]},
     {otherUnit_maskInput_lo[2655:2640]},
     {otherUnit_maskInput_lo[2639:2624]},
     {otherUnit_maskInput_lo[2623:2608]},
     {otherUnit_maskInput_lo[2607:2592]},
     {otherUnit_maskInput_lo[2591:2576]},
     {otherUnit_maskInput_lo[2575:2560]},
     {otherUnit_maskInput_lo[2559:2544]},
     {otherUnit_maskInput_lo[2543:2528]},
     {otherUnit_maskInput_lo[2527:2512]},
     {otherUnit_maskInput_lo[2511:2496]},
     {otherUnit_maskInput_lo[2495:2480]},
     {otherUnit_maskInput_lo[2479:2464]},
     {otherUnit_maskInput_lo[2463:2448]},
     {otherUnit_maskInput_lo[2447:2432]},
     {otherUnit_maskInput_lo[2431:2416]},
     {otherUnit_maskInput_lo[2415:2400]},
     {otherUnit_maskInput_lo[2399:2384]},
     {otherUnit_maskInput_lo[2383:2368]},
     {otherUnit_maskInput_lo[2367:2352]},
     {otherUnit_maskInput_lo[2351:2336]},
     {otherUnit_maskInput_lo[2335:2320]},
     {otherUnit_maskInput_lo[2319:2304]},
     {otherUnit_maskInput_lo[2303:2288]},
     {otherUnit_maskInput_lo[2287:2272]},
     {otherUnit_maskInput_lo[2271:2256]},
     {otherUnit_maskInput_lo[2255:2240]},
     {otherUnit_maskInput_lo[2239:2224]},
     {otherUnit_maskInput_lo[2223:2208]},
     {otherUnit_maskInput_lo[2207:2192]},
     {otherUnit_maskInput_lo[2191:2176]},
     {otherUnit_maskInput_lo[2175:2160]},
     {otherUnit_maskInput_lo[2159:2144]},
     {otherUnit_maskInput_lo[2143:2128]},
     {otherUnit_maskInput_lo[2127:2112]},
     {otherUnit_maskInput_lo[2111:2096]},
     {otherUnit_maskInput_lo[2095:2080]},
     {otherUnit_maskInput_lo[2079:2064]},
     {otherUnit_maskInput_lo[2063:2048]},
     {otherUnit_maskInput_lo[2047:2032]},
     {otherUnit_maskInput_lo[2031:2016]},
     {otherUnit_maskInput_lo[2015:2000]},
     {otherUnit_maskInput_lo[1999:1984]},
     {otherUnit_maskInput_lo[1983:1968]},
     {otherUnit_maskInput_lo[1967:1952]},
     {otherUnit_maskInput_lo[1951:1936]},
     {otherUnit_maskInput_lo[1935:1920]},
     {otherUnit_maskInput_lo[1919:1904]},
     {otherUnit_maskInput_lo[1903:1888]},
     {otherUnit_maskInput_lo[1887:1872]},
     {otherUnit_maskInput_lo[1871:1856]},
     {otherUnit_maskInput_lo[1855:1840]},
     {otherUnit_maskInput_lo[1839:1824]},
     {otherUnit_maskInput_lo[1823:1808]},
     {otherUnit_maskInput_lo[1807:1792]},
     {otherUnit_maskInput_lo[1791:1776]},
     {otherUnit_maskInput_lo[1775:1760]},
     {otherUnit_maskInput_lo[1759:1744]},
     {otherUnit_maskInput_lo[1743:1728]},
     {otherUnit_maskInput_lo[1727:1712]},
     {otherUnit_maskInput_lo[1711:1696]},
     {otherUnit_maskInput_lo[1695:1680]},
     {otherUnit_maskInput_lo[1679:1664]},
     {otherUnit_maskInput_lo[1663:1648]},
     {otherUnit_maskInput_lo[1647:1632]},
     {otherUnit_maskInput_lo[1631:1616]},
     {otherUnit_maskInput_lo[1615:1600]},
     {otherUnit_maskInput_lo[1599:1584]},
     {otherUnit_maskInput_lo[1583:1568]},
     {otherUnit_maskInput_lo[1567:1552]},
     {otherUnit_maskInput_lo[1551:1536]},
     {otherUnit_maskInput_lo[1535:1520]},
     {otherUnit_maskInput_lo[1519:1504]},
     {otherUnit_maskInput_lo[1503:1488]},
     {otherUnit_maskInput_lo[1487:1472]},
     {otherUnit_maskInput_lo[1471:1456]},
     {otherUnit_maskInput_lo[1455:1440]},
     {otherUnit_maskInput_lo[1439:1424]},
     {otherUnit_maskInput_lo[1423:1408]},
     {otherUnit_maskInput_lo[1407:1392]},
     {otherUnit_maskInput_lo[1391:1376]},
     {otherUnit_maskInput_lo[1375:1360]},
     {otherUnit_maskInput_lo[1359:1344]},
     {otherUnit_maskInput_lo[1343:1328]},
     {otherUnit_maskInput_lo[1327:1312]},
     {otherUnit_maskInput_lo[1311:1296]},
     {otherUnit_maskInput_lo[1295:1280]},
     {otherUnit_maskInput_lo[1279:1264]},
     {otherUnit_maskInput_lo[1263:1248]},
     {otherUnit_maskInput_lo[1247:1232]},
     {otherUnit_maskInput_lo[1231:1216]},
     {otherUnit_maskInput_lo[1215:1200]},
     {otherUnit_maskInput_lo[1199:1184]},
     {otherUnit_maskInput_lo[1183:1168]},
     {otherUnit_maskInput_lo[1167:1152]},
     {otherUnit_maskInput_lo[1151:1136]},
     {otherUnit_maskInput_lo[1135:1120]},
     {otherUnit_maskInput_lo[1119:1104]},
     {otherUnit_maskInput_lo[1103:1088]},
     {otherUnit_maskInput_lo[1087:1072]},
     {otherUnit_maskInput_lo[1071:1056]},
     {otherUnit_maskInput_lo[1055:1040]},
     {otherUnit_maskInput_lo[1039:1024]},
     {otherUnit_maskInput_lo[1023:1008]},
     {otherUnit_maskInput_lo[1007:992]},
     {otherUnit_maskInput_lo[991:976]},
     {otherUnit_maskInput_lo[975:960]},
     {otherUnit_maskInput_lo[959:944]},
     {otherUnit_maskInput_lo[943:928]},
     {otherUnit_maskInput_lo[927:912]},
     {otherUnit_maskInput_lo[911:896]},
     {otherUnit_maskInput_lo[895:880]},
     {otherUnit_maskInput_lo[879:864]},
     {otherUnit_maskInput_lo[863:848]},
     {otherUnit_maskInput_lo[847:832]},
     {otherUnit_maskInput_lo[831:816]},
     {otherUnit_maskInput_lo[815:800]},
     {otherUnit_maskInput_lo[799:784]},
     {otherUnit_maskInput_lo[783:768]},
     {otherUnit_maskInput_lo[767:752]},
     {otherUnit_maskInput_lo[751:736]},
     {otherUnit_maskInput_lo[735:720]},
     {otherUnit_maskInput_lo[719:704]},
     {otherUnit_maskInput_lo[703:688]},
     {otherUnit_maskInput_lo[687:672]},
     {otherUnit_maskInput_lo[671:656]},
     {otherUnit_maskInput_lo[655:640]},
     {otherUnit_maskInput_lo[639:624]},
     {otherUnit_maskInput_lo[623:608]},
     {otherUnit_maskInput_lo[607:592]},
     {otherUnit_maskInput_lo[591:576]},
     {otherUnit_maskInput_lo[575:560]},
     {otherUnit_maskInput_lo[559:544]},
     {otherUnit_maskInput_lo[543:528]},
     {otherUnit_maskInput_lo[527:512]},
     {otherUnit_maskInput_lo[511:496]},
     {otherUnit_maskInput_lo[495:480]},
     {otherUnit_maskInput_lo[479:464]},
     {otherUnit_maskInput_lo[463:448]},
     {otherUnit_maskInput_lo[447:432]},
     {otherUnit_maskInput_lo[431:416]},
     {otherUnit_maskInput_lo[415:400]},
     {otherUnit_maskInput_lo[399:384]},
     {otherUnit_maskInput_lo[383:368]},
     {otherUnit_maskInput_lo[367:352]},
     {otherUnit_maskInput_lo[351:336]},
     {otherUnit_maskInput_lo[335:320]},
     {otherUnit_maskInput_lo[319:304]},
     {otherUnit_maskInput_lo[303:288]},
     {otherUnit_maskInput_lo[287:272]},
     {otherUnit_maskInput_lo[271:256]},
     {otherUnit_maskInput_lo[255:240]},
     {otherUnit_maskInput_lo[239:224]},
     {otherUnit_maskInput_lo[223:208]},
     {otherUnit_maskInput_lo[207:192]},
     {otherUnit_maskInput_lo[191:176]},
     {otherUnit_maskInput_lo[175:160]},
     {otherUnit_maskInput_lo[159:144]},
     {otherUnit_maskInput_lo[143:128]},
     {otherUnit_maskInput_lo[127:112]},
     {otherUnit_maskInput_lo[111:96]},
     {otherUnit_maskInput_lo[95:80]},
     {otherUnit_maskInput_lo[79:64]},
     {otherUnit_maskInput_lo[63:48]},
     {otherUnit_maskInput_lo[47:32]},
     {otherUnit_maskInput_lo[31:16]},
     {otherUnit_maskInput_lo[15:0]}};
  wire               vrfWritePort_0_valid_0 = writeQueueVec_0_deq_valid;
  wire [4:0]         vrfWritePort_0_bits_vd_0 = writeQueueVec_0_deq_bits_data_vd;
  wire [5:0]         vrfWritePort_0_bits_offset_0 = writeQueueVec_0_deq_bits_data_offset;
  wire [3:0]         vrfWritePort_0_bits_mask_0 = writeQueueVec_0_deq_bits_data_mask;
  wire [31:0]        vrfWritePort_0_bits_data_0 = writeQueueVec_0_deq_bits_data_data;
  wire               vrfWritePort_0_bits_last_0 = writeQueueVec_0_deq_bits_data_last;
  wire [2:0]         vrfWritePort_0_bits_instructionIndex_0 = writeQueueVec_0_deq_bits_data_instructionIndex;
  wire [2:0]         writeIndexQueue_enq_bits = writeQueueVec_0_deq_bits_data_instructionIndex;
  wire [31:0]        writeQueueVec_0_enq_bits_data_data;
  wire               writeQueueVec_0_enq_bits_data_last;
  wire [32:0]        writeQueueVec_dataIn_lo_hi = {writeQueueVec_0_enq_bits_data_data, writeQueueVec_0_enq_bits_data_last};
  wire [2:0]         writeQueueVec_0_enq_bits_data_instructionIndex;
  wire [35:0]        writeQueueVec_dataIn_lo = {writeQueueVec_dataIn_lo_hi, writeQueueVec_0_enq_bits_data_instructionIndex};
  wire [4:0]         writeQueueVec_0_enq_bits_data_vd;
  wire [5:0]         writeQueueVec_0_enq_bits_data_offset;
  wire [10:0]        writeQueueVec_dataIn_hi_hi = {writeQueueVec_0_enq_bits_data_vd, writeQueueVec_0_enq_bits_data_offset};
  wire [3:0]         writeQueueVec_0_enq_bits_data_mask;
  wire [14:0]        writeQueueVec_dataIn_hi = {writeQueueVec_dataIn_hi_hi, writeQueueVec_0_enq_bits_data_mask};
  wire [54:0]        writeQueueVec_dataIn = {writeQueueVec_dataIn_hi, writeQueueVec_dataIn_lo, 4'h1};
  wire [3:0]         writeQueueVec_dataOut_targetLane = _writeQueueVec_fifo_data_out[3:0];
  wire [2:0]         writeQueueVec_dataOut_data_instructionIndex = _writeQueueVec_fifo_data_out[6:4];
  wire               writeQueueVec_dataOut_data_last = _writeQueueVec_fifo_data_out[7];
  wire [31:0]        writeQueueVec_dataOut_data_data = _writeQueueVec_fifo_data_out[39:8];
  wire [3:0]         writeQueueVec_dataOut_data_mask = _writeQueueVec_fifo_data_out[43:40];
  wire [5:0]         writeQueueVec_dataOut_data_offset = _writeQueueVec_fifo_data_out[49:44];
  wire [4:0]         writeQueueVec_dataOut_data_vd = _writeQueueVec_fifo_data_out[54:50];
  wire               writeQueueVec_0_enq_ready = ~_writeQueueVec_fifo_full;
  wire               writeQueueVec_0_enq_valid;
  wire               _probeWire_slots_0_writeValid_T = writeQueueVec_0_enq_ready & writeQueueVec_0_enq_valid;
  assign writeQueueVec_0_deq_valid = ~_writeQueueVec_fifo_empty | writeQueueVec_0_enq_valid;
  assign writeQueueVec_0_deq_bits_data_vd = _writeQueueVec_fifo_empty ? writeQueueVec_0_enq_bits_data_vd : writeQueueVec_dataOut_data_vd;
  assign writeQueueVec_0_deq_bits_data_offset = _writeQueueVec_fifo_empty ? writeQueueVec_0_enq_bits_data_offset : writeQueueVec_dataOut_data_offset;
  assign writeQueueVec_0_deq_bits_data_mask = _writeQueueVec_fifo_empty ? writeQueueVec_0_enq_bits_data_mask : writeQueueVec_dataOut_data_mask;
  assign writeQueueVec_0_deq_bits_data_data = _writeQueueVec_fifo_empty ? writeQueueVec_0_enq_bits_data_data : writeQueueVec_dataOut_data_data;
  assign writeQueueVec_0_deq_bits_data_last = _writeQueueVec_fifo_empty ? writeQueueVec_0_enq_bits_data_last : writeQueueVec_dataOut_data_last;
  assign writeQueueVec_0_deq_bits_data_instructionIndex = _writeQueueVec_fifo_empty ? writeQueueVec_0_enq_bits_data_instructionIndex : writeQueueVec_dataOut_data_instructionIndex;
  wire [3:0]         writeQueueVec_0_deq_bits_targetLane = _writeQueueVec_fifo_empty ? 4'h1 : writeQueueVec_dataOut_targetLane;
  wire               vrfWritePort_1_valid_0 = writeQueueVec_1_deq_valid;
  wire [4:0]         vrfWritePort_1_bits_vd_0 = writeQueueVec_1_deq_bits_data_vd;
  wire [5:0]         vrfWritePort_1_bits_offset_0 = writeQueueVec_1_deq_bits_data_offset;
  wire [3:0]         vrfWritePort_1_bits_mask_0 = writeQueueVec_1_deq_bits_data_mask;
  wire [31:0]        vrfWritePort_1_bits_data_0 = writeQueueVec_1_deq_bits_data_data;
  wire               vrfWritePort_1_bits_last_0 = writeQueueVec_1_deq_bits_data_last;
  wire [2:0]         vrfWritePort_1_bits_instructionIndex_0 = writeQueueVec_1_deq_bits_data_instructionIndex;
  wire [2:0]         writeIndexQueue_1_enq_bits = writeQueueVec_1_deq_bits_data_instructionIndex;
  wire [31:0]        writeQueueVec_1_enq_bits_data_data;
  wire               writeQueueVec_1_enq_bits_data_last;
  wire [32:0]        writeQueueVec_dataIn_lo_hi_1 = {writeQueueVec_1_enq_bits_data_data, writeQueueVec_1_enq_bits_data_last};
  wire [2:0]         writeQueueVec_1_enq_bits_data_instructionIndex;
  wire [35:0]        writeQueueVec_dataIn_lo_1 = {writeQueueVec_dataIn_lo_hi_1, writeQueueVec_1_enq_bits_data_instructionIndex};
  wire [4:0]         writeQueueVec_1_enq_bits_data_vd;
  wire [5:0]         writeQueueVec_1_enq_bits_data_offset;
  wire [10:0]        writeQueueVec_dataIn_hi_hi_1 = {writeQueueVec_1_enq_bits_data_vd, writeQueueVec_1_enq_bits_data_offset};
  wire [3:0]         writeQueueVec_1_enq_bits_data_mask;
  wire [14:0]        writeQueueVec_dataIn_hi_1 = {writeQueueVec_dataIn_hi_hi_1, writeQueueVec_1_enq_bits_data_mask};
  wire [54:0]        writeQueueVec_dataIn_1 = {writeQueueVec_dataIn_hi_1, writeQueueVec_dataIn_lo_1, 4'h2};
  wire [3:0]         writeQueueVec_dataOut_1_targetLane = _writeQueueVec_fifo_1_data_out[3:0];
  wire [2:0]         writeQueueVec_dataOut_1_data_instructionIndex = _writeQueueVec_fifo_1_data_out[6:4];
  wire               writeQueueVec_dataOut_1_data_last = _writeQueueVec_fifo_1_data_out[7];
  wire [31:0]        writeQueueVec_dataOut_1_data_data = _writeQueueVec_fifo_1_data_out[39:8];
  wire [3:0]         writeQueueVec_dataOut_1_data_mask = _writeQueueVec_fifo_1_data_out[43:40];
  wire [5:0]         writeQueueVec_dataOut_1_data_offset = _writeQueueVec_fifo_1_data_out[49:44];
  wire [4:0]         writeQueueVec_dataOut_1_data_vd = _writeQueueVec_fifo_1_data_out[54:50];
  wire               writeQueueVec_1_enq_ready = ~_writeQueueVec_fifo_1_full;
  wire               writeQueueVec_1_enq_valid;
  wire               _probeWire_slots_1_writeValid_T = writeQueueVec_1_enq_ready & writeQueueVec_1_enq_valid;
  assign writeQueueVec_1_deq_valid = ~_writeQueueVec_fifo_1_empty | writeQueueVec_1_enq_valid;
  assign writeQueueVec_1_deq_bits_data_vd = _writeQueueVec_fifo_1_empty ? writeQueueVec_1_enq_bits_data_vd : writeQueueVec_dataOut_1_data_vd;
  assign writeQueueVec_1_deq_bits_data_offset = _writeQueueVec_fifo_1_empty ? writeQueueVec_1_enq_bits_data_offset : writeQueueVec_dataOut_1_data_offset;
  assign writeQueueVec_1_deq_bits_data_mask = _writeQueueVec_fifo_1_empty ? writeQueueVec_1_enq_bits_data_mask : writeQueueVec_dataOut_1_data_mask;
  assign writeQueueVec_1_deq_bits_data_data = _writeQueueVec_fifo_1_empty ? writeQueueVec_1_enq_bits_data_data : writeQueueVec_dataOut_1_data_data;
  assign writeQueueVec_1_deq_bits_data_last = _writeQueueVec_fifo_1_empty ? writeQueueVec_1_enq_bits_data_last : writeQueueVec_dataOut_1_data_last;
  assign writeQueueVec_1_deq_bits_data_instructionIndex = _writeQueueVec_fifo_1_empty ? writeQueueVec_1_enq_bits_data_instructionIndex : writeQueueVec_dataOut_1_data_instructionIndex;
  wire [3:0]         writeQueueVec_1_deq_bits_targetLane = _writeQueueVec_fifo_1_empty ? 4'h2 : writeQueueVec_dataOut_1_targetLane;
  wire               vrfWritePort_2_valid_0 = writeQueueVec_2_deq_valid;
  wire [4:0]         vrfWritePort_2_bits_vd_0 = writeQueueVec_2_deq_bits_data_vd;
  wire [5:0]         vrfWritePort_2_bits_offset_0 = writeQueueVec_2_deq_bits_data_offset;
  wire [3:0]         vrfWritePort_2_bits_mask_0 = writeQueueVec_2_deq_bits_data_mask;
  wire [31:0]        vrfWritePort_2_bits_data_0 = writeQueueVec_2_deq_bits_data_data;
  wire               vrfWritePort_2_bits_last_0 = writeQueueVec_2_deq_bits_data_last;
  wire [2:0]         vrfWritePort_2_bits_instructionIndex_0 = writeQueueVec_2_deq_bits_data_instructionIndex;
  wire [2:0]         writeIndexQueue_2_enq_bits = writeQueueVec_2_deq_bits_data_instructionIndex;
  wire [31:0]        writeQueueVec_2_enq_bits_data_data;
  wire               writeQueueVec_2_enq_bits_data_last;
  wire [32:0]        writeQueueVec_dataIn_lo_hi_2 = {writeQueueVec_2_enq_bits_data_data, writeQueueVec_2_enq_bits_data_last};
  wire [2:0]         writeQueueVec_2_enq_bits_data_instructionIndex;
  wire [35:0]        writeQueueVec_dataIn_lo_2 = {writeQueueVec_dataIn_lo_hi_2, writeQueueVec_2_enq_bits_data_instructionIndex};
  wire [4:0]         writeQueueVec_2_enq_bits_data_vd;
  wire [5:0]         writeQueueVec_2_enq_bits_data_offset;
  wire [10:0]        writeQueueVec_dataIn_hi_hi_2 = {writeQueueVec_2_enq_bits_data_vd, writeQueueVec_2_enq_bits_data_offset};
  wire [3:0]         writeQueueVec_2_enq_bits_data_mask;
  wire [14:0]        writeQueueVec_dataIn_hi_2 = {writeQueueVec_dataIn_hi_hi_2, writeQueueVec_2_enq_bits_data_mask};
  wire [54:0]        writeQueueVec_dataIn_2 = {writeQueueVec_dataIn_hi_2, writeQueueVec_dataIn_lo_2, 4'h4};
  wire [3:0]         writeQueueVec_dataOut_2_targetLane = _writeQueueVec_fifo_2_data_out[3:0];
  wire [2:0]         writeQueueVec_dataOut_2_data_instructionIndex = _writeQueueVec_fifo_2_data_out[6:4];
  wire               writeQueueVec_dataOut_2_data_last = _writeQueueVec_fifo_2_data_out[7];
  wire [31:0]        writeQueueVec_dataOut_2_data_data = _writeQueueVec_fifo_2_data_out[39:8];
  wire [3:0]         writeQueueVec_dataOut_2_data_mask = _writeQueueVec_fifo_2_data_out[43:40];
  wire [5:0]         writeQueueVec_dataOut_2_data_offset = _writeQueueVec_fifo_2_data_out[49:44];
  wire [4:0]         writeQueueVec_dataOut_2_data_vd = _writeQueueVec_fifo_2_data_out[54:50];
  wire               writeQueueVec_2_enq_ready = ~_writeQueueVec_fifo_2_full;
  wire               writeQueueVec_2_enq_valid;
  wire               _probeWire_slots_2_writeValid_T = writeQueueVec_2_enq_ready & writeQueueVec_2_enq_valid;
  assign writeQueueVec_2_deq_valid = ~_writeQueueVec_fifo_2_empty | writeQueueVec_2_enq_valid;
  assign writeQueueVec_2_deq_bits_data_vd = _writeQueueVec_fifo_2_empty ? writeQueueVec_2_enq_bits_data_vd : writeQueueVec_dataOut_2_data_vd;
  assign writeQueueVec_2_deq_bits_data_offset = _writeQueueVec_fifo_2_empty ? writeQueueVec_2_enq_bits_data_offset : writeQueueVec_dataOut_2_data_offset;
  assign writeQueueVec_2_deq_bits_data_mask = _writeQueueVec_fifo_2_empty ? writeQueueVec_2_enq_bits_data_mask : writeQueueVec_dataOut_2_data_mask;
  assign writeQueueVec_2_deq_bits_data_data = _writeQueueVec_fifo_2_empty ? writeQueueVec_2_enq_bits_data_data : writeQueueVec_dataOut_2_data_data;
  assign writeQueueVec_2_deq_bits_data_last = _writeQueueVec_fifo_2_empty ? writeQueueVec_2_enq_bits_data_last : writeQueueVec_dataOut_2_data_last;
  assign writeQueueVec_2_deq_bits_data_instructionIndex = _writeQueueVec_fifo_2_empty ? writeQueueVec_2_enq_bits_data_instructionIndex : writeQueueVec_dataOut_2_data_instructionIndex;
  wire [3:0]         writeQueueVec_2_deq_bits_targetLane = _writeQueueVec_fifo_2_empty ? 4'h4 : writeQueueVec_dataOut_2_targetLane;
  wire               vrfWritePort_3_valid_0 = writeQueueVec_3_deq_valid;
  wire [4:0]         vrfWritePort_3_bits_vd_0 = writeQueueVec_3_deq_bits_data_vd;
  wire [5:0]         vrfWritePort_3_bits_offset_0 = writeQueueVec_3_deq_bits_data_offset;
  wire [3:0]         vrfWritePort_3_bits_mask_0 = writeQueueVec_3_deq_bits_data_mask;
  wire [31:0]        vrfWritePort_3_bits_data_0 = writeQueueVec_3_deq_bits_data_data;
  wire               vrfWritePort_3_bits_last_0 = writeQueueVec_3_deq_bits_data_last;
  wire [2:0]         vrfWritePort_3_bits_instructionIndex_0 = writeQueueVec_3_deq_bits_data_instructionIndex;
  wire [2:0]         writeIndexQueue_3_enq_bits = writeQueueVec_3_deq_bits_data_instructionIndex;
  wire [31:0]        writeQueueVec_3_enq_bits_data_data;
  wire               writeQueueVec_3_enq_bits_data_last;
  wire [32:0]        writeQueueVec_dataIn_lo_hi_3 = {writeQueueVec_3_enq_bits_data_data, writeQueueVec_3_enq_bits_data_last};
  wire [2:0]         writeQueueVec_3_enq_bits_data_instructionIndex;
  wire [35:0]        writeQueueVec_dataIn_lo_3 = {writeQueueVec_dataIn_lo_hi_3, writeQueueVec_3_enq_bits_data_instructionIndex};
  wire [4:0]         writeQueueVec_3_enq_bits_data_vd;
  wire [5:0]         writeQueueVec_3_enq_bits_data_offset;
  wire [10:0]        writeQueueVec_dataIn_hi_hi_3 = {writeQueueVec_3_enq_bits_data_vd, writeQueueVec_3_enq_bits_data_offset};
  wire [3:0]         writeQueueVec_3_enq_bits_data_mask;
  wire [14:0]        writeQueueVec_dataIn_hi_3 = {writeQueueVec_dataIn_hi_hi_3, writeQueueVec_3_enq_bits_data_mask};
  wire [54:0]        writeQueueVec_dataIn_3 = {writeQueueVec_dataIn_hi_3, writeQueueVec_dataIn_lo_3, 4'h8};
  wire [3:0]         writeQueueVec_dataOut_3_targetLane = _writeQueueVec_fifo_3_data_out[3:0];
  wire [2:0]         writeQueueVec_dataOut_3_data_instructionIndex = _writeQueueVec_fifo_3_data_out[6:4];
  wire               writeQueueVec_dataOut_3_data_last = _writeQueueVec_fifo_3_data_out[7];
  wire [31:0]        writeQueueVec_dataOut_3_data_data = _writeQueueVec_fifo_3_data_out[39:8];
  wire [3:0]         writeQueueVec_dataOut_3_data_mask = _writeQueueVec_fifo_3_data_out[43:40];
  wire [5:0]         writeQueueVec_dataOut_3_data_offset = _writeQueueVec_fifo_3_data_out[49:44];
  wire [4:0]         writeQueueVec_dataOut_3_data_vd = _writeQueueVec_fifo_3_data_out[54:50];
  wire               writeQueueVec_3_enq_ready = ~_writeQueueVec_fifo_3_full;
  wire               writeQueueVec_3_enq_valid;
  wire               _probeWire_slots_3_writeValid_T = writeQueueVec_3_enq_ready & writeQueueVec_3_enq_valid;
  assign writeQueueVec_3_deq_valid = ~_writeQueueVec_fifo_3_empty | writeQueueVec_3_enq_valid;
  assign writeQueueVec_3_deq_bits_data_vd = _writeQueueVec_fifo_3_empty ? writeQueueVec_3_enq_bits_data_vd : writeQueueVec_dataOut_3_data_vd;
  assign writeQueueVec_3_deq_bits_data_offset = _writeQueueVec_fifo_3_empty ? writeQueueVec_3_enq_bits_data_offset : writeQueueVec_dataOut_3_data_offset;
  assign writeQueueVec_3_deq_bits_data_mask = _writeQueueVec_fifo_3_empty ? writeQueueVec_3_enq_bits_data_mask : writeQueueVec_dataOut_3_data_mask;
  assign writeQueueVec_3_deq_bits_data_data = _writeQueueVec_fifo_3_empty ? writeQueueVec_3_enq_bits_data_data : writeQueueVec_dataOut_3_data_data;
  assign writeQueueVec_3_deq_bits_data_last = _writeQueueVec_fifo_3_empty ? writeQueueVec_3_enq_bits_data_last : writeQueueVec_dataOut_3_data_last;
  assign writeQueueVec_3_deq_bits_data_instructionIndex = _writeQueueVec_fifo_3_empty ? writeQueueVec_3_enq_bits_data_instructionIndex : writeQueueVec_dataOut_3_data_instructionIndex;
  wire [3:0]         writeQueueVec_3_deq_bits_targetLane = _writeQueueVec_fifo_3_empty ? 4'h8 : writeQueueVec_dataOut_3_targetLane;
  wire               otherUnitTargetQueue_deq_valid;
  assign otherUnitTargetQueue_deq_valid = ~_otherUnitTargetQueue_fifo_empty;
  wire               otherUnitTargetQueue_deq_ready;
  wire               otherUnitTargetQueue_enq_ready = ~_otherUnitTargetQueue_fifo_full | otherUnitTargetQueue_deq_ready;
  wire               otherUnitTargetQueue_enq_valid;
  wire               otherUnitDataQueueVec_0_enq_ready = ~_otherUnitDataQueueVec_fifo_full;
  wire               otherUnitDataQueueVec_0_deq_ready;
  wire               otherUnitDataQueueVec_0_enq_valid;
  wire               otherUnitDataQueueVec_0_deq_valid = ~_otherUnitDataQueueVec_fifo_empty | otherUnitDataQueueVec_0_enq_valid;
  wire [31:0]        otherUnitDataQueueVec_0_deq_bits = _otherUnitDataQueueVec_fifo_empty ? otherUnitDataQueueVec_0_enq_bits : _otherUnitDataQueueVec_fifo_data_out;
  wire               otherUnitDataQueueVec_1_enq_ready = ~_otherUnitDataQueueVec_fifo_1_full;
  wire               otherUnitDataQueueVec_1_deq_ready;
  wire               otherUnitDataQueueVec_1_enq_valid;
  wire               otherUnitDataQueueVec_1_deq_valid = ~_otherUnitDataQueueVec_fifo_1_empty | otherUnitDataQueueVec_1_enq_valid;
  wire [31:0]        otherUnitDataQueueVec_1_deq_bits = _otherUnitDataQueueVec_fifo_1_empty ? otherUnitDataQueueVec_1_enq_bits : _otherUnitDataQueueVec_fifo_1_data_out;
  wire               otherUnitDataQueueVec_2_enq_ready = ~_otherUnitDataQueueVec_fifo_2_full;
  wire               otherUnitDataQueueVec_2_deq_ready;
  wire               otherUnitDataQueueVec_2_enq_valid;
  wire               otherUnitDataQueueVec_2_deq_valid = ~_otherUnitDataQueueVec_fifo_2_empty | otherUnitDataQueueVec_2_enq_valid;
  wire [31:0]        otherUnitDataQueueVec_2_deq_bits = _otherUnitDataQueueVec_fifo_2_empty ? otherUnitDataQueueVec_2_enq_bits : _otherUnitDataQueueVec_fifo_2_data_out;
  wire               otherUnitDataQueueVec_3_enq_ready = ~_otherUnitDataQueueVec_fifo_3_full;
  wire               otherUnitDataQueueVec_3_deq_ready;
  wire               otherUnitDataQueueVec_3_enq_valid;
  wire               otherUnitDataQueueVec_3_deq_valid = ~_otherUnitDataQueueVec_fifo_3_empty | otherUnitDataQueueVec_3_enq_valid;
  wire [31:0]        otherUnitDataQueueVec_3_deq_bits = _otherUnitDataQueueVec_fifo_3_empty ? otherUnitDataQueueVec_3_enq_bits : _otherUnitDataQueueVec_fifo_3_data_out;
  wire [3:0]         otherTryReadVrf = _otherUnit_vrfReadDataPorts_valid ? _otherUnit_status_targetLane : 4'h0;
  wire               vrfReadDataPorts_0_valid_0 = otherTryReadVrf[0] | _storeUnit_vrfReadDataPorts_0_valid;
  wire [4:0]         vrfReadDataPorts_0_bits_vs_0 = otherTryReadVrf[0] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_0_bits_vs;
  wire [5:0]         vrfReadDataPorts_0_bits_offset_0 = otherTryReadVrf[0] ? _otherUnit_vrfReadDataPorts_bits_offset : _storeUnit_vrfReadDataPorts_0_bits_offset;
  wire [2:0]         vrfReadDataPorts_0_bits_instructionIndex_0 = otherTryReadVrf[0] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_0_bits_instructionIndex;
  wire               otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_0_enq_valid = vrfReadResults_0_valid & ~otherUnitTargetQueue_empty;
  wire [3:0]         dataDeqFire;
  assign otherUnitDataQueueVec_0_deq_ready = dataDeqFire[0];
  wire               vrfReadDataPorts_1_valid_0 = otherTryReadVrf[1] | _storeUnit_vrfReadDataPorts_1_valid;
  wire [4:0]         vrfReadDataPorts_1_bits_vs_0 = otherTryReadVrf[1] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_1_bits_vs;
  wire [5:0]         vrfReadDataPorts_1_bits_offset_0 = otherTryReadVrf[1] ? _otherUnit_vrfReadDataPorts_bits_offset : _storeUnit_vrfReadDataPorts_1_bits_offset;
  wire [2:0]         vrfReadDataPorts_1_bits_instructionIndex_0 = otherTryReadVrf[1] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_1_bits_instructionIndex;
  assign otherUnitDataQueueVec_1_enq_valid = vrfReadResults_1_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_1_deq_ready = dataDeqFire[1];
  wire               vrfReadDataPorts_2_valid_0 = otherTryReadVrf[2] | _storeUnit_vrfReadDataPorts_2_valid;
  wire [4:0]         vrfReadDataPorts_2_bits_vs_0 = otherTryReadVrf[2] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_2_bits_vs;
  wire [5:0]         vrfReadDataPorts_2_bits_offset_0 = otherTryReadVrf[2] ? _otherUnit_vrfReadDataPorts_bits_offset : _storeUnit_vrfReadDataPorts_2_bits_offset;
  wire [2:0]         vrfReadDataPorts_2_bits_instructionIndex_0 = otherTryReadVrf[2] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_2_bits_instructionIndex;
  assign otherUnitDataQueueVec_2_enq_valid = vrfReadResults_2_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_2_deq_ready = dataDeqFire[2];
  wire               vrfReadDataPorts_3_valid_0 = otherTryReadVrf[3] | _storeUnit_vrfReadDataPorts_3_valid;
  wire [4:0]         vrfReadDataPorts_3_bits_vs_0 = otherTryReadVrf[3] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_3_bits_vs;
  wire [5:0]         vrfReadDataPorts_3_bits_offset_0 = otherTryReadVrf[3] ? _otherUnit_vrfReadDataPorts_bits_offset : _storeUnit_vrfReadDataPorts_3_bits_offset;
  wire [2:0]         vrfReadDataPorts_3_bits_instructionIndex_0 = otherTryReadVrf[3] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_3_bits_instructionIndex;
  assign otherUnitDataQueueVec_3_enq_valid = vrfReadResults_3_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_3_deq_ready = dataDeqFire[3];
  wire [1:0]         otherUnit_vrfReadDataPorts_ready_lo = {vrfReadDataPorts_1_ready_0, vrfReadDataPorts_0_ready_0};
  wire [1:0]         otherUnit_vrfReadDataPorts_ready_hi = {vrfReadDataPorts_3_ready_0, vrfReadDataPorts_2_ready_0};
  wire               otherUnit_vrfReadDataPorts_ready = (|(otherTryReadVrf & {otherUnit_vrfReadDataPorts_ready_hi, otherUnit_vrfReadDataPorts_ready_lo})) & otherUnitTargetQueue_enq_ready;
  assign otherUnitTargetQueue_enq_valid = otherUnit_vrfReadDataPorts_ready & _otherUnit_vrfReadDataPorts_valid;
  wire [3:0]         otherUnitTargetQueue_deq_bits;
  wire [1:0]         otherUnit_vrfReadResults_valid_lo = {otherUnitDataQueueVec_1_deq_valid, otherUnitDataQueueVec_0_deq_valid};
  wire [1:0]         otherUnit_vrfReadResults_valid_hi = {otherUnitDataQueueVec_3_deq_valid, otherUnitDataQueueVec_2_deq_valid};
  assign otherUnitTargetQueue_deq_ready = otherUnitTargetQueue_deq_valid & (|(otherUnitTargetQueue_deq_bits & {otherUnit_vrfReadResults_valid_hi, otherUnit_vrfReadResults_valid_lo}));
  assign dataDeqFire = otherUnitTargetQueue_deq_ready ? otherUnitTargetQueue_deq_bits : 4'h0;
  wire [3:0]         otherTryToWrite = _otherUnit_vrfWritePort_valid ? _otherUnit_status_targetLane : 4'h0;
  wire [1:0]         otherUnit_vrfWritePort_ready_lo = {writeQueueVec_1_enq_ready, writeQueueVec_0_enq_ready};
  wire [1:0]         otherUnit_vrfWritePort_ready_hi = {writeQueueVec_3_enq_ready, writeQueueVec_2_enq_ready};
  assign writeQueueVec_0_enq_valid = otherTryToWrite[0] | _loadUnit_vrfWritePort_0_valid;
  assign writeQueueVec_0_enq_bits_data_vd = otherTryToWrite[0] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_0_bits_vd;
  assign writeQueueVec_0_enq_bits_data_offset = otherTryToWrite[0] ? _otherUnit_vrfWritePort_bits_offset : _loadUnit_vrfWritePort_0_bits_offset;
  assign writeQueueVec_0_enq_bits_data_mask = otherTryToWrite[0] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_0_bits_mask;
  assign writeQueueVec_0_enq_bits_data_data = otherTryToWrite[0] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_0_bits_data;
  assign writeQueueVec_0_enq_bits_data_last = otherTryToWrite[0] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_0_enq_bits_data_instructionIndex = otherTryToWrite[0] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_0_bits_instructionIndex;
  assign writeQueueVec_1_enq_valid = otherTryToWrite[1] | _loadUnit_vrfWritePort_1_valid;
  assign writeQueueVec_1_enq_bits_data_vd = otherTryToWrite[1] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_1_bits_vd;
  assign writeQueueVec_1_enq_bits_data_offset = otherTryToWrite[1] ? _otherUnit_vrfWritePort_bits_offset : _loadUnit_vrfWritePort_1_bits_offset;
  assign writeQueueVec_1_enq_bits_data_mask = otherTryToWrite[1] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_1_bits_mask;
  assign writeQueueVec_1_enq_bits_data_data = otherTryToWrite[1] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_1_bits_data;
  assign writeQueueVec_1_enq_bits_data_last = otherTryToWrite[1] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_1_enq_bits_data_instructionIndex = otherTryToWrite[1] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_1_bits_instructionIndex;
  assign writeQueueVec_2_enq_valid = otherTryToWrite[2] | _loadUnit_vrfWritePort_2_valid;
  assign writeQueueVec_2_enq_bits_data_vd = otherTryToWrite[2] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_2_bits_vd;
  assign writeQueueVec_2_enq_bits_data_offset = otherTryToWrite[2] ? _otherUnit_vrfWritePort_bits_offset : _loadUnit_vrfWritePort_2_bits_offset;
  assign writeQueueVec_2_enq_bits_data_mask = otherTryToWrite[2] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_2_bits_mask;
  assign writeQueueVec_2_enq_bits_data_data = otherTryToWrite[2] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_2_bits_data;
  assign writeQueueVec_2_enq_bits_data_last = otherTryToWrite[2] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_2_enq_bits_data_instructionIndex = otherTryToWrite[2] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_2_bits_instructionIndex;
  assign writeQueueVec_3_enq_valid = otherTryToWrite[3] | _loadUnit_vrfWritePort_3_valid;
  assign writeQueueVec_3_enq_bits_data_vd = otherTryToWrite[3] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_3_bits_vd;
  assign writeQueueVec_3_enq_bits_data_offset = otherTryToWrite[3] ? _otherUnit_vrfWritePort_bits_offset : _loadUnit_vrfWritePort_3_bits_offset;
  assign writeQueueVec_3_enq_bits_data_mask = otherTryToWrite[3] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_3_bits_mask;
  assign writeQueueVec_3_enq_bits_data_data = otherTryToWrite[3] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_3_bits_data;
  assign writeQueueVec_3_enq_bits_data_last = otherTryToWrite[3] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_3_enq_bits_data_instructionIndex = otherTryToWrite[3] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_3_bits_instructionIndex;
  wire [7:0]         _GEN_130 = {5'h0, _loadUnit_status_instructionIndex};
  wire [7:0]         _GEN_131 = {5'h0, _otherUnit_status_instructionIndex};
  wire [7:0]         dataInMSHR = (_loadUnit_status_idle ? 8'h0 : 8'h1 << _GEN_130) | (_otherUnit_status_idle | _otherUnit_status_isStore ? 8'h0 : 8'h1 << _GEN_131);
  reg  [6:0]         queueCount_0;
  reg  [6:0]         queueCount_1;
  reg  [6:0]         queueCount_2;
  reg  [6:0]         queueCount_3;
  reg  [6:0]         queueCount_4;
  reg  [6:0]         queueCount_5;
  reg  [6:0]         queueCount_6;
  reg  [6:0]         queueCount_7;
  wire [7:0]         enqOH = 8'h1 << writeQueueVec_0_enq_bits_data_instructionIndex;
  wire [7:0]         queueEnq = _probeWire_slots_0_writeValid_T ? enqOH : 8'h0;
  wire               writeIndexQueue_deq_valid;
  assign writeIndexQueue_deq_valid = ~_writeIndexQueue_fifo_empty;
  wire               writeIndexQueue_enq_ready = ~_writeIndexQueue_fifo_full;
  wire               writeIndexQueue_enq_valid;
  assign writeIndexQueue_enq_valid = writeQueueVec_0_deq_ready & writeQueueVec_0_deq_valid;
  wire [2:0]         writeIndexQueue_deq_bits;
  wire [7:0]         queueDeq = writeIndexQueue_deq_ready & writeIndexQueue_deq_valid ? 8'h1 << writeIndexQueue_deq_bits : 8'h0;
  wire [6:0]         counterUpdate = queueEnq[0] ? 7'h1 : 7'h7F;
  wire [6:0]         counterUpdate_1 = queueEnq[1] ? 7'h1 : 7'h7F;
  wire [6:0]         counterUpdate_2 = queueEnq[2] ? 7'h1 : 7'h7F;
  wire [6:0]         counterUpdate_3 = queueEnq[3] ? 7'h1 : 7'h7F;
  wire [6:0]         counterUpdate_4 = queueEnq[4] ? 7'h1 : 7'h7F;
  wire [6:0]         counterUpdate_5 = queueEnq[5] ? 7'h1 : 7'h7F;
  wire [6:0]         counterUpdate_6 = queueEnq[6] ? 7'h1 : 7'h7F;
  wire [6:0]         counterUpdate_7 = queueEnq[7] ? 7'h1 : 7'h7F;
  wire [1:0]         dataInWriteQueue_0_lo_lo = {|queueCount_1, |queueCount_0};
  wire [1:0]         dataInWriteQueue_0_lo_hi = {|queueCount_3, |queueCount_2};
  wire [3:0]         dataInWriteQueue_0_lo = {dataInWriteQueue_0_lo_hi, dataInWriteQueue_0_lo_lo};
  wire [1:0]         dataInWriteQueue_0_hi_lo = {|queueCount_5, |queueCount_4};
  wire [1:0]         dataInWriteQueue_0_hi_hi = {|queueCount_7, |queueCount_6};
  wire [3:0]         dataInWriteQueue_0_hi = {dataInWriteQueue_0_hi_hi, dataInWriteQueue_0_hi_lo};
  reg  [6:0]         queueCount_0_1;
  reg  [6:0]         queueCount_1_1;
  reg  [6:0]         queueCount_2_1;
  reg  [6:0]         queueCount_3_1;
  reg  [6:0]         queueCount_4_1;
  reg  [6:0]         queueCount_5_1;
  reg  [6:0]         queueCount_6_1;
  reg  [6:0]         queueCount_7_1;
  wire [7:0]         enqOH_1 = 8'h1 << writeQueueVec_1_enq_bits_data_instructionIndex;
  wire [7:0]         queueEnq_1 = _probeWire_slots_1_writeValid_T ? enqOH_1 : 8'h0;
  wire               writeIndexQueue_1_deq_valid;
  assign writeIndexQueue_1_deq_valid = ~_writeIndexQueue_fifo_1_empty;
  wire               writeIndexQueue_1_enq_ready = ~_writeIndexQueue_fifo_1_full;
  wire               writeIndexQueue_1_enq_valid;
  assign writeIndexQueue_1_enq_valid = writeQueueVec_1_deq_ready & writeQueueVec_1_deq_valid;
  wire [2:0]         writeIndexQueue_1_deq_bits;
  wire [7:0]         queueDeq_1 = writeIndexQueue_1_deq_ready & writeIndexQueue_1_deq_valid ? 8'h1 << writeIndexQueue_1_deq_bits : 8'h0;
  wire [6:0]         counterUpdate_8 = queueEnq_1[0] ? 7'h1 : 7'h7F;
  wire [6:0]         counterUpdate_9 = queueEnq_1[1] ? 7'h1 : 7'h7F;
  wire [6:0]         counterUpdate_10 = queueEnq_1[2] ? 7'h1 : 7'h7F;
  wire [6:0]         counterUpdate_11 = queueEnq_1[3] ? 7'h1 : 7'h7F;
  wire [6:0]         counterUpdate_12 = queueEnq_1[4] ? 7'h1 : 7'h7F;
  wire [6:0]         counterUpdate_13 = queueEnq_1[5] ? 7'h1 : 7'h7F;
  wire [6:0]         counterUpdate_14 = queueEnq_1[6] ? 7'h1 : 7'h7F;
  wire [6:0]         counterUpdate_15 = queueEnq_1[7] ? 7'h1 : 7'h7F;
  wire [1:0]         dataInWriteQueue_1_lo_lo = {|queueCount_1_1, |queueCount_0_1};
  wire [1:0]         dataInWriteQueue_1_lo_hi = {|queueCount_3_1, |queueCount_2_1};
  wire [3:0]         dataInWriteQueue_1_lo = {dataInWriteQueue_1_lo_hi, dataInWriteQueue_1_lo_lo};
  wire [1:0]         dataInWriteQueue_1_hi_lo = {|queueCount_5_1, |queueCount_4_1};
  wire [1:0]         dataInWriteQueue_1_hi_hi = {|queueCount_7_1, |queueCount_6_1};
  wire [3:0]         dataInWriteQueue_1_hi = {dataInWriteQueue_1_hi_hi, dataInWriteQueue_1_hi_lo};
  reg  [6:0]         queueCount_0_2;
  reg  [6:0]         queueCount_1_2;
  reg  [6:0]         queueCount_2_2;
  reg  [6:0]         queueCount_3_2;
  reg  [6:0]         queueCount_4_2;
  reg  [6:0]         queueCount_5_2;
  reg  [6:0]         queueCount_6_2;
  reg  [6:0]         queueCount_7_2;
  wire [7:0]         enqOH_2 = 8'h1 << writeQueueVec_2_enq_bits_data_instructionIndex;
  wire [7:0]         queueEnq_2 = _probeWire_slots_2_writeValid_T ? enqOH_2 : 8'h0;
  wire               writeIndexQueue_2_deq_valid;
  assign writeIndexQueue_2_deq_valid = ~_writeIndexQueue_fifo_2_empty;
  wire               writeIndexQueue_2_enq_ready = ~_writeIndexQueue_fifo_2_full;
  wire               writeIndexQueue_2_enq_valid;
  assign writeIndexQueue_2_enq_valid = writeQueueVec_2_deq_ready & writeQueueVec_2_deq_valid;
  wire [2:0]         writeIndexQueue_2_deq_bits;
  wire [7:0]         queueDeq_2 = writeIndexQueue_2_deq_ready & writeIndexQueue_2_deq_valid ? 8'h1 << writeIndexQueue_2_deq_bits : 8'h0;
  wire [6:0]         counterUpdate_16 = queueEnq_2[0] ? 7'h1 : 7'h7F;
  wire [6:0]         counterUpdate_17 = queueEnq_2[1] ? 7'h1 : 7'h7F;
  wire [6:0]         counterUpdate_18 = queueEnq_2[2] ? 7'h1 : 7'h7F;
  wire [6:0]         counterUpdate_19 = queueEnq_2[3] ? 7'h1 : 7'h7F;
  wire [6:0]         counterUpdate_20 = queueEnq_2[4] ? 7'h1 : 7'h7F;
  wire [6:0]         counterUpdate_21 = queueEnq_2[5] ? 7'h1 : 7'h7F;
  wire [6:0]         counterUpdate_22 = queueEnq_2[6] ? 7'h1 : 7'h7F;
  wire [6:0]         counterUpdate_23 = queueEnq_2[7] ? 7'h1 : 7'h7F;
  wire [1:0]         dataInWriteQueue_2_lo_lo = {|queueCount_1_2, |queueCount_0_2};
  wire [1:0]         dataInWriteQueue_2_lo_hi = {|queueCount_3_2, |queueCount_2_2};
  wire [3:0]         dataInWriteQueue_2_lo = {dataInWriteQueue_2_lo_hi, dataInWriteQueue_2_lo_lo};
  wire [1:0]         dataInWriteQueue_2_hi_lo = {|queueCount_5_2, |queueCount_4_2};
  wire [1:0]         dataInWriteQueue_2_hi_hi = {|queueCount_7_2, |queueCount_6_2};
  wire [3:0]         dataInWriteQueue_2_hi = {dataInWriteQueue_2_hi_hi, dataInWriteQueue_2_hi_lo};
  reg  [6:0]         queueCount_0_3;
  reg  [6:0]         queueCount_1_3;
  reg  [6:0]         queueCount_2_3;
  reg  [6:0]         queueCount_3_3;
  reg  [6:0]         queueCount_4_3;
  reg  [6:0]         queueCount_5_3;
  reg  [6:0]         queueCount_6_3;
  reg  [6:0]         queueCount_7_3;
  wire [7:0]         enqOH_3 = 8'h1 << writeQueueVec_3_enq_bits_data_instructionIndex;
  wire [7:0]         queueEnq_3 = _probeWire_slots_3_writeValid_T ? enqOH_3 : 8'h0;
  wire               writeIndexQueue_3_deq_valid;
  assign writeIndexQueue_3_deq_valid = ~_writeIndexQueue_fifo_3_empty;
  wire               writeIndexQueue_3_enq_ready = ~_writeIndexQueue_fifo_3_full;
  wire               writeIndexQueue_3_enq_valid;
  assign writeIndexQueue_3_enq_valid = writeQueueVec_3_deq_ready & writeQueueVec_3_deq_valid;
  wire [2:0]         writeIndexQueue_3_deq_bits;
  wire [7:0]         queueDeq_3 = writeIndexQueue_3_deq_ready & writeIndexQueue_3_deq_valid ? 8'h1 << writeIndexQueue_3_deq_bits : 8'h0;
  wire [6:0]         counterUpdate_24 = queueEnq_3[0] ? 7'h1 : 7'h7F;
  wire [6:0]         counterUpdate_25 = queueEnq_3[1] ? 7'h1 : 7'h7F;
  wire [6:0]         counterUpdate_26 = queueEnq_3[2] ? 7'h1 : 7'h7F;
  wire [6:0]         counterUpdate_27 = queueEnq_3[3] ? 7'h1 : 7'h7F;
  wire [6:0]         counterUpdate_28 = queueEnq_3[4] ? 7'h1 : 7'h7F;
  wire [6:0]         counterUpdate_29 = queueEnq_3[5] ? 7'h1 : 7'h7F;
  wire [6:0]         counterUpdate_30 = queueEnq_3[6] ? 7'h1 : 7'h7F;
  wire [6:0]         counterUpdate_31 = queueEnq_3[7] ? 7'h1 : 7'h7F;
  wire [1:0]         dataInWriteQueue_3_lo_lo = {|queueCount_1_3, |queueCount_0_3};
  wire [1:0]         dataInWriteQueue_3_lo_hi = {|queueCount_3_3, |queueCount_2_3};
  wire [3:0]         dataInWriteQueue_3_lo = {dataInWriteQueue_3_lo_hi, dataInWriteQueue_3_lo_lo};
  wire [1:0]         dataInWriteQueue_3_hi_lo = {|queueCount_5_3, |queueCount_4_3};
  wire [1:0]         dataInWriteQueue_3_hi_hi = {|queueCount_7_3, |queueCount_6_3};
  wire [3:0]         dataInWriteQueue_3_hi = {dataInWriteQueue_3_hi_hi, dataInWriteQueue_3_hi_lo};
  wire               sourceQueue_deq_valid;
  assign sourceQueue_deq_valid = ~_sourceQueue_fifo_empty;
  wire               sourceQueue_enq_ready = ~_sourceQueue_fifo_full;
  wire               sourceQueue_enq_valid;
  wire               sourceQueue_deq_ready;
  wire               axi4Port_ar_valid_0 = _loadUnit_memRequest_valid & sourceQueue_enq_ready;
  wire               axi4Port_r_ready_0;
  assign sourceQueue_enq_valid = _loadUnit_memRequest_valid & axi4Port_ar_ready_0;
  assign sourceQueue_deq_ready = axi4Port_r_ready_0 & axi4Port_r_valid_0;
  assign dataQueue_deq_valid = ~_dataQueue_fifo_empty;
  wire               axi4Port_w_valid_0 = dataQueue_deq_valid;
  wire [127:0]       dataQueue_dataOut_data;
  wire [127:0]       axi4Port_w_bits_data_0 = dataQueue_deq_bits_data;
  wire [15:0]        dataQueue_dataOut_mask;
  wire [15:0]        axi4Port_w_bits_strb_0 = dataQueue_deq_bits_mask;
  wire [9:0]         dataQueue_dataOut_index;
  wire [31:0]        dataQueue_dataOut_address;
  wire [9:0]         dataQueue_enq_bits_index;
  wire [31:0]        dataQueue_enq_bits_address;
  wire [41:0]        dataQueue_dataIn_lo = {dataQueue_enq_bits_index, dataQueue_enq_bits_address};
  wire [127:0]       dataQueue_enq_bits_data;
  wire [15:0]        dataQueue_enq_bits_mask;
  wire [143:0]       dataQueue_dataIn_hi = {dataQueue_enq_bits_data, dataQueue_enq_bits_mask};
  wire [185:0]       dataQueue_dataIn = {dataQueue_dataIn_hi, dataQueue_dataIn_lo};
  assign dataQueue_dataOut_address = _dataQueue_fifo_data_out[31:0];
  assign dataQueue_dataOut_index = _dataQueue_fifo_data_out[41:32];
  assign dataQueue_dataOut_mask = _dataQueue_fifo_data_out[57:42];
  assign dataQueue_dataOut_data = _dataQueue_fifo_data_out[185:58];
  assign dataQueue_deq_bits_data = dataQueue_dataOut_data;
  assign dataQueue_deq_bits_mask = dataQueue_dataOut_mask;
  wire [9:0]         dataQueue_deq_bits_index = dataQueue_dataOut_index;
  wire [31:0]        dataQueue_deq_bits_address = dataQueue_dataOut_address;
  wire               dataQueue_enq_ready = ~_dataQueue_fifo_full;
  wire               dataQueue_enq_valid;
  wire               axi4Port_aw_valid_0 = _storeUnit_memRequest_valid & dataQueue_enq_ready;
  wire [1:0]         axi4Port_aw_bits_id_0 = _storeUnit_memRequest_bits_index[1:0];
  assign dataQueue_enq_valid = _storeUnit_memRequest_valid & axi4Port_aw_ready_0;
  wire               simpleSourceQueue_deq_valid;
  assign simpleSourceQueue_deq_valid = ~_simpleSourceQueue_fifo_empty;
  wire               simpleSourceQueue_enq_ready = ~_simpleSourceQueue_fifo_full;
  wire               simpleSourceQueue_enq_valid;
  wire               simpleSourceQueue_deq_ready;
  wire               simpleAccessPorts_ar_valid_0 = _otherUnit_memReadRequest_valid & simpleSourceQueue_enq_ready;
  wire               simpleAccessPorts_r_ready_0;
  assign simpleSourceQueue_enq_valid = _otherUnit_memReadRequest_valid & simpleAccessPorts_ar_ready_0;
  assign simpleSourceQueue_deq_ready = simpleAccessPorts_r_ready_0 & simpleAccessPorts_r_valid_0;
  assign simpleDataQueue_deq_valid = ~_simpleDataQueue_fifo_empty;
  wire               simpleAccessPorts_w_valid_0 = simpleDataQueue_deq_valid;
  wire [31:0]        simpleDataQueue_dataOut_data;
  wire [31:0]        simpleAccessPorts_w_bits_data_0 = simpleDataQueue_deq_bits_data;
  wire [3:0]         simpleDataQueue_dataOut_mask;
  wire [3:0]         simpleAccessPorts_w_bits_strb_0 = simpleDataQueue_deq_bits_mask;
  wire [7:0]         simpleDataQueue_dataOut_source;
  wire [31:0]        simpleDataQueue_dataOut_address;
  wire [1:0]         simpleDataQueue_dataOut_size;
  wire [31:0]        simpleDataQueue_enq_bits_address;
  wire [1:0]         simpleDataQueue_enq_bits_size;
  wire [33:0]        simpleDataQueue_dataIn_lo = {simpleDataQueue_enq_bits_address, simpleDataQueue_enq_bits_size};
  wire [31:0]        simpleDataQueue_enq_bits_data;
  wire [3:0]         simpleDataQueue_enq_bits_mask;
  wire [35:0]        simpleDataQueue_dataIn_hi_hi = {simpleDataQueue_enq_bits_data, simpleDataQueue_enq_bits_mask};
  wire [7:0]         simpleDataQueue_enq_bits_source;
  wire [43:0]        simpleDataQueue_dataIn_hi = {simpleDataQueue_dataIn_hi_hi, simpleDataQueue_enq_bits_source};
  wire [77:0]        simpleDataQueue_dataIn = {simpleDataQueue_dataIn_hi, simpleDataQueue_dataIn_lo};
  assign simpleDataQueue_dataOut_size = _simpleDataQueue_fifo_data_out[1:0];
  assign simpleDataQueue_dataOut_address = _simpleDataQueue_fifo_data_out[33:2];
  assign simpleDataQueue_dataOut_source = _simpleDataQueue_fifo_data_out[41:34];
  assign simpleDataQueue_dataOut_mask = _simpleDataQueue_fifo_data_out[45:42];
  assign simpleDataQueue_dataOut_data = _simpleDataQueue_fifo_data_out[77:46];
  assign simpleDataQueue_deq_bits_data = simpleDataQueue_dataOut_data;
  assign simpleDataQueue_deq_bits_mask = simpleDataQueue_dataOut_mask;
  wire [7:0]         simpleDataQueue_deq_bits_source = simpleDataQueue_dataOut_source;
  wire [31:0]        simpleDataQueue_deq_bits_address = simpleDataQueue_dataOut_address;
  wire [1:0]         simpleDataQueue_deq_bits_size = simpleDataQueue_dataOut_size;
  wire               simpleDataQueue_enq_ready = ~_simpleDataQueue_fifo_full;
  wire               simpleDataQueue_enq_valid;
  wire               simpleAccessPorts_aw_valid_0 = _otherUnit_memWriteRequest_valid & dataQueue_enq_ready;
  wire [2:0]         simpleAccessPorts_aw_bits_size_0 = {1'h0, _otherUnit_memWriteRequest_bits_size};
  wire [1:0]         simpleAccessPorts_aw_bits_id_0 = _otherUnit_memWriteRequest_bits_source[1:0];
  assign simpleDataQueue_enq_valid = _otherUnit_memWriteRequest_valid & simpleAccessPorts_aw_ready_0;
  wire [1:0]         tokenIO_offsetGroupRelease_lo = {_otherUnit_offsetRelease_1, _otherUnit_offsetRelease_0};
  wire [1:0]         tokenIO_offsetGroupRelease_hi = {_otherUnit_offsetRelease_3, _otherUnit_offsetRelease_2};
  wire               unitOrder =
    _loadUnit_status_instructionIndex == _storeUnit_status_instructionIndex | _loadUnit_status_instructionIndex[1:0] < _storeUnit_status_instructionIndex[1:0] ^ _loadUnit_status_instructionIndex[2] ^ _storeUnit_status_instructionIndex[2];
  wire               loadAddressConflict = _loadUnit_status_startAddress >= _storeUnit_status_startAddress & _loadUnit_status_startAddress <= _storeUnit_status_endAddress;
  wire               storeAddressConflict = _storeUnit_status_startAddress >= _loadUnit_status_startAddress & _storeUnit_status_startAddress <= _loadUnit_status_endAddress;
  wire               stallLoad = ~unitOrder & loadAddressConflict & ~_storeUnit_status_idle;
  wire               stallStore = unitOrder & storeAddressConflict & ~_loadUnit_status_idle;
  always @(posedge clock) begin
    if (reset) begin
      v0_0 <= 32'h0;
      v0_1 <= 32'h0;
      v0_2 <= 32'h0;
      v0_3 <= 32'h0;
      v0_4 <= 32'h0;
      v0_5 <= 32'h0;
      v0_6 <= 32'h0;
      v0_7 <= 32'h0;
      v0_8 <= 32'h0;
      v0_9 <= 32'h0;
      v0_10 <= 32'h0;
      v0_11 <= 32'h0;
      v0_12 <= 32'h0;
      v0_13 <= 32'h0;
      v0_14 <= 32'h0;
      v0_15 <= 32'h0;
      v0_16 <= 32'h0;
      v0_17 <= 32'h0;
      v0_18 <= 32'h0;
      v0_19 <= 32'h0;
      v0_20 <= 32'h0;
      v0_21 <= 32'h0;
      v0_22 <= 32'h0;
      v0_23 <= 32'h0;
      v0_24 <= 32'h0;
      v0_25 <= 32'h0;
      v0_26 <= 32'h0;
      v0_27 <= 32'h0;
      v0_28 <= 32'h0;
      v0_29 <= 32'h0;
      v0_30 <= 32'h0;
      v0_31 <= 32'h0;
      v0_32 <= 32'h0;
      v0_33 <= 32'h0;
      v0_34 <= 32'h0;
      v0_35 <= 32'h0;
      v0_36 <= 32'h0;
      v0_37 <= 32'h0;
      v0_38 <= 32'h0;
      v0_39 <= 32'h0;
      v0_40 <= 32'h0;
      v0_41 <= 32'h0;
      v0_42 <= 32'h0;
      v0_43 <= 32'h0;
      v0_44 <= 32'h0;
      v0_45 <= 32'h0;
      v0_46 <= 32'h0;
      v0_47 <= 32'h0;
      v0_48 <= 32'h0;
      v0_49 <= 32'h0;
      v0_50 <= 32'h0;
      v0_51 <= 32'h0;
      v0_52 <= 32'h0;
      v0_53 <= 32'h0;
      v0_54 <= 32'h0;
      v0_55 <= 32'h0;
      v0_56 <= 32'h0;
      v0_57 <= 32'h0;
      v0_58 <= 32'h0;
      v0_59 <= 32'h0;
      v0_60 <= 32'h0;
      v0_61 <= 32'h0;
      v0_62 <= 32'h0;
      v0_63 <= 32'h0;
      v0_64 <= 32'h0;
      v0_65 <= 32'h0;
      v0_66 <= 32'h0;
      v0_67 <= 32'h0;
      v0_68 <= 32'h0;
      v0_69 <= 32'h0;
      v0_70 <= 32'h0;
      v0_71 <= 32'h0;
      v0_72 <= 32'h0;
      v0_73 <= 32'h0;
      v0_74 <= 32'h0;
      v0_75 <= 32'h0;
      v0_76 <= 32'h0;
      v0_77 <= 32'h0;
      v0_78 <= 32'h0;
      v0_79 <= 32'h0;
      v0_80 <= 32'h0;
      v0_81 <= 32'h0;
      v0_82 <= 32'h0;
      v0_83 <= 32'h0;
      v0_84 <= 32'h0;
      v0_85 <= 32'h0;
      v0_86 <= 32'h0;
      v0_87 <= 32'h0;
      v0_88 <= 32'h0;
      v0_89 <= 32'h0;
      v0_90 <= 32'h0;
      v0_91 <= 32'h0;
      v0_92 <= 32'h0;
      v0_93 <= 32'h0;
      v0_94 <= 32'h0;
      v0_95 <= 32'h0;
      v0_96 <= 32'h0;
      v0_97 <= 32'h0;
      v0_98 <= 32'h0;
      v0_99 <= 32'h0;
      v0_100 <= 32'h0;
      v0_101 <= 32'h0;
      v0_102 <= 32'h0;
      v0_103 <= 32'h0;
      v0_104 <= 32'h0;
      v0_105 <= 32'h0;
      v0_106 <= 32'h0;
      v0_107 <= 32'h0;
      v0_108 <= 32'h0;
      v0_109 <= 32'h0;
      v0_110 <= 32'h0;
      v0_111 <= 32'h0;
      v0_112 <= 32'h0;
      v0_113 <= 32'h0;
      v0_114 <= 32'h0;
      v0_115 <= 32'h0;
      v0_116 <= 32'h0;
      v0_117 <= 32'h0;
      v0_118 <= 32'h0;
      v0_119 <= 32'h0;
      v0_120 <= 32'h0;
      v0_121 <= 32'h0;
      v0_122 <= 32'h0;
      v0_123 <= 32'h0;
      v0_124 <= 32'h0;
      v0_125 <= 32'h0;
      v0_126 <= 32'h0;
      v0_127 <= 32'h0;
      v0_128 <= 32'h0;
      v0_129 <= 32'h0;
      v0_130 <= 32'h0;
      v0_131 <= 32'h0;
      v0_132 <= 32'h0;
      v0_133 <= 32'h0;
      v0_134 <= 32'h0;
      v0_135 <= 32'h0;
      v0_136 <= 32'h0;
      v0_137 <= 32'h0;
      v0_138 <= 32'h0;
      v0_139 <= 32'h0;
      v0_140 <= 32'h0;
      v0_141 <= 32'h0;
      v0_142 <= 32'h0;
      v0_143 <= 32'h0;
      v0_144 <= 32'h0;
      v0_145 <= 32'h0;
      v0_146 <= 32'h0;
      v0_147 <= 32'h0;
      v0_148 <= 32'h0;
      v0_149 <= 32'h0;
      v0_150 <= 32'h0;
      v0_151 <= 32'h0;
      v0_152 <= 32'h0;
      v0_153 <= 32'h0;
      v0_154 <= 32'h0;
      v0_155 <= 32'h0;
      v0_156 <= 32'h0;
      v0_157 <= 32'h0;
      v0_158 <= 32'h0;
      v0_159 <= 32'h0;
      v0_160 <= 32'h0;
      v0_161 <= 32'h0;
      v0_162 <= 32'h0;
      v0_163 <= 32'h0;
      v0_164 <= 32'h0;
      v0_165 <= 32'h0;
      v0_166 <= 32'h0;
      v0_167 <= 32'h0;
      v0_168 <= 32'h0;
      v0_169 <= 32'h0;
      v0_170 <= 32'h0;
      v0_171 <= 32'h0;
      v0_172 <= 32'h0;
      v0_173 <= 32'h0;
      v0_174 <= 32'h0;
      v0_175 <= 32'h0;
      v0_176 <= 32'h0;
      v0_177 <= 32'h0;
      v0_178 <= 32'h0;
      v0_179 <= 32'h0;
      v0_180 <= 32'h0;
      v0_181 <= 32'h0;
      v0_182 <= 32'h0;
      v0_183 <= 32'h0;
      v0_184 <= 32'h0;
      v0_185 <= 32'h0;
      v0_186 <= 32'h0;
      v0_187 <= 32'h0;
      v0_188 <= 32'h0;
      v0_189 <= 32'h0;
      v0_190 <= 32'h0;
      v0_191 <= 32'h0;
      v0_192 <= 32'h0;
      v0_193 <= 32'h0;
      v0_194 <= 32'h0;
      v0_195 <= 32'h0;
      v0_196 <= 32'h0;
      v0_197 <= 32'h0;
      v0_198 <= 32'h0;
      v0_199 <= 32'h0;
      v0_200 <= 32'h0;
      v0_201 <= 32'h0;
      v0_202 <= 32'h0;
      v0_203 <= 32'h0;
      v0_204 <= 32'h0;
      v0_205 <= 32'h0;
      v0_206 <= 32'h0;
      v0_207 <= 32'h0;
      v0_208 <= 32'h0;
      v0_209 <= 32'h0;
      v0_210 <= 32'h0;
      v0_211 <= 32'h0;
      v0_212 <= 32'h0;
      v0_213 <= 32'h0;
      v0_214 <= 32'h0;
      v0_215 <= 32'h0;
      v0_216 <= 32'h0;
      v0_217 <= 32'h0;
      v0_218 <= 32'h0;
      v0_219 <= 32'h0;
      v0_220 <= 32'h0;
      v0_221 <= 32'h0;
      v0_222 <= 32'h0;
      v0_223 <= 32'h0;
      v0_224 <= 32'h0;
      v0_225 <= 32'h0;
      v0_226 <= 32'h0;
      v0_227 <= 32'h0;
      v0_228 <= 32'h0;
      v0_229 <= 32'h0;
      v0_230 <= 32'h0;
      v0_231 <= 32'h0;
      v0_232 <= 32'h0;
      v0_233 <= 32'h0;
      v0_234 <= 32'h0;
      v0_235 <= 32'h0;
      v0_236 <= 32'h0;
      v0_237 <= 32'h0;
      v0_238 <= 32'h0;
      v0_239 <= 32'h0;
      v0_240 <= 32'h0;
      v0_241 <= 32'h0;
      v0_242 <= 32'h0;
      v0_243 <= 32'h0;
      v0_244 <= 32'h0;
      v0_245 <= 32'h0;
      v0_246 <= 32'h0;
      v0_247 <= 32'h0;
      v0_248 <= 32'h0;
      v0_249 <= 32'h0;
      v0_250 <= 32'h0;
      v0_251 <= 32'h0;
      v0_252 <= 32'h0;
      v0_253 <= 32'h0;
      v0_254 <= 32'h0;
      v0_255 <= 32'h0;
      queueCount_0 <= 7'h0;
      queueCount_1 <= 7'h0;
      queueCount_2 <= 7'h0;
      queueCount_3 <= 7'h0;
      queueCount_4 <= 7'h0;
      queueCount_5 <= 7'h0;
      queueCount_6 <= 7'h0;
      queueCount_7 <= 7'h0;
      queueCount_0_1 <= 7'h0;
      queueCount_1_1 <= 7'h0;
      queueCount_2_1 <= 7'h0;
      queueCount_3_1 <= 7'h0;
      queueCount_4_1 <= 7'h0;
      queueCount_5_1 <= 7'h0;
      queueCount_6_1 <= 7'h0;
      queueCount_7_1 <= 7'h0;
      queueCount_0_2 <= 7'h0;
      queueCount_1_2 <= 7'h0;
      queueCount_2_2 <= 7'h0;
      queueCount_3_2 <= 7'h0;
      queueCount_4_2 <= 7'h0;
      queueCount_5_2 <= 7'h0;
      queueCount_6_2 <= 7'h0;
      queueCount_7_2 <= 7'h0;
      queueCount_0_3 <= 7'h0;
      queueCount_1_3 <= 7'h0;
      queueCount_2_3 <= 7'h0;
      queueCount_3_3 <= 7'h0;
      queueCount_4_3 <= 7'h0;
      queueCount_5_3 <= 7'h0;
      queueCount_6_3 <= 7'h0;
      queueCount_7_3 <= 7'h0;
    end
    else begin
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h0)
        v0_0 <= v0_0 & ~maskExt | maskExt & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h0)
        v0_1 <= v0_1 & ~maskExt_1 | maskExt_1 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h0)
        v0_2 <= v0_2 & ~maskExt_2 | maskExt_2 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h0)
        v0_3 <= v0_3 & ~maskExt_3 | maskExt_3 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h1)
        v0_4 <= v0_4 & ~maskExt_4 | maskExt_4 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h1)
        v0_5 <= v0_5 & ~maskExt_5 | maskExt_5 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h1)
        v0_6 <= v0_6 & ~maskExt_6 | maskExt_6 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h1)
        v0_7 <= v0_7 & ~maskExt_7 | maskExt_7 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h2)
        v0_8 <= v0_8 & ~maskExt_8 | maskExt_8 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h2)
        v0_9 <= v0_9 & ~maskExt_9 | maskExt_9 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h2)
        v0_10 <= v0_10 & ~maskExt_10 | maskExt_10 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h2)
        v0_11 <= v0_11 & ~maskExt_11 | maskExt_11 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h3)
        v0_12 <= v0_12 & ~maskExt_12 | maskExt_12 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h3)
        v0_13 <= v0_13 & ~maskExt_13 | maskExt_13 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h3)
        v0_14 <= v0_14 & ~maskExt_14 | maskExt_14 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h3)
        v0_15 <= v0_15 & ~maskExt_15 | maskExt_15 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h4)
        v0_16 <= v0_16 & ~maskExt_16 | maskExt_16 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h4)
        v0_17 <= v0_17 & ~maskExt_17 | maskExt_17 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h4)
        v0_18 <= v0_18 & ~maskExt_18 | maskExt_18 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h4)
        v0_19 <= v0_19 & ~maskExt_19 | maskExt_19 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h5)
        v0_20 <= v0_20 & ~maskExt_20 | maskExt_20 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h5)
        v0_21 <= v0_21 & ~maskExt_21 | maskExt_21 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h5)
        v0_22 <= v0_22 & ~maskExt_22 | maskExt_22 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h5)
        v0_23 <= v0_23 & ~maskExt_23 | maskExt_23 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h6)
        v0_24 <= v0_24 & ~maskExt_24 | maskExt_24 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h6)
        v0_25 <= v0_25 & ~maskExt_25 | maskExt_25 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h6)
        v0_26 <= v0_26 & ~maskExt_26 | maskExt_26 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h6)
        v0_27 <= v0_27 & ~maskExt_27 | maskExt_27 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h7)
        v0_28 <= v0_28 & ~maskExt_28 | maskExt_28 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h7)
        v0_29 <= v0_29 & ~maskExt_29 | maskExt_29 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h7)
        v0_30 <= v0_30 & ~maskExt_30 | maskExt_30 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h7)
        v0_31 <= v0_31 & ~maskExt_31 | maskExt_31 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h8)
        v0_32 <= v0_32 & ~maskExt_32 | maskExt_32 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h8)
        v0_33 <= v0_33 & ~maskExt_33 | maskExt_33 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h8)
        v0_34 <= v0_34 & ~maskExt_34 | maskExt_34 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h8)
        v0_35 <= v0_35 & ~maskExt_35 | maskExt_35 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h9)
        v0_36 <= v0_36 & ~maskExt_36 | maskExt_36 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h9)
        v0_37 <= v0_37 & ~maskExt_37 | maskExt_37 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h9)
        v0_38 <= v0_38 & ~maskExt_38 | maskExt_38 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h9)
        v0_39 <= v0_39 & ~maskExt_39 | maskExt_39 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'hA)
        v0_40 <= v0_40 & ~maskExt_40 | maskExt_40 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'hA)
        v0_41 <= v0_41 & ~maskExt_41 | maskExt_41 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'hA)
        v0_42 <= v0_42 & ~maskExt_42 | maskExt_42 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'hA)
        v0_43 <= v0_43 & ~maskExt_43 | maskExt_43 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'hB)
        v0_44 <= v0_44 & ~maskExt_44 | maskExt_44 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'hB)
        v0_45 <= v0_45 & ~maskExt_45 | maskExt_45 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'hB)
        v0_46 <= v0_46 & ~maskExt_46 | maskExt_46 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'hB)
        v0_47 <= v0_47 & ~maskExt_47 | maskExt_47 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'hC)
        v0_48 <= v0_48 & ~maskExt_48 | maskExt_48 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'hC)
        v0_49 <= v0_49 & ~maskExt_49 | maskExt_49 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'hC)
        v0_50 <= v0_50 & ~maskExt_50 | maskExt_50 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'hC)
        v0_51 <= v0_51 & ~maskExt_51 | maskExt_51 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'hD)
        v0_52 <= v0_52 & ~maskExt_52 | maskExt_52 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'hD)
        v0_53 <= v0_53 & ~maskExt_53 | maskExt_53 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'hD)
        v0_54 <= v0_54 & ~maskExt_54 | maskExt_54 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'hD)
        v0_55 <= v0_55 & ~maskExt_55 | maskExt_55 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'hE)
        v0_56 <= v0_56 & ~maskExt_56 | maskExt_56 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'hE)
        v0_57 <= v0_57 & ~maskExt_57 | maskExt_57 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'hE)
        v0_58 <= v0_58 & ~maskExt_58 | maskExt_58 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'hE)
        v0_59 <= v0_59 & ~maskExt_59 | maskExt_59 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'hF)
        v0_60 <= v0_60 & ~maskExt_60 | maskExt_60 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'hF)
        v0_61 <= v0_61 & ~maskExt_61 | maskExt_61 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'hF)
        v0_62 <= v0_62 & ~maskExt_62 | maskExt_62 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'hF)
        v0_63 <= v0_63 & ~maskExt_63 | maskExt_63 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h10)
        v0_64 <= v0_64 & ~maskExt_64 | maskExt_64 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h10)
        v0_65 <= v0_65 & ~maskExt_65 | maskExt_65 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h10)
        v0_66 <= v0_66 & ~maskExt_66 | maskExt_66 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h10)
        v0_67 <= v0_67 & ~maskExt_67 | maskExt_67 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h11)
        v0_68 <= v0_68 & ~maskExt_68 | maskExt_68 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h11)
        v0_69 <= v0_69 & ~maskExt_69 | maskExt_69 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h11)
        v0_70 <= v0_70 & ~maskExt_70 | maskExt_70 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h11)
        v0_71 <= v0_71 & ~maskExt_71 | maskExt_71 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h12)
        v0_72 <= v0_72 & ~maskExt_72 | maskExt_72 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h12)
        v0_73 <= v0_73 & ~maskExt_73 | maskExt_73 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h12)
        v0_74 <= v0_74 & ~maskExt_74 | maskExt_74 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h12)
        v0_75 <= v0_75 & ~maskExt_75 | maskExt_75 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h13)
        v0_76 <= v0_76 & ~maskExt_76 | maskExt_76 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h13)
        v0_77 <= v0_77 & ~maskExt_77 | maskExt_77 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h13)
        v0_78 <= v0_78 & ~maskExt_78 | maskExt_78 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h13)
        v0_79 <= v0_79 & ~maskExt_79 | maskExt_79 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h14)
        v0_80 <= v0_80 & ~maskExt_80 | maskExt_80 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h14)
        v0_81 <= v0_81 & ~maskExt_81 | maskExt_81 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h14)
        v0_82 <= v0_82 & ~maskExt_82 | maskExt_82 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h14)
        v0_83 <= v0_83 & ~maskExt_83 | maskExt_83 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h15)
        v0_84 <= v0_84 & ~maskExt_84 | maskExt_84 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h15)
        v0_85 <= v0_85 & ~maskExt_85 | maskExt_85 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h15)
        v0_86 <= v0_86 & ~maskExt_86 | maskExt_86 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h15)
        v0_87 <= v0_87 & ~maskExt_87 | maskExt_87 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h16)
        v0_88 <= v0_88 & ~maskExt_88 | maskExt_88 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h16)
        v0_89 <= v0_89 & ~maskExt_89 | maskExt_89 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h16)
        v0_90 <= v0_90 & ~maskExt_90 | maskExt_90 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h16)
        v0_91 <= v0_91 & ~maskExt_91 | maskExt_91 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h17)
        v0_92 <= v0_92 & ~maskExt_92 | maskExt_92 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h17)
        v0_93 <= v0_93 & ~maskExt_93 | maskExt_93 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h17)
        v0_94 <= v0_94 & ~maskExt_94 | maskExt_94 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h17)
        v0_95 <= v0_95 & ~maskExt_95 | maskExt_95 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h18)
        v0_96 <= v0_96 & ~maskExt_96 | maskExt_96 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h18)
        v0_97 <= v0_97 & ~maskExt_97 | maskExt_97 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h18)
        v0_98 <= v0_98 & ~maskExt_98 | maskExt_98 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h18)
        v0_99 <= v0_99 & ~maskExt_99 | maskExt_99 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h19)
        v0_100 <= v0_100 & ~maskExt_100 | maskExt_100 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h19)
        v0_101 <= v0_101 & ~maskExt_101 | maskExt_101 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h19)
        v0_102 <= v0_102 & ~maskExt_102 | maskExt_102 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h19)
        v0_103 <= v0_103 & ~maskExt_103 | maskExt_103 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h1A)
        v0_104 <= v0_104 & ~maskExt_104 | maskExt_104 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h1A)
        v0_105 <= v0_105 & ~maskExt_105 | maskExt_105 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h1A)
        v0_106 <= v0_106 & ~maskExt_106 | maskExt_106 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h1A)
        v0_107 <= v0_107 & ~maskExt_107 | maskExt_107 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h1B)
        v0_108 <= v0_108 & ~maskExt_108 | maskExt_108 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h1B)
        v0_109 <= v0_109 & ~maskExt_109 | maskExt_109 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h1B)
        v0_110 <= v0_110 & ~maskExt_110 | maskExt_110 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h1B)
        v0_111 <= v0_111 & ~maskExt_111 | maskExt_111 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h1C)
        v0_112 <= v0_112 & ~maskExt_112 | maskExt_112 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h1C)
        v0_113 <= v0_113 & ~maskExt_113 | maskExt_113 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h1C)
        v0_114 <= v0_114 & ~maskExt_114 | maskExt_114 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h1C)
        v0_115 <= v0_115 & ~maskExt_115 | maskExt_115 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h1D)
        v0_116 <= v0_116 & ~maskExt_116 | maskExt_116 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h1D)
        v0_117 <= v0_117 & ~maskExt_117 | maskExt_117 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h1D)
        v0_118 <= v0_118 & ~maskExt_118 | maskExt_118 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h1D)
        v0_119 <= v0_119 & ~maskExt_119 | maskExt_119 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h1E)
        v0_120 <= v0_120 & ~maskExt_120 | maskExt_120 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h1E)
        v0_121 <= v0_121 & ~maskExt_121 | maskExt_121 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h1E)
        v0_122 <= v0_122 & ~maskExt_122 | maskExt_122 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h1E)
        v0_123 <= v0_123 & ~maskExt_123 | maskExt_123 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h1F)
        v0_124 <= v0_124 & ~maskExt_124 | maskExt_124 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h1F)
        v0_125 <= v0_125 & ~maskExt_125 | maskExt_125 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h1F)
        v0_126 <= v0_126 & ~maskExt_126 | maskExt_126 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h1F)
        v0_127 <= v0_127 & ~maskExt_127 | maskExt_127 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h20)
        v0_128 <= v0_128 & ~maskExt_128 | maskExt_128 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h20)
        v0_129 <= v0_129 & ~maskExt_129 | maskExt_129 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h20)
        v0_130 <= v0_130 & ~maskExt_130 | maskExt_130 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h20)
        v0_131 <= v0_131 & ~maskExt_131 | maskExt_131 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h21)
        v0_132 <= v0_132 & ~maskExt_132 | maskExt_132 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h21)
        v0_133 <= v0_133 & ~maskExt_133 | maskExt_133 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h21)
        v0_134 <= v0_134 & ~maskExt_134 | maskExt_134 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h21)
        v0_135 <= v0_135 & ~maskExt_135 | maskExt_135 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h22)
        v0_136 <= v0_136 & ~maskExt_136 | maskExt_136 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h22)
        v0_137 <= v0_137 & ~maskExt_137 | maskExt_137 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h22)
        v0_138 <= v0_138 & ~maskExt_138 | maskExt_138 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h22)
        v0_139 <= v0_139 & ~maskExt_139 | maskExt_139 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h23)
        v0_140 <= v0_140 & ~maskExt_140 | maskExt_140 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h23)
        v0_141 <= v0_141 & ~maskExt_141 | maskExt_141 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h23)
        v0_142 <= v0_142 & ~maskExt_142 | maskExt_142 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h23)
        v0_143 <= v0_143 & ~maskExt_143 | maskExt_143 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h24)
        v0_144 <= v0_144 & ~maskExt_144 | maskExt_144 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h24)
        v0_145 <= v0_145 & ~maskExt_145 | maskExt_145 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h24)
        v0_146 <= v0_146 & ~maskExt_146 | maskExt_146 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h24)
        v0_147 <= v0_147 & ~maskExt_147 | maskExt_147 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h25)
        v0_148 <= v0_148 & ~maskExt_148 | maskExt_148 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h25)
        v0_149 <= v0_149 & ~maskExt_149 | maskExt_149 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h25)
        v0_150 <= v0_150 & ~maskExt_150 | maskExt_150 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h25)
        v0_151 <= v0_151 & ~maskExt_151 | maskExt_151 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h26)
        v0_152 <= v0_152 & ~maskExt_152 | maskExt_152 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h26)
        v0_153 <= v0_153 & ~maskExt_153 | maskExt_153 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h26)
        v0_154 <= v0_154 & ~maskExt_154 | maskExt_154 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h26)
        v0_155 <= v0_155 & ~maskExt_155 | maskExt_155 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h27)
        v0_156 <= v0_156 & ~maskExt_156 | maskExt_156 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h27)
        v0_157 <= v0_157 & ~maskExt_157 | maskExt_157 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h27)
        v0_158 <= v0_158 & ~maskExt_158 | maskExt_158 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h27)
        v0_159 <= v0_159 & ~maskExt_159 | maskExt_159 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h28)
        v0_160 <= v0_160 & ~maskExt_160 | maskExt_160 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h28)
        v0_161 <= v0_161 & ~maskExt_161 | maskExt_161 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h28)
        v0_162 <= v0_162 & ~maskExt_162 | maskExt_162 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h28)
        v0_163 <= v0_163 & ~maskExt_163 | maskExt_163 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h29)
        v0_164 <= v0_164 & ~maskExt_164 | maskExt_164 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h29)
        v0_165 <= v0_165 & ~maskExt_165 | maskExt_165 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h29)
        v0_166 <= v0_166 & ~maskExt_166 | maskExt_166 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h29)
        v0_167 <= v0_167 & ~maskExt_167 | maskExt_167 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h2A)
        v0_168 <= v0_168 & ~maskExt_168 | maskExt_168 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h2A)
        v0_169 <= v0_169 & ~maskExt_169 | maskExt_169 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h2A)
        v0_170 <= v0_170 & ~maskExt_170 | maskExt_170 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h2A)
        v0_171 <= v0_171 & ~maskExt_171 | maskExt_171 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h2B)
        v0_172 <= v0_172 & ~maskExt_172 | maskExt_172 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h2B)
        v0_173 <= v0_173 & ~maskExt_173 | maskExt_173 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h2B)
        v0_174 <= v0_174 & ~maskExt_174 | maskExt_174 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h2B)
        v0_175 <= v0_175 & ~maskExt_175 | maskExt_175 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h2C)
        v0_176 <= v0_176 & ~maskExt_176 | maskExt_176 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h2C)
        v0_177 <= v0_177 & ~maskExt_177 | maskExt_177 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h2C)
        v0_178 <= v0_178 & ~maskExt_178 | maskExt_178 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h2C)
        v0_179 <= v0_179 & ~maskExt_179 | maskExt_179 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h2D)
        v0_180 <= v0_180 & ~maskExt_180 | maskExt_180 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h2D)
        v0_181 <= v0_181 & ~maskExt_181 | maskExt_181 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h2D)
        v0_182 <= v0_182 & ~maskExt_182 | maskExt_182 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h2D)
        v0_183 <= v0_183 & ~maskExt_183 | maskExt_183 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h2E)
        v0_184 <= v0_184 & ~maskExt_184 | maskExt_184 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h2E)
        v0_185 <= v0_185 & ~maskExt_185 | maskExt_185 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h2E)
        v0_186 <= v0_186 & ~maskExt_186 | maskExt_186 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h2E)
        v0_187 <= v0_187 & ~maskExt_187 | maskExt_187 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h2F)
        v0_188 <= v0_188 & ~maskExt_188 | maskExt_188 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h2F)
        v0_189 <= v0_189 & ~maskExt_189 | maskExt_189 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h2F)
        v0_190 <= v0_190 & ~maskExt_190 | maskExt_190 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h2F)
        v0_191 <= v0_191 & ~maskExt_191 | maskExt_191 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h30)
        v0_192 <= v0_192 & ~maskExt_192 | maskExt_192 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h30)
        v0_193 <= v0_193 & ~maskExt_193 | maskExt_193 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h30)
        v0_194 <= v0_194 & ~maskExt_194 | maskExt_194 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h30)
        v0_195 <= v0_195 & ~maskExt_195 | maskExt_195 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h31)
        v0_196 <= v0_196 & ~maskExt_196 | maskExt_196 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h31)
        v0_197 <= v0_197 & ~maskExt_197 | maskExt_197 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h31)
        v0_198 <= v0_198 & ~maskExt_198 | maskExt_198 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h31)
        v0_199 <= v0_199 & ~maskExt_199 | maskExt_199 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h32)
        v0_200 <= v0_200 & ~maskExt_200 | maskExt_200 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h32)
        v0_201 <= v0_201 & ~maskExt_201 | maskExt_201 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h32)
        v0_202 <= v0_202 & ~maskExt_202 | maskExt_202 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h32)
        v0_203 <= v0_203 & ~maskExt_203 | maskExt_203 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h33)
        v0_204 <= v0_204 & ~maskExt_204 | maskExt_204 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h33)
        v0_205 <= v0_205 & ~maskExt_205 | maskExt_205 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h33)
        v0_206 <= v0_206 & ~maskExt_206 | maskExt_206 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h33)
        v0_207 <= v0_207 & ~maskExt_207 | maskExt_207 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h34)
        v0_208 <= v0_208 & ~maskExt_208 | maskExt_208 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h34)
        v0_209 <= v0_209 & ~maskExt_209 | maskExt_209 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h34)
        v0_210 <= v0_210 & ~maskExt_210 | maskExt_210 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h34)
        v0_211 <= v0_211 & ~maskExt_211 | maskExt_211 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h35)
        v0_212 <= v0_212 & ~maskExt_212 | maskExt_212 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h35)
        v0_213 <= v0_213 & ~maskExt_213 | maskExt_213 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h35)
        v0_214 <= v0_214 & ~maskExt_214 | maskExt_214 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h35)
        v0_215 <= v0_215 & ~maskExt_215 | maskExt_215 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h36)
        v0_216 <= v0_216 & ~maskExt_216 | maskExt_216 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h36)
        v0_217 <= v0_217 & ~maskExt_217 | maskExt_217 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h36)
        v0_218 <= v0_218 & ~maskExt_218 | maskExt_218 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h36)
        v0_219 <= v0_219 & ~maskExt_219 | maskExt_219 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h37)
        v0_220 <= v0_220 & ~maskExt_220 | maskExt_220 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h37)
        v0_221 <= v0_221 & ~maskExt_221 | maskExt_221 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h37)
        v0_222 <= v0_222 & ~maskExt_222 | maskExt_222 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h37)
        v0_223 <= v0_223 & ~maskExt_223 | maskExt_223 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h38)
        v0_224 <= v0_224 & ~maskExt_224 | maskExt_224 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h38)
        v0_225 <= v0_225 & ~maskExt_225 | maskExt_225 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h38)
        v0_226 <= v0_226 & ~maskExt_226 | maskExt_226 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h38)
        v0_227 <= v0_227 & ~maskExt_227 | maskExt_227 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h39)
        v0_228 <= v0_228 & ~maskExt_228 | maskExt_228 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h39)
        v0_229 <= v0_229 & ~maskExt_229 | maskExt_229 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h39)
        v0_230 <= v0_230 & ~maskExt_230 | maskExt_230 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h39)
        v0_231 <= v0_231 & ~maskExt_231 | maskExt_231 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h3A)
        v0_232 <= v0_232 & ~maskExt_232 | maskExt_232 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h3A)
        v0_233 <= v0_233 & ~maskExt_233 | maskExt_233 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h3A)
        v0_234 <= v0_234 & ~maskExt_234 | maskExt_234 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h3A)
        v0_235 <= v0_235 & ~maskExt_235 | maskExt_235 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h3B)
        v0_236 <= v0_236 & ~maskExt_236 | maskExt_236 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h3B)
        v0_237 <= v0_237 & ~maskExt_237 | maskExt_237 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h3B)
        v0_238 <= v0_238 & ~maskExt_238 | maskExt_238 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h3B)
        v0_239 <= v0_239 & ~maskExt_239 | maskExt_239 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h3C)
        v0_240 <= v0_240 & ~maskExt_240 | maskExt_240 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h3C)
        v0_241 <= v0_241 & ~maskExt_241 | maskExt_241 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h3C)
        v0_242 <= v0_242 & ~maskExt_242 | maskExt_242 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h3C)
        v0_243 <= v0_243 & ~maskExt_243 | maskExt_243 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h3D)
        v0_244 <= v0_244 & ~maskExt_244 | maskExt_244 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h3D)
        v0_245 <= v0_245 & ~maskExt_245 | maskExt_245 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h3D)
        v0_246 <= v0_246 & ~maskExt_246 | maskExt_246 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h3D)
        v0_247 <= v0_247 & ~maskExt_247 | maskExt_247 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h3E)
        v0_248 <= v0_248 & ~maskExt_248 | maskExt_248 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h3E)
        v0_249 <= v0_249 & ~maskExt_249 | maskExt_249 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h3E)
        v0_250 <= v0_250 & ~maskExt_250 | maskExt_250 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h3E)
        v0_251 <= v0_251 & ~maskExt_251 | maskExt_251 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & (&v0UpdateVec_0_bits_offset))
        v0_252 <= v0_252 & ~maskExt_252 | maskExt_252 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & (&v0UpdateVec_1_bits_offset))
        v0_253 <= v0_253 & ~maskExt_253 | maskExt_253 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & (&v0UpdateVec_2_bits_offset))
        v0_254 <= v0_254 & ~maskExt_254 | maskExt_254 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & (&v0UpdateVec_3_bits_offset))
        v0_255 <= v0_255 & ~maskExt_255 | maskExt_255 & v0UpdateVec_3_bits_data;
      if (queueEnq[0] ^ queueDeq[0])
        queueCount_0 <= queueCount_0 + counterUpdate;
      if (queueEnq[1] ^ queueDeq[1])
        queueCount_1 <= queueCount_1 + counterUpdate_1;
      if (queueEnq[2] ^ queueDeq[2])
        queueCount_2 <= queueCount_2 + counterUpdate_2;
      if (queueEnq[3] ^ queueDeq[3])
        queueCount_3 <= queueCount_3 + counterUpdate_3;
      if (queueEnq[4] ^ queueDeq[4])
        queueCount_4 <= queueCount_4 + counterUpdate_4;
      if (queueEnq[5] ^ queueDeq[5])
        queueCount_5 <= queueCount_5 + counterUpdate_5;
      if (queueEnq[6] ^ queueDeq[6])
        queueCount_6 <= queueCount_6 + counterUpdate_6;
      if (queueEnq[7] ^ queueDeq[7])
        queueCount_7 <= queueCount_7 + counterUpdate_7;
      if (queueEnq_1[0] ^ queueDeq_1[0])
        queueCount_0_1 <= queueCount_0_1 + counterUpdate_8;
      if (queueEnq_1[1] ^ queueDeq_1[1])
        queueCount_1_1 <= queueCount_1_1 + counterUpdate_9;
      if (queueEnq_1[2] ^ queueDeq_1[2])
        queueCount_2_1 <= queueCount_2_1 + counterUpdate_10;
      if (queueEnq_1[3] ^ queueDeq_1[3])
        queueCount_3_1 <= queueCount_3_1 + counterUpdate_11;
      if (queueEnq_1[4] ^ queueDeq_1[4])
        queueCount_4_1 <= queueCount_4_1 + counterUpdate_12;
      if (queueEnq_1[5] ^ queueDeq_1[5])
        queueCount_5_1 <= queueCount_5_1 + counterUpdate_13;
      if (queueEnq_1[6] ^ queueDeq_1[6])
        queueCount_6_1 <= queueCount_6_1 + counterUpdate_14;
      if (queueEnq_1[7] ^ queueDeq_1[7])
        queueCount_7_1 <= queueCount_7_1 + counterUpdate_15;
      if (queueEnq_2[0] ^ queueDeq_2[0])
        queueCount_0_2 <= queueCount_0_2 + counterUpdate_16;
      if (queueEnq_2[1] ^ queueDeq_2[1])
        queueCount_1_2 <= queueCount_1_2 + counterUpdate_17;
      if (queueEnq_2[2] ^ queueDeq_2[2])
        queueCount_2_2 <= queueCount_2_2 + counterUpdate_18;
      if (queueEnq_2[3] ^ queueDeq_2[3])
        queueCount_3_2 <= queueCount_3_2 + counterUpdate_19;
      if (queueEnq_2[4] ^ queueDeq_2[4])
        queueCount_4_2 <= queueCount_4_2 + counterUpdate_20;
      if (queueEnq_2[5] ^ queueDeq_2[5])
        queueCount_5_2 <= queueCount_5_2 + counterUpdate_21;
      if (queueEnq_2[6] ^ queueDeq_2[6])
        queueCount_6_2 <= queueCount_6_2 + counterUpdate_22;
      if (queueEnq_2[7] ^ queueDeq_2[7])
        queueCount_7_2 <= queueCount_7_2 + counterUpdate_23;
      if (queueEnq_3[0] ^ queueDeq_3[0])
        queueCount_0_3 <= queueCount_0_3 + counterUpdate_24;
      if (queueEnq_3[1] ^ queueDeq_3[1])
        queueCount_1_3 <= queueCount_1_3 + counterUpdate_25;
      if (queueEnq_3[2] ^ queueDeq_3[2])
        queueCount_2_3 <= queueCount_2_3 + counterUpdate_26;
      if (queueEnq_3[3] ^ queueDeq_3[3])
        queueCount_3_3 <= queueCount_3_3 + counterUpdate_27;
      if (queueEnq_3[4] ^ queueDeq_3[4])
        queueCount_4_3 <= queueCount_4_3 + counterUpdate_28;
      if (queueEnq_3[5] ^ queueDeq_3[5])
        queueCount_5_3 <= queueCount_5_3 + counterUpdate_29;
      if (queueEnq_3[6] ^ queueDeq_3[6])
        queueCount_6_3 <= queueCount_6_3 + counterUpdate_30;
      if (queueEnq_3[7] ^ queueDeq_3[7])
        queueCount_7_3 <= queueCount_7_3 + counterUpdate_31;
    end
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:262];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [8:0] i = 9'h0; i < 9'h107; i += 9'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        v0_0 = _RANDOM[9'h0];
        v0_1 = _RANDOM[9'h1];
        v0_2 = _RANDOM[9'h2];
        v0_3 = _RANDOM[9'h3];
        v0_4 = _RANDOM[9'h4];
        v0_5 = _RANDOM[9'h5];
        v0_6 = _RANDOM[9'h6];
        v0_7 = _RANDOM[9'h7];
        v0_8 = _RANDOM[9'h8];
        v0_9 = _RANDOM[9'h9];
        v0_10 = _RANDOM[9'hA];
        v0_11 = _RANDOM[9'hB];
        v0_12 = _RANDOM[9'hC];
        v0_13 = _RANDOM[9'hD];
        v0_14 = _RANDOM[9'hE];
        v0_15 = _RANDOM[9'hF];
        v0_16 = _RANDOM[9'h10];
        v0_17 = _RANDOM[9'h11];
        v0_18 = _RANDOM[9'h12];
        v0_19 = _RANDOM[9'h13];
        v0_20 = _RANDOM[9'h14];
        v0_21 = _RANDOM[9'h15];
        v0_22 = _RANDOM[9'h16];
        v0_23 = _RANDOM[9'h17];
        v0_24 = _RANDOM[9'h18];
        v0_25 = _RANDOM[9'h19];
        v0_26 = _RANDOM[9'h1A];
        v0_27 = _RANDOM[9'h1B];
        v0_28 = _RANDOM[9'h1C];
        v0_29 = _RANDOM[9'h1D];
        v0_30 = _RANDOM[9'h1E];
        v0_31 = _RANDOM[9'h1F];
        v0_32 = _RANDOM[9'h20];
        v0_33 = _RANDOM[9'h21];
        v0_34 = _RANDOM[9'h22];
        v0_35 = _RANDOM[9'h23];
        v0_36 = _RANDOM[9'h24];
        v0_37 = _RANDOM[9'h25];
        v0_38 = _RANDOM[9'h26];
        v0_39 = _RANDOM[9'h27];
        v0_40 = _RANDOM[9'h28];
        v0_41 = _RANDOM[9'h29];
        v0_42 = _RANDOM[9'h2A];
        v0_43 = _RANDOM[9'h2B];
        v0_44 = _RANDOM[9'h2C];
        v0_45 = _RANDOM[9'h2D];
        v0_46 = _RANDOM[9'h2E];
        v0_47 = _RANDOM[9'h2F];
        v0_48 = _RANDOM[9'h30];
        v0_49 = _RANDOM[9'h31];
        v0_50 = _RANDOM[9'h32];
        v0_51 = _RANDOM[9'h33];
        v0_52 = _RANDOM[9'h34];
        v0_53 = _RANDOM[9'h35];
        v0_54 = _RANDOM[9'h36];
        v0_55 = _RANDOM[9'h37];
        v0_56 = _RANDOM[9'h38];
        v0_57 = _RANDOM[9'h39];
        v0_58 = _RANDOM[9'h3A];
        v0_59 = _RANDOM[9'h3B];
        v0_60 = _RANDOM[9'h3C];
        v0_61 = _RANDOM[9'h3D];
        v0_62 = _RANDOM[9'h3E];
        v0_63 = _RANDOM[9'h3F];
        v0_64 = _RANDOM[9'h40];
        v0_65 = _RANDOM[9'h41];
        v0_66 = _RANDOM[9'h42];
        v0_67 = _RANDOM[9'h43];
        v0_68 = _RANDOM[9'h44];
        v0_69 = _RANDOM[9'h45];
        v0_70 = _RANDOM[9'h46];
        v0_71 = _RANDOM[9'h47];
        v0_72 = _RANDOM[9'h48];
        v0_73 = _RANDOM[9'h49];
        v0_74 = _RANDOM[9'h4A];
        v0_75 = _RANDOM[9'h4B];
        v0_76 = _RANDOM[9'h4C];
        v0_77 = _RANDOM[9'h4D];
        v0_78 = _RANDOM[9'h4E];
        v0_79 = _RANDOM[9'h4F];
        v0_80 = _RANDOM[9'h50];
        v0_81 = _RANDOM[9'h51];
        v0_82 = _RANDOM[9'h52];
        v0_83 = _RANDOM[9'h53];
        v0_84 = _RANDOM[9'h54];
        v0_85 = _RANDOM[9'h55];
        v0_86 = _RANDOM[9'h56];
        v0_87 = _RANDOM[9'h57];
        v0_88 = _RANDOM[9'h58];
        v0_89 = _RANDOM[9'h59];
        v0_90 = _RANDOM[9'h5A];
        v0_91 = _RANDOM[9'h5B];
        v0_92 = _RANDOM[9'h5C];
        v0_93 = _RANDOM[9'h5D];
        v0_94 = _RANDOM[9'h5E];
        v0_95 = _RANDOM[9'h5F];
        v0_96 = _RANDOM[9'h60];
        v0_97 = _RANDOM[9'h61];
        v0_98 = _RANDOM[9'h62];
        v0_99 = _RANDOM[9'h63];
        v0_100 = _RANDOM[9'h64];
        v0_101 = _RANDOM[9'h65];
        v0_102 = _RANDOM[9'h66];
        v0_103 = _RANDOM[9'h67];
        v0_104 = _RANDOM[9'h68];
        v0_105 = _RANDOM[9'h69];
        v0_106 = _RANDOM[9'h6A];
        v0_107 = _RANDOM[9'h6B];
        v0_108 = _RANDOM[9'h6C];
        v0_109 = _RANDOM[9'h6D];
        v0_110 = _RANDOM[9'h6E];
        v0_111 = _RANDOM[9'h6F];
        v0_112 = _RANDOM[9'h70];
        v0_113 = _RANDOM[9'h71];
        v0_114 = _RANDOM[9'h72];
        v0_115 = _RANDOM[9'h73];
        v0_116 = _RANDOM[9'h74];
        v0_117 = _RANDOM[9'h75];
        v0_118 = _RANDOM[9'h76];
        v0_119 = _RANDOM[9'h77];
        v0_120 = _RANDOM[9'h78];
        v0_121 = _RANDOM[9'h79];
        v0_122 = _RANDOM[9'h7A];
        v0_123 = _RANDOM[9'h7B];
        v0_124 = _RANDOM[9'h7C];
        v0_125 = _RANDOM[9'h7D];
        v0_126 = _RANDOM[9'h7E];
        v0_127 = _RANDOM[9'h7F];
        v0_128 = _RANDOM[9'h80];
        v0_129 = _RANDOM[9'h81];
        v0_130 = _RANDOM[9'h82];
        v0_131 = _RANDOM[9'h83];
        v0_132 = _RANDOM[9'h84];
        v0_133 = _RANDOM[9'h85];
        v0_134 = _RANDOM[9'h86];
        v0_135 = _RANDOM[9'h87];
        v0_136 = _RANDOM[9'h88];
        v0_137 = _RANDOM[9'h89];
        v0_138 = _RANDOM[9'h8A];
        v0_139 = _RANDOM[9'h8B];
        v0_140 = _RANDOM[9'h8C];
        v0_141 = _RANDOM[9'h8D];
        v0_142 = _RANDOM[9'h8E];
        v0_143 = _RANDOM[9'h8F];
        v0_144 = _RANDOM[9'h90];
        v0_145 = _RANDOM[9'h91];
        v0_146 = _RANDOM[9'h92];
        v0_147 = _RANDOM[9'h93];
        v0_148 = _RANDOM[9'h94];
        v0_149 = _RANDOM[9'h95];
        v0_150 = _RANDOM[9'h96];
        v0_151 = _RANDOM[9'h97];
        v0_152 = _RANDOM[9'h98];
        v0_153 = _RANDOM[9'h99];
        v0_154 = _RANDOM[9'h9A];
        v0_155 = _RANDOM[9'h9B];
        v0_156 = _RANDOM[9'h9C];
        v0_157 = _RANDOM[9'h9D];
        v0_158 = _RANDOM[9'h9E];
        v0_159 = _RANDOM[9'h9F];
        v0_160 = _RANDOM[9'hA0];
        v0_161 = _RANDOM[9'hA1];
        v0_162 = _RANDOM[9'hA2];
        v0_163 = _RANDOM[9'hA3];
        v0_164 = _RANDOM[9'hA4];
        v0_165 = _RANDOM[9'hA5];
        v0_166 = _RANDOM[9'hA6];
        v0_167 = _RANDOM[9'hA7];
        v0_168 = _RANDOM[9'hA8];
        v0_169 = _RANDOM[9'hA9];
        v0_170 = _RANDOM[9'hAA];
        v0_171 = _RANDOM[9'hAB];
        v0_172 = _RANDOM[9'hAC];
        v0_173 = _RANDOM[9'hAD];
        v0_174 = _RANDOM[9'hAE];
        v0_175 = _RANDOM[9'hAF];
        v0_176 = _RANDOM[9'hB0];
        v0_177 = _RANDOM[9'hB1];
        v0_178 = _RANDOM[9'hB2];
        v0_179 = _RANDOM[9'hB3];
        v0_180 = _RANDOM[9'hB4];
        v0_181 = _RANDOM[9'hB5];
        v0_182 = _RANDOM[9'hB6];
        v0_183 = _RANDOM[9'hB7];
        v0_184 = _RANDOM[9'hB8];
        v0_185 = _RANDOM[9'hB9];
        v0_186 = _RANDOM[9'hBA];
        v0_187 = _RANDOM[9'hBB];
        v0_188 = _RANDOM[9'hBC];
        v0_189 = _RANDOM[9'hBD];
        v0_190 = _RANDOM[9'hBE];
        v0_191 = _RANDOM[9'hBF];
        v0_192 = _RANDOM[9'hC0];
        v0_193 = _RANDOM[9'hC1];
        v0_194 = _RANDOM[9'hC2];
        v0_195 = _RANDOM[9'hC3];
        v0_196 = _RANDOM[9'hC4];
        v0_197 = _RANDOM[9'hC5];
        v0_198 = _RANDOM[9'hC6];
        v0_199 = _RANDOM[9'hC7];
        v0_200 = _RANDOM[9'hC8];
        v0_201 = _RANDOM[9'hC9];
        v0_202 = _RANDOM[9'hCA];
        v0_203 = _RANDOM[9'hCB];
        v0_204 = _RANDOM[9'hCC];
        v0_205 = _RANDOM[9'hCD];
        v0_206 = _RANDOM[9'hCE];
        v0_207 = _RANDOM[9'hCF];
        v0_208 = _RANDOM[9'hD0];
        v0_209 = _RANDOM[9'hD1];
        v0_210 = _RANDOM[9'hD2];
        v0_211 = _RANDOM[9'hD3];
        v0_212 = _RANDOM[9'hD4];
        v0_213 = _RANDOM[9'hD5];
        v0_214 = _RANDOM[9'hD6];
        v0_215 = _RANDOM[9'hD7];
        v0_216 = _RANDOM[9'hD8];
        v0_217 = _RANDOM[9'hD9];
        v0_218 = _RANDOM[9'hDA];
        v0_219 = _RANDOM[9'hDB];
        v0_220 = _RANDOM[9'hDC];
        v0_221 = _RANDOM[9'hDD];
        v0_222 = _RANDOM[9'hDE];
        v0_223 = _RANDOM[9'hDF];
        v0_224 = _RANDOM[9'hE0];
        v0_225 = _RANDOM[9'hE1];
        v0_226 = _RANDOM[9'hE2];
        v0_227 = _RANDOM[9'hE3];
        v0_228 = _RANDOM[9'hE4];
        v0_229 = _RANDOM[9'hE5];
        v0_230 = _RANDOM[9'hE6];
        v0_231 = _RANDOM[9'hE7];
        v0_232 = _RANDOM[9'hE8];
        v0_233 = _RANDOM[9'hE9];
        v0_234 = _RANDOM[9'hEA];
        v0_235 = _RANDOM[9'hEB];
        v0_236 = _RANDOM[9'hEC];
        v0_237 = _RANDOM[9'hED];
        v0_238 = _RANDOM[9'hEE];
        v0_239 = _RANDOM[9'hEF];
        v0_240 = _RANDOM[9'hF0];
        v0_241 = _RANDOM[9'hF1];
        v0_242 = _RANDOM[9'hF2];
        v0_243 = _RANDOM[9'hF3];
        v0_244 = _RANDOM[9'hF4];
        v0_245 = _RANDOM[9'hF5];
        v0_246 = _RANDOM[9'hF6];
        v0_247 = _RANDOM[9'hF7];
        v0_248 = _RANDOM[9'hF8];
        v0_249 = _RANDOM[9'hF9];
        v0_250 = _RANDOM[9'hFA];
        v0_251 = _RANDOM[9'hFB];
        v0_252 = _RANDOM[9'hFC];
        v0_253 = _RANDOM[9'hFD];
        v0_254 = _RANDOM[9'hFE];
        v0_255 = _RANDOM[9'hFF];
        queueCount_0 = _RANDOM[9'h100][6:0];
        queueCount_1 = _RANDOM[9'h100][13:7];
        queueCount_2 = _RANDOM[9'h100][20:14];
        queueCount_3 = _RANDOM[9'h100][27:21];
        queueCount_4 = {_RANDOM[9'h100][31:28], _RANDOM[9'h101][2:0]};
        queueCount_5 = _RANDOM[9'h101][9:3];
        queueCount_6 = _RANDOM[9'h101][16:10];
        queueCount_7 = _RANDOM[9'h101][23:17];
        queueCount_0_1 = _RANDOM[9'h101][30:24];
        queueCount_1_1 = {_RANDOM[9'h101][31], _RANDOM[9'h102][5:0]};
        queueCount_2_1 = _RANDOM[9'h102][12:6];
        queueCount_3_1 = _RANDOM[9'h102][19:13];
        queueCount_4_1 = _RANDOM[9'h102][26:20];
        queueCount_5_1 = {_RANDOM[9'h102][31:27], _RANDOM[9'h103][1:0]};
        queueCount_6_1 = _RANDOM[9'h103][8:2];
        queueCount_7_1 = _RANDOM[9'h103][15:9];
        queueCount_0_2 = _RANDOM[9'h103][22:16];
        queueCount_1_2 = _RANDOM[9'h103][29:23];
        queueCount_2_2 = {_RANDOM[9'h103][31:30], _RANDOM[9'h104][4:0]};
        queueCount_3_2 = _RANDOM[9'h104][11:5];
        queueCount_4_2 = _RANDOM[9'h104][18:12];
        queueCount_5_2 = _RANDOM[9'h104][25:19];
        queueCount_6_2 = {_RANDOM[9'h104][31:26], _RANDOM[9'h105][0]};
        queueCount_7_2 = _RANDOM[9'h105][7:1];
        queueCount_0_3 = _RANDOM[9'h105][14:8];
        queueCount_1_3 = _RANDOM[9'h105][21:15];
        queueCount_2_3 = _RANDOM[9'h105][28:22];
        queueCount_3_3 = {_RANDOM[9'h105][31:29], _RANDOM[9'h106][3:0]};
        queueCount_4_3 = _RANDOM[9'h106][10:4];
        queueCount_5_3 = _RANDOM[9'h106][17:11];
        queueCount_6_3 = _RANDOM[9'h106][24:18];
        queueCount_7_3 = _RANDOM[9'h106][31:25];
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  wire [9:0]         sourceQueue_deq_bits;
  wire [31:0]        axi4Port_aw_bits_addr_0;
  assign axi4Port_aw_bits_addr_0 = _storeUnit_memRequest_bits_address;
  assign dataQueue_enq_bits_index = _storeUnit_memRequest_bits_index;
  assign dataQueue_enq_bits_address = _storeUnit_memRequest_bits_address;
  wire [6:0]         simpleSourceQueue_deq_bits;
  wire [31:0]        simpleAccessPorts_aw_bits_addr_0;
  assign simpleAccessPorts_aw_bits_addr_0 = _otherUnit_memWriteRequest_bits_address;
  wire [3:0]         otherUnitTargetQueue_enq_bits;
  assign otherUnitTargetQueue_enq_bits = _otherUnit_status_targetLane;
  assign simpleDataQueue_enq_bits_source = _otherUnit_memWriteRequest_bits_source;
  assign simpleDataQueue_enq_bits_address = _otherUnit_memWriteRequest_bits_address;
  assign simpleDataQueue_enq_bits_size = _otherUnit_memWriteRequest_bits_size;
  wire               writeQueueVec_0_empty;
  assign writeQueueVec_0_empty = _writeQueueVec_fifo_empty;
  wire               writeQueueVec_0_full;
  assign writeQueueVec_0_full = _writeQueueVec_fifo_full;
  wire               writeQueueVec_1_empty;
  assign writeQueueVec_1_empty = _writeQueueVec_fifo_1_empty;
  wire               writeQueueVec_1_full;
  assign writeQueueVec_1_full = _writeQueueVec_fifo_1_full;
  wire               writeQueueVec_2_empty;
  assign writeQueueVec_2_empty = _writeQueueVec_fifo_2_empty;
  wire               writeQueueVec_2_full;
  assign writeQueueVec_2_full = _writeQueueVec_fifo_2_full;
  wire               writeQueueVec_3_empty;
  assign writeQueueVec_3_empty = _writeQueueVec_fifo_3_empty;
  wire               writeQueueVec_3_full;
  assign writeQueueVec_3_full = _writeQueueVec_fifo_3_full;
  assign otherUnitTargetQueue_empty = _otherUnitTargetQueue_fifo_empty;
  wire               otherUnitTargetQueue_full;
  assign otherUnitTargetQueue_full = _otherUnitTargetQueue_fifo_full;
  wire               otherUnitDataQueueVec_0_empty;
  assign otherUnitDataQueueVec_0_empty = _otherUnitDataQueueVec_fifo_empty;
  wire               otherUnitDataQueueVec_0_full;
  assign otherUnitDataQueueVec_0_full = _otherUnitDataQueueVec_fifo_full;
  wire               otherUnitDataQueueVec_1_empty;
  assign otherUnitDataQueueVec_1_empty = _otherUnitDataQueueVec_fifo_1_empty;
  wire               otherUnitDataQueueVec_1_full;
  assign otherUnitDataQueueVec_1_full = _otherUnitDataQueueVec_fifo_1_full;
  wire               otherUnitDataQueueVec_2_empty;
  assign otherUnitDataQueueVec_2_empty = _otherUnitDataQueueVec_fifo_2_empty;
  wire               otherUnitDataQueueVec_2_full;
  assign otherUnitDataQueueVec_2_full = _otherUnitDataQueueVec_fifo_2_full;
  wire               otherUnitDataQueueVec_3_empty;
  assign otherUnitDataQueueVec_3_empty = _otherUnitDataQueueVec_fifo_3_empty;
  wire               otherUnitDataQueueVec_3_full;
  assign otherUnitDataQueueVec_3_full = _otherUnitDataQueueVec_fifo_3_full;
  wire               writeIndexQueue_empty;
  assign writeIndexQueue_empty = _writeIndexQueue_fifo_empty;
  wire               writeIndexQueue_full;
  assign writeIndexQueue_full = _writeIndexQueue_fifo_full;
  wire               writeIndexQueue_1_empty;
  assign writeIndexQueue_1_empty = _writeIndexQueue_fifo_1_empty;
  wire               writeIndexQueue_1_full;
  assign writeIndexQueue_1_full = _writeIndexQueue_fifo_1_full;
  wire               writeIndexQueue_2_empty;
  assign writeIndexQueue_2_empty = _writeIndexQueue_fifo_2_empty;
  wire               writeIndexQueue_2_full;
  assign writeIndexQueue_2_full = _writeIndexQueue_fifo_2_full;
  wire               writeIndexQueue_3_empty;
  assign writeIndexQueue_3_empty = _writeIndexQueue_fifo_3_empty;
  wire               writeIndexQueue_3_full;
  assign writeIndexQueue_3_full = _writeIndexQueue_fifo_3_full;
  wire               sourceQueue_empty;
  assign sourceQueue_empty = _sourceQueue_fifo_empty;
  wire               sourceQueue_full;
  assign sourceQueue_full = _sourceQueue_fifo_full;
  wire               dataQueue_empty;
  assign dataQueue_empty = _dataQueue_fifo_empty;
  wire               dataQueue_full;
  assign dataQueue_full = _dataQueue_fifo_full;
  wire               simpleSourceQueue_empty;
  assign simpleSourceQueue_empty = _simpleSourceQueue_fifo_empty;
  wire               simpleSourceQueue_full;
  assign simpleSourceQueue_full = _simpleSourceQueue_fifo_full;
  wire               simpleDataQueue_empty;
  assign simpleDataQueue_empty = _simpleDataQueue_fifo_empty;
  wire               simpleDataQueue_full;
  assign simpleDataQueue_full = _simpleDataQueue_fifo_full;
  LoadUnit loadUnit (
    .clock                                                  (clock),
    .reset                                                  (reset),
    .lsuRequest_valid                                       (reqEnq_0),
    .lsuRequest_bits_instructionInformation_nf              (request_bits_instructionInformation_nf_0),
    .lsuRequest_bits_instructionInformation_mew             (request_bits_instructionInformation_mew_0),
    .lsuRequest_bits_instructionInformation_mop             (request_bits_instructionInformation_mop_0),
    .lsuRequest_bits_instructionInformation_lumop           (request_bits_instructionInformation_lumop_0),
    .lsuRequest_bits_instructionInformation_eew             (request_bits_instructionInformation_eew_0),
    .lsuRequest_bits_instructionInformation_vs3             (request_bits_instructionInformation_vs3_0),
    .lsuRequest_bits_instructionInformation_isStore         (request_bits_instructionInformation_isStore_0),
    .lsuRequest_bits_instructionInformation_maskedLoadStore (request_bits_instructionInformation_maskedLoadStore_0),
    .lsuRequest_bits_rs1Data                                (request_bits_rs1Data_0),
    .lsuRequest_bits_rs2Data                                (request_bits_rs2Data_0),
    .lsuRequest_bits_instructionIndex                       (request_bits_instructionIndex_0),
    .csrInterface_vl                                        (csrInterface_vl),
    .csrInterface_vStart                                    (csrInterface_vStart),
    .csrInterface_vlmul                                     (csrInterface_vlmul),
    .csrInterface_vSew                                      (csrInterface_vSew),
    .csrInterface_vxrm                                      (csrInterface_vxrm),
    .csrInterface_vta                                       (csrInterface_vta),
    .csrInterface_vma                                       (csrInterface_vma),
    .maskInput                                              (_GEN_127[maskSelect]),
    .maskSelect_valid                                       (_loadUnit_maskSelect_valid),
    .maskSelect_bits                                        (_loadUnit_maskSelect_bits),
    .addressConflict                                        (stallLoad),
    .memRequest_ready                                       (sourceQueue_enq_ready & axi4Port_ar_ready_0),
    .memRequest_valid                                       (_loadUnit_memRequest_valid),
    .memRequest_bits_src                                    (sourceQueue_enq_bits),
    .memRequest_bits_address                                (axi4Port_ar_bits_addr_0),
    .memResponse_ready                                      (axi4Port_r_ready_0),
    .memResponse_valid                                      (axi4Port_r_valid_0),
    .memResponse_bits_data                                  (axi4Port_r_bits_data_0),
    .memResponse_bits_index                                 (sourceQueue_deq_bits),
    .status_idle                                            (_loadUnit_status_idle),
    .status_last                                            (_loadUnit_status_last),
    .status_instructionIndex                                (_loadUnit_status_instructionIndex),
    .status_changeMaskGroup                                 (/* unused */),
    .status_startAddress                                    (_loadUnit_status_startAddress),
    .status_endAddress                                      (_loadUnit_status_endAddress),
    .vrfWritePort_0_ready                                   (writeQueueVec_0_enq_ready & ~(otherTryToWrite[0])),
    .vrfWritePort_0_valid                                   (_loadUnit_vrfWritePort_0_valid),
    .vrfWritePort_0_bits_vd                                 (_loadUnit_vrfWritePort_0_bits_vd),
    .vrfWritePort_0_bits_offset                             (_loadUnit_vrfWritePort_0_bits_offset),
    .vrfWritePort_0_bits_mask                               (_loadUnit_vrfWritePort_0_bits_mask),
    .vrfWritePort_0_bits_data                               (_loadUnit_vrfWritePort_0_bits_data),
    .vrfWritePort_0_bits_instructionIndex                   (_loadUnit_vrfWritePort_0_bits_instructionIndex),
    .vrfWritePort_1_ready                                   (writeQueueVec_1_enq_ready & ~(otherTryToWrite[1])),
    .vrfWritePort_1_valid                                   (_loadUnit_vrfWritePort_1_valid),
    .vrfWritePort_1_bits_vd                                 (_loadUnit_vrfWritePort_1_bits_vd),
    .vrfWritePort_1_bits_offset                             (_loadUnit_vrfWritePort_1_bits_offset),
    .vrfWritePort_1_bits_mask                               (_loadUnit_vrfWritePort_1_bits_mask),
    .vrfWritePort_1_bits_data                               (_loadUnit_vrfWritePort_1_bits_data),
    .vrfWritePort_1_bits_instructionIndex                   (_loadUnit_vrfWritePort_1_bits_instructionIndex),
    .vrfWritePort_2_ready                                   (writeQueueVec_2_enq_ready & ~(otherTryToWrite[2])),
    .vrfWritePort_2_valid                                   (_loadUnit_vrfWritePort_2_valid),
    .vrfWritePort_2_bits_vd                                 (_loadUnit_vrfWritePort_2_bits_vd),
    .vrfWritePort_2_bits_offset                             (_loadUnit_vrfWritePort_2_bits_offset),
    .vrfWritePort_2_bits_mask                               (_loadUnit_vrfWritePort_2_bits_mask),
    .vrfWritePort_2_bits_data                               (_loadUnit_vrfWritePort_2_bits_data),
    .vrfWritePort_2_bits_instructionIndex                   (_loadUnit_vrfWritePort_2_bits_instructionIndex),
    .vrfWritePort_3_ready                                   (writeQueueVec_3_enq_ready & ~(otherTryToWrite[3])),
    .vrfWritePort_3_valid                                   (_loadUnit_vrfWritePort_3_valid),
    .vrfWritePort_3_bits_vd                                 (_loadUnit_vrfWritePort_3_bits_vd),
    .vrfWritePort_3_bits_offset                             (_loadUnit_vrfWritePort_3_bits_offset),
    .vrfWritePort_3_bits_mask                               (_loadUnit_vrfWritePort_3_bits_mask),
    .vrfWritePort_3_bits_data                               (_loadUnit_vrfWritePort_3_bits_data),
    .vrfWritePort_3_bits_instructionIndex                   (_loadUnit_vrfWritePort_3_bits_instructionIndex)
  );
  StoreUnit storeUnit (
    .clock                                                  (clock),
    .reset                                                  (reset),
    .lsuRequest_valid                                       (reqEnq_1),
    .lsuRequest_bits_instructionInformation_nf              (request_bits_instructionInformation_nf_0),
    .lsuRequest_bits_instructionInformation_mew             (request_bits_instructionInformation_mew_0),
    .lsuRequest_bits_instructionInformation_mop             (request_bits_instructionInformation_mop_0),
    .lsuRequest_bits_instructionInformation_lumop           (request_bits_instructionInformation_lumop_0),
    .lsuRequest_bits_instructionInformation_eew             (request_bits_instructionInformation_eew_0),
    .lsuRequest_bits_instructionInformation_vs3             (request_bits_instructionInformation_vs3_0),
    .lsuRequest_bits_instructionInformation_isStore         (request_bits_instructionInformation_isStore_0),
    .lsuRequest_bits_instructionInformation_maskedLoadStore (request_bits_instructionInformation_maskedLoadStore_0),
    .lsuRequest_bits_rs1Data                                (request_bits_rs1Data_0),
    .lsuRequest_bits_rs2Data                                (request_bits_rs2Data_0),
    .lsuRequest_bits_instructionIndex                       (request_bits_instructionIndex_0),
    .csrInterface_vl                                        (csrInterface_vl),
    .csrInterface_vStart                                    (csrInterface_vStart),
    .csrInterface_vlmul                                     (csrInterface_vlmul),
    .csrInterface_vSew                                      (csrInterface_vSew),
    .csrInterface_vxrm                                      (csrInterface_vxrm),
    .csrInterface_vta                                       (csrInterface_vta),
    .csrInterface_vma                                       (csrInterface_vma),
    .maskInput                                              (_GEN_128[maskSelect_1]),
    .maskSelect_valid                                       (_storeUnit_maskSelect_valid),
    .maskSelect_bits                                        (_storeUnit_maskSelect_bits),
    .memRequest_ready                                       (axi4Port_aw_ready_0 & dataQueue_enq_ready),
    .memRequest_valid                                       (_storeUnit_memRequest_valid),
    .memRequest_bits_data                                   (dataQueue_enq_bits_data),
    .memRequest_bits_mask                                   (dataQueue_enq_bits_mask),
    .memRequest_bits_index                                  (_storeUnit_memRequest_bits_index),
    .memRequest_bits_address                                (_storeUnit_memRequest_bits_address),
    .status_idle                                            (_storeUnit_status_idle),
    .status_last                                            (_storeUnit_status_last),
    .status_instructionIndex                                (_storeUnit_status_instructionIndex),
    .status_changeMaskGroup                                 (/* unused */),
    .status_startAddress                                    (_storeUnit_status_startAddress),
    .status_endAddress                                      (_storeUnit_status_endAddress),
    .vrfReadDataPorts_0_ready                               (vrfReadDataPorts_0_ready_0 & ~(otherTryReadVrf[0])),
    .vrfReadDataPorts_0_valid                               (_storeUnit_vrfReadDataPorts_0_valid),
    .vrfReadDataPorts_0_bits_vs                             (_storeUnit_vrfReadDataPorts_0_bits_vs),
    .vrfReadDataPorts_0_bits_offset                         (_storeUnit_vrfReadDataPorts_0_bits_offset),
    .vrfReadDataPorts_0_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_0_bits_instructionIndex),
    .vrfReadDataPorts_1_ready                               (vrfReadDataPorts_1_ready_0 & ~(otherTryReadVrf[1])),
    .vrfReadDataPorts_1_valid                               (_storeUnit_vrfReadDataPorts_1_valid),
    .vrfReadDataPorts_1_bits_vs                             (_storeUnit_vrfReadDataPorts_1_bits_vs),
    .vrfReadDataPorts_1_bits_offset                         (_storeUnit_vrfReadDataPorts_1_bits_offset),
    .vrfReadDataPorts_1_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_1_bits_instructionIndex),
    .vrfReadDataPorts_2_ready                               (vrfReadDataPorts_2_ready_0 & ~(otherTryReadVrf[2])),
    .vrfReadDataPorts_2_valid                               (_storeUnit_vrfReadDataPorts_2_valid),
    .vrfReadDataPorts_2_bits_vs                             (_storeUnit_vrfReadDataPorts_2_bits_vs),
    .vrfReadDataPorts_2_bits_offset                         (_storeUnit_vrfReadDataPorts_2_bits_offset),
    .vrfReadDataPorts_2_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_2_bits_instructionIndex),
    .vrfReadDataPorts_3_ready                               (vrfReadDataPorts_3_ready_0 & ~(otherTryReadVrf[3])),
    .vrfReadDataPorts_3_valid                               (_storeUnit_vrfReadDataPorts_3_valid),
    .vrfReadDataPorts_3_bits_vs                             (_storeUnit_vrfReadDataPorts_3_bits_vs),
    .vrfReadDataPorts_3_bits_offset                         (_storeUnit_vrfReadDataPorts_3_bits_offset),
    .vrfReadDataPorts_3_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_3_bits_instructionIndex),
    .vrfReadResults_0_valid                                 (vrfReadResults_0_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_0_bits                                  (vrfReadResults_0_bits),
    .vrfReadResults_1_valid                                 (vrfReadResults_1_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_1_bits                                  (vrfReadResults_1_bits),
    .vrfReadResults_2_valid                                 (vrfReadResults_2_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_2_bits                                  (vrfReadResults_2_bits),
    .vrfReadResults_3_valid                                 (vrfReadResults_3_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_3_bits                                  (vrfReadResults_3_bits),
    .storeResponse                                          (axi4Port_b_valid_0)
  );
  SimpleAccessUnit otherUnit (
    .clock                                                  (clock),
    .reset                                                  (reset),
    .lsuRequest_valid                                       (reqEnq_2),
    .lsuRequest_bits_instructionInformation_nf              (request_bits_instructionInformation_nf_0),
    .lsuRequest_bits_instructionInformation_mew             (request_bits_instructionInformation_mew_0),
    .lsuRequest_bits_instructionInformation_mop             (request_bits_instructionInformation_mop_0),
    .lsuRequest_bits_instructionInformation_lumop           (request_bits_instructionInformation_lumop_0),
    .lsuRequest_bits_instructionInformation_eew             (request_bits_instructionInformation_eew_0),
    .lsuRequest_bits_instructionInformation_vs3             (request_bits_instructionInformation_vs3_0),
    .lsuRequest_bits_instructionInformation_isStore         (request_bits_instructionInformation_isStore_0),
    .lsuRequest_bits_instructionInformation_maskedLoadStore (request_bits_instructionInformation_maskedLoadStore_0),
    .lsuRequest_bits_rs1Data                                (request_bits_rs1Data_0),
    .lsuRequest_bits_rs2Data                                (request_bits_rs2Data_0),
    .lsuRequest_bits_instructionIndex                       (request_bits_instructionIndex_0),
    .vrfReadDataPorts_ready                                 (otherUnit_vrfReadDataPorts_ready),
    .vrfReadDataPorts_valid                                 (_otherUnit_vrfReadDataPorts_valid),
    .vrfReadDataPorts_bits_vs                               (_otherUnit_vrfReadDataPorts_bits_vs),
    .vrfReadDataPorts_bits_offset                           (_otherUnit_vrfReadDataPorts_bits_offset),
    .vrfReadDataPorts_bits_instructionIndex                 (_otherUnit_vrfReadDataPorts_bits_instructionIndex),
    .vrfReadResults_valid                                   (otherUnitTargetQueue_deq_ready),
    .vrfReadResults_bits
      ((otherUnitTargetQueue_deq_bits[0] ? otherUnitDataQueueVec_0_deq_bits : 32'h0) | (otherUnitTargetQueue_deq_bits[1] ? otherUnitDataQueueVec_1_deq_bits : 32'h0)
       | (otherUnitTargetQueue_deq_bits[2] ? otherUnitDataQueueVec_2_deq_bits : 32'h0) | (otherUnitTargetQueue_deq_bits[3] ? otherUnitDataQueueVec_3_deq_bits : 32'h0)),
    .offsetReadResult_0_valid                               (offsetReadResult_0_valid),
    .offsetReadResult_0_bits                                (offsetReadResult_0_bits),
    .offsetReadResult_1_valid                               (offsetReadResult_1_valid),
    .offsetReadResult_1_bits                                (offsetReadResult_1_bits),
    .offsetReadResult_2_valid                               (offsetReadResult_2_valid),
    .offsetReadResult_2_bits                                (offsetReadResult_2_bits),
    .offsetReadResult_3_valid                               (offsetReadResult_3_valid),
    .offsetReadResult_3_bits                                (offsetReadResult_3_bits),
    .maskInput                                              (_GEN_129[maskSelect_2]),
    .maskSelect_valid                                       (_otherUnit_maskSelect_valid),
    .maskSelect_bits                                        (_otherUnit_maskSelect_bits),
    .memReadRequest_ready                                   (simpleSourceQueue_enq_ready & simpleAccessPorts_ar_ready_0),
    .memReadRequest_valid                                   (_otherUnit_memReadRequest_valid),
    .memReadRequest_bits_address                            (simpleAccessPorts_ar_bits_addr_0),
    .memReadRequest_bits_source                             (simpleSourceQueue_enq_bits),
    .memReadResponse_ready                                  (simpleAccessPorts_r_ready_0),
    .memReadResponse_valid                                  (simpleAccessPorts_r_valid_0),
    .memReadResponse_bits_data                              (simpleAccessPorts_r_bits_data_0),
    .memReadResponse_bits_source                            (simpleSourceQueue_deq_bits),
    .memWriteRequest_ready                                  (simpleAccessPorts_aw_ready_0 & simpleDataQueue_enq_ready),
    .memWriteRequest_valid                                  (_otherUnit_memWriteRequest_valid),
    .memWriteRequest_bits_data                              (simpleDataQueue_enq_bits_data),
    .memWriteRequest_bits_mask                              (simpleDataQueue_enq_bits_mask),
    .memWriteRequest_bits_source                            (_otherUnit_memWriteRequest_bits_source),
    .memWriteRequest_bits_address                           (_otherUnit_memWriteRequest_bits_address),
    .memWriteRequest_bits_size                              (_otherUnit_memWriteRequest_bits_size),
    .vrfWritePort_ready                                     (|(_otherUnit_status_targetLane & {otherUnit_vrfWritePort_ready_hi, otherUnit_vrfWritePort_ready_lo})),
    .vrfWritePort_valid                                     (_otherUnit_vrfWritePort_valid),
    .vrfWritePort_bits_vd                                   (_otherUnit_vrfWritePort_bits_vd),
    .vrfWritePort_bits_offset                               (_otherUnit_vrfWritePort_bits_offset),
    .vrfWritePort_bits_mask                                 (_otherUnit_vrfWritePort_bits_mask),
    .vrfWritePort_bits_data                                 (_otherUnit_vrfWritePort_bits_data),
    .vrfWritePort_bits_last                                 (_otherUnit_vrfWritePort_bits_last),
    .vrfWritePort_bits_instructionIndex                     (_otherUnit_vrfWritePort_bits_instructionIndex),
    .csrInterface_vl                                        (csrInterface_vl),
    .csrInterface_vStart                                    (csrInterface_vStart),
    .csrInterface_vlmul                                     (csrInterface_vlmul),
    .csrInterface_vSew                                      (csrInterface_vSew),
    .csrInterface_vxrm                                      (csrInterface_vxrm),
    .csrInterface_vta                                       (csrInterface_vta),
    .csrInterface_vma                                       (csrInterface_vma),
    .status_idle                                            (_otherUnit_status_idle),
    .status_last                                            (_otherUnit_status_last),
    .status_instructionIndex                                (_otherUnit_status_instructionIndex),
    .status_targetLane                                      (_otherUnit_status_targetLane),
    .status_isStore                                         (_otherUnit_status_isStore),
    .offsetRelease_0                                        (_otherUnit_offsetRelease_0),
    .offsetRelease_1                                        (_otherUnit_offsetRelease_1),
    .offsetRelease_2                                        (_otherUnit_offsetRelease_2),
    .offsetRelease_3                                        (_otherUnit_offsetRelease_3)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(55)
  ) writeQueueVec_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_0_writeValid_T & ~(_writeQueueVec_fifo_empty & writeQueueVec_0_deq_ready))),
    .pop_req_n    (~(writeQueueVec_0_deq_ready & ~_writeQueueVec_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn),
    .empty        (_writeQueueVec_fifo_empty),
    .almost_empty (writeQueueVec_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_0_almostFull),
    .full         (_writeQueueVec_fifo_full),
    .error        (_writeQueueVec_fifo_error),
    .data_out     (_writeQueueVec_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(55)
  ) writeQueueVec_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_1_writeValid_T & ~(_writeQueueVec_fifo_1_empty & writeQueueVec_1_deq_ready))),
    .pop_req_n    (~(writeQueueVec_1_deq_ready & ~_writeQueueVec_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_1),
    .empty        (_writeQueueVec_fifo_1_empty),
    .almost_empty (writeQueueVec_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_1_almostFull),
    .full         (_writeQueueVec_fifo_1_full),
    .error        (_writeQueueVec_fifo_1_error),
    .data_out     (_writeQueueVec_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(55)
  ) writeQueueVec_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_2_writeValid_T & ~(_writeQueueVec_fifo_2_empty & writeQueueVec_2_deq_ready))),
    .pop_req_n    (~(writeQueueVec_2_deq_ready & ~_writeQueueVec_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_2),
    .empty        (_writeQueueVec_fifo_2_empty),
    .almost_empty (writeQueueVec_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_2_almostFull),
    .full         (_writeQueueVec_fifo_2_full),
    .error        (_writeQueueVec_fifo_2_error),
    .data_out     (_writeQueueVec_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(55)
  ) writeQueueVec_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_3_writeValid_T & ~(_writeQueueVec_fifo_3_empty & writeQueueVec_3_deq_ready))),
    .pop_req_n    (~(writeQueueVec_3_deq_ready & ~_writeQueueVec_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_3),
    .empty        (_writeQueueVec_fifo_3_empty),
    .almost_empty (writeQueueVec_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_3_almostFull),
    .full         (_writeQueueVec_fifo_3_full),
    .error        (_writeQueueVec_fifo_3_error),
    .data_out     (_writeQueueVec_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(4)
  ) otherUnitTargetQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitTargetQueue_enq_ready & otherUnitTargetQueue_enq_valid)),
    .pop_req_n    (~(otherUnitTargetQueue_deq_ready & ~_otherUnitTargetQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitTargetQueue_enq_bits),
    .empty        (_otherUnitTargetQueue_fifo_empty),
    .almost_empty (otherUnitTargetQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitTargetQueue_almostFull),
    .full         (_otherUnitTargetQueue_fifo_full),
    .error        (_otherUnitTargetQueue_fifo_error),
    .data_out     (otherUnitTargetQueue_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_0_enq_ready & otherUnitDataQueueVec_0_enq_valid & ~(_otherUnitDataQueueVec_fifo_empty & otherUnitDataQueueVec_0_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_0_deq_ready & ~_otherUnitDataQueueVec_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_0_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_empty),
    .almost_empty (otherUnitDataQueueVec_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_0_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_full),
    .error        (_otherUnitDataQueueVec_fifo_error),
    .data_out     (_otherUnitDataQueueVec_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_1_enq_ready & otherUnitDataQueueVec_1_enq_valid & ~(_otherUnitDataQueueVec_fifo_1_empty & otherUnitDataQueueVec_1_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_1_deq_ready & ~_otherUnitDataQueueVec_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_1_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_1_empty),
    .almost_empty (otherUnitDataQueueVec_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_1_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_1_full),
    .error        (_otherUnitDataQueueVec_fifo_1_error),
    .data_out     (_otherUnitDataQueueVec_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_2_enq_ready & otherUnitDataQueueVec_2_enq_valid & ~(_otherUnitDataQueueVec_fifo_2_empty & otherUnitDataQueueVec_2_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_2_deq_ready & ~_otherUnitDataQueueVec_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_2_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_2_empty),
    .almost_empty (otherUnitDataQueueVec_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_2_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_2_full),
    .error        (_otherUnitDataQueueVec_fifo_2_error),
    .data_out     (_otherUnitDataQueueVec_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_3_enq_ready & otherUnitDataQueueVec_3_enq_valid & ~(_otherUnitDataQueueVec_fifo_3_empty & otherUnitDataQueueVec_3_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_3_deq_ready & ~_otherUnitDataQueueVec_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_3_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_3_empty),
    .almost_empty (otherUnitDataQueueVec_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_3_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_3_full),
    .error        (_otherUnitDataQueueVec_fifo_3_error),
    .data_out     (_otherUnitDataQueueVec_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_enq_ready & writeIndexQueue_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_deq_ready & ~_writeIndexQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_enq_bits),
    .empty        (_writeIndexQueue_fifo_empty),
    .almost_empty (writeIndexQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_almostFull),
    .full         (_writeIndexQueue_fifo_full),
    .error        (_writeIndexQueue_fifo_error),
    .data_out     (writeIndexQueue_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_1_enq_ready & writeIndexQueue_1_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_1_deq_ready & ~_writeIndexQueue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_1_enq_bits),
    .empty        (_writeIndexQueue_fifo_1_empty),
    .almost_empty (writeIndexQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_1_almostFull),
    .full         (_writeIndexQueue_fifo_1_full),
    .error        (_writeIndexQueue_fifo_1_error),
    .data_out     (writeIndexQueue_1_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_2_enq_ready & writeIndexQueue_2_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_2_deq_ready & ~_writeIndexQueue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_2_enq_bits),
    .empty        (_writeIndexQueue_fifo_2_empty),
    .almost_empty (writeIndexQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_2_almostFull),
    .full         (_writeIndexQueue_fifo_2_full),
    .error        (_writeIndexQueue_fifo_2_error),
    .data_out     (writeIndexQueue_2_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_3_enq_ready & writeIndexQueue_3_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_3_deq_ready & ~_writeIndexQueue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_3_enq_bits),
    .empty        (_writeIndexQueue_fifo_3_empty),
    .almost_empty (writeIndexQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_3_almostFull),
    .full         (_writeIndexQueue_fifo_3_full),
    .error        (_writeIndexQueue_fifo_3_error),
    .data_out     (writeIndexQueue_3_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(32),
    .err_mode(2),
    .rst_mode(3),
    .width(10)
  ) sourceQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sourceQueue_enq_ready & sourceQueue_enq_valid)),
    .pop_req_n    (~(sourceQueue_deq_ready & ~_sourceQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (sourceQueue_enq_bits),
    .empty        (_sourceQueue_fifo_empty),
    .almost_empty (sourceQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sourceQueue_almostFull),
    .full         (_sourceQueue_fifo_full),
    .error        (_sourceQueue_fifo_error),
    .data_out     (sourceQueue_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(2),
    .err_mode(2),
    .rst_mode(3),
    .width(186)
  ) dataQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(dataQueue_enq_ready & dataQueue_enq_valid)),
    .pop_req_n    (~(dataQueue_deq_ready & ~_dataQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (dataQueue_dataIn),
    .empty        (_dataQueue_fifo_empty),
    .almost_empty (dataQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (dataQueue_almostFull),
    .full         (_dataQueue_fifo_full),
    .error        (_dataQueue_fifo_error),
    .data_out     (_dataQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(32),
    .err_mode(2),
    .rst_mode(3),
    .width(7)
  ) simpleSourceQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(simpleSourceQueue_enq_ready & simpleSourceQueue_enq_valid)),
    .pop_req_n    (~(simpleSourceQueue_deq_ready & ~_simpleSourceQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (simpleSourceQueue_enq_bits),
    .empty        (_simpleSourceQueue_fifo_empty),
    .almost_empty (simpleSourceQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (simpleSourceQueue_almostFull),
    .full         (_simpleSourceQueue_fifo_full),
    .error        (_simpleSourceQueue_fifo_error),
    .data_out     (simpleSourceQueue_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(2),
    .err_mode(2),
    .rst_mode(3),
    .width(78)
  ) simpleDataQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(simpleDataQueue_enq_ready & simpleDataQueue_enq_valid)),
    .pop_req_n    (~(simpleDataQueue_deq_ready & ~_simpleDataQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (simpleDataQueue_dataIn),
    .empty        (_simpleDataQueue_fifo_empty),
    .almost_empty (simpleDataQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (simpleDataQueue_almostFull),
    .full         (_simpleDataQueue_fifo_full),
    .error        (_simpleDataQueue_fifo_error),
    .data_out     (_simpleDataQueue_fifo_data_out)
  );
  assign request_ready = request_ready_0;
  assign axi4Port_aw_valid = axi4Port_aw_valid_0;
  assign axi4Port_aw_bits_id = axi4Port_aw_bits_id_0;
  assign axi4Port_aw_bits_addr = axi4Port_aw_bits_addr_0;
  assign axi4Port_w_valid = axi4Port_w_valid_0;
  assign axi4Port_w_bits_data = axi4Port_w_bits_data_0;
  assign axi4Port_w_bits_strb = axi4Port_w_bits_strb_0;
  assign axi4Port_ar_valid = axi4Port_ar_valid_0;
  assign axi4Port_ar_bits_addr = axi4Port_ar_bits_addr_0;
  assign axi4Port_r_ready = axi4Port_r_ready_0;
  assign simpleAccessPorts_aw_valid = simpleAccessPorts_aw_valid_0;
  assign simpleAccessPorts_aw_bits_id = simpleAccessPorts_aw_bits_id_0;
  assign simpleAccessPorts_aw_bits_addr = simpleAccessPorts_aw_bits_addr_0;
  assign simpleAccessPorts_aw_bits_size = simpleAccessPorts_aw_bits_size_0;
  assign simpleAccessPorts_w_valid = simpleAccessPorts_w_valid_0;
  assign simpleAccessPorts_w_bits_data = simpleAccessPorts_w_bits_data_0;
  assign simpleAccessPorts_w_bits_strb = simpleAccessPorts_w_bits_strb_0;
  assign simpleAccessPorts_ar_valid = simpleAccessPorts_ar_valid_0;
  assign simpleAccessPorts_ar_bits_addr = simpleAccessPorts_ar_bits_addr_0;
  assign simpleAccessPorts_r_ready = simpleAccessPorts_r_ready_0;
  assign vrfReadDataPorts_0_valid = vrfReadDataPorts_0_valid_0;
  assign vrfReadDataPorts_0_bits_vs = vrfReadDataPorts_0_bits_vs_0;
  assign vrfReadDataPorts_0_bits_offset = vrfReadDataPorts_0_bits_offset_0;
  assign vrfReadDataPorts_0_bits_instructionIndex = vrfReadDataPorts_0_bits_instructionIndex_0;
  assign vrfReadDataPorts_1_valid = vrfReadDataPorts_1_valid_0;
  assign vrfReadDataPorts_1_bits_vs = vrfReadDataPorts_1_bits_vs_0;
  assign vrfReadDataPorts_1_bits_offset = vrfReadDataPorts_1_bits_offset_0;
  assign vrfReadDataPorts_1_bits_instructionIndex = vrfReadDataPorts_1_bits_instructionIndex_0;
  assign vrfReadDataPorts_2_valid = vrfReadDataPorts_2_valid_0;
  assign vrfReadDataPorts_2_bits_vs = vrfReadDataPorts_2_bits_vs_0;
  assign vrfReadDataPorts_2_bits_offset = vrfReadDataPorts_2_bits_offset_0;
  assign vrfReadDataPorts_2_bits_instructionIndex = vrfReadDataPorts_2_bits_instructionIndex_0;
  assign vrfReadDataPorts_3_valid = vrfReadDataPorts_3_valid_0;
  assign vrfReadDataPorts_3_bits_vs = vrfReadDataPorts_3_bits_vs_0;
  assign vrfReadDataPorts_3_bits_offset = vrfReadDataPorts_3_bits_offset_0;
  assign vrfReadDataPorts_3_bits_instructionIndex = vrfReadDataPorts_3_bits_instructionIndex_0;
  assign vrfWritePort_0_valid = vrfWritePort_0_valid_0;
  assign vrfWritePort_0_bits_vd = vrfWritePort_0_bits_vd_0;
  assign vrfWritePort_0_bits_offset = vrfWritePort_0_bits_offset_0;
  assign vrfWritePort_0_bits_mask = vrfWritePort_0_bits_mask_0;
  assign vrfWritePort_0_bits_data = vrfWritePort_0_bits_data_0;
  assign vrfWritePort_0_bits_last = vrfWritePort_0_bits_last_0;
  assign vrfWritePort_0_bits_instructionIndex = vrfWritePort_0_bits_instructionIndex_0;
  assign vrfWritePort_1_valid = vrfWritePort_1_valid_0;
  assign vrfWritePort_1_bits_vd = vrfWritePort_1_bits_vd_0;
  assign vrfWritePort_1_bits_offset = vrfWritePort_1_bits_offset_0;
  assign vrfWritePort_1_bits_mask = vrfWritePort_1_bits_mask_0;
  assign vrfWritePort_1_bits_data = vrfWritePort_1_bits_data_0;
  assign vrfWritePort_1_bits_last = vrfWritePort_1_bits_last_0;
  assign vrfWritePort_1_bits_instructionIndex = vrfWritePort_1_bits_instructionIndex_0;
  assign vrfWritePort_2_valid = vrfWritePort_2_valid_0;
  assign vrfWritePort_2_bits_vd = vrfWritePort_2_bits_vd_0;
  assign vrfWritePort_2_bits_offset = vrfWritePort_2_bits_offset_0;
  assign vrfWritePort_2_bits_mask = vrfWritePort_2_bits_mask_0;
  assign vrfWritePort_2_bits_data = vrfWritePort_2_bits_data_0;
  assign vrfWritePort_2_bits_last = vrfWritePort_2_bits_last_0;
  assign vrfWritePort_2_bits_instructionIndex = vrfWritePort_2_bits_instructionIndex_0;
  assign vrfWritePort_3_valid = vrfWritePort_3_valid_0;
  assign vrfWritePort_3_bits_vd = vrfWritePort_3_bits_vd_0;
  assign vrfWritePort_3_bits_offset = vrfWritePort_3_bits_offset_0;
  assign vrfWritePort_3_bits_mask = vrfWritePort_3_bits_mask_0;
  assign vrfWritePort_3_bits_data = vrfWritePort_3_bits_data_0;
  assign vrfWritePort_3_bits_last = vrfWritePort_3_bits_last_0;
  assign vrfWritePort_3_bits_instructionIndex = vrfWritePort_3_bits_instructionIndex_0;
  assign dataInWriteQueue_0 = {dataInWriteQueue_0_hi, dataInWriteQueue_0_lo} | dataInMSHR;
  assign dataInWriteQueue_1 = {dataInWriteQueue_1_hi, dataInWriteQueue_1_lo} | dataInMSHR;
  assign dataInWriteQueue_2 = {dataInWriteQueue_2_hi, dataInWriteQueue_2_lo} | dataInMSHR;
  assign dataInWriteQueue_3 = {dataInWriteQueue_3_hi, dataInWriteQueue_3_lo} | dataInMSHR;
  assign lastReport = (_loadUnit_status_last ? 8'h1 << _GEN_130 : 8'h0) | (_storeUnit_status_last ? 8'h1 << _storeUnit_status_instructionIndex : 8'h0) | (_otherUnit_status_last ? 8'h1 << _GEN_131 : 8'h0);
  assign tokenIO_offsetGroupRelease = {tokenIO_offsetGroupRelease_hi, tokenIO_offsetGroupRelease_lo};
endmodule

