module LaneLogic(
  input  [31:0] req_src_0,
                req_src_1,
  input  [3:0]  req_opcode,
  output [31:0] resp
);

  wire [4:0]  view__resp_plaInput;
  wire [4:0]  view__resp_invInputs = ~view__resp_plaInput;
  wire        view__resp_invMatrixOutputs;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0 = view__resp_plaInput[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_1 = view__resp_plaInput[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_3 = view__resp_plaInput[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1 = view__resp_plaInput[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_2 = view__resp_plaInput[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_4 = view__resp_plaInput[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2 = view__resp_invInputs[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_1 = view__resp_invInputs[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_2 = view__resp_invInputs[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3 = view__resp_invInputs[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_1 = view__resp_invInputs[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_2 = view__resp_invInputs[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4 = view__resp_invInputs[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_1 = view__resp_invInputs[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo = {view__resp_andMatrixOutputs_andMatrixInput_2, view__resp_andMatrixOutputs_andMatrixInput_3};
  wire [1:0]  view__resp_andMatrixOutputs_hi = {view__resp_andMatrixOutputs_andMatrixInput_0, view__resp_andMatrixOutputs_andMatrixInput_1};
  wire        view__resp_andMatrixOutputs_4_2 = &{view__resp_andMatrixOutputs_hi, view__resp_andMatrixOutputs_lo};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_1 = view__resp_plaInput[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_2 = view__resp_plaInput[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_1 = {view__resp_andMatrixOutputs_andMatrixInput_2_1, view__resp_andMatrixOutputs_andMatrixInput_3_1};
  wire [1:0]  view__resp_andMatrixOutputs_hi_1 = {view__resp_andMatrixOutputs_andMatrixInput_0_1, view__resp_andMatrixOutputs_andMatrixInput_1_1};
  wire        view__resp_andMatrixOutputs_1_2 = &{view__resp_andMatrixOutputs_hi_1, view__resp_andMatrixOutputs_lo_1};
  wire [1:0]  view__resp_andMatrixOutputs_lo_2 = {view__resp_andMatrixOutputs_andMatrixInput_2_2, view__resp_andMatrixOutputs_andMatrixInput_3_2};
  wire [1:0]  view__resp_andMatrixOutputs_hi_2 = {view__resp_andMatrixOutputs_andMatrixInput_0_2, view__resp_andMatrixOutputs_andMatrixInput_1_2};
  wire        view__resp_andMatrixOutputs_3_2 = &{view__resp_andMatrixOutputs_hi_2, view__resp_andMatrixOutputs_lo_2};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_3 = view__resp_invInputs[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_3 = view__resp_invInputs[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_4 = view__resp_invInputs[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_3 = view__resp_plaInput[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_4 = view__resp_plaInput[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_3 = {view__resp_andMatrixOutputs_andMatrixInput_3_3, view__resp_andMatrixOutputs_andMatrixInput_4};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi = {view__resp_andMatrixOutputs_andMatrixInput_0_3, view__resp_andMatrixOutputs_andMatrixInput_1_3};
  wire [2:0]  view__resp_andMatrixOutputs_hi_3 = {view__resp_andMatrixOutputs_hi_hi, view__resp_andMatrixOutputs_andMatrixInput_2_3};
  wire        view__resp_andMatrixOutputs_0_2 = &{view__resp_andMatrixOutputs_hi_3, view__resp_andMatrixOutputs_lo_3};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_4 = view__resp_invInputs[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_4 = {view__resp_andMatrixOutputs_andMatrixInput_3_4, view__resp_andMatrixOutputs_andMatrixInput_4_1};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_1 = {view__resp_andMatrixOutputs_andMatrixInput_0_4, view__resp_andMatrixOutputs_andMatrixInput_1_4};
  wire [2:0]  view__resp_andMatrixOutputs_hi_4 = {view__resp_andMatrixOutputs_hi_hi_1, view__resp_andMatrixOutputs_andMatrixInput_2_4};
  wire        view__resp_andMatrixOutputs_2_2 = &{view__resp_andMatrixOutputs_hi_4, view__resp_andMatrixOutputs_lo_4};
  wire [1:0]  view__resp_orMatrixOutputs_lo = {view__resp_andMatrixOutputs_0_2, view__resp_andMatrixOutputs_2_2};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi = {view__resp_andMatrixOutputs_4_2, view__resp_andMatrixOutputs_1_2};
  wire [2:0]  view__resp_orMatrixOutputs_hi = {view__resp_orMatrixOutputs_hi_hi, view__resp_andMatrixOutputs_3_2};
  wire        view__resp_orMatrixOutputs = |{view__resp_orMatrixOutputs_hi, view__resp_orMatrixOutputs_lo};
  assign view__resp_invMatrixOutputs = view__resp_orMatrixOutputs;
  wire        view__resp_plaOutput = view__resp_invMatrixOutputs;
  assign view__resp_plaInput = {1'h0, req_opcode[1:0], req_src_0[0], req_opcode[2] ^ req_src_1[0]};
  wire [4:0]  view__resp_plaInput_1;
  wire [4:0]  view__resp_invInputs_1 = ~view__resp_plaInput_1;
  wire        view__resp_invMatrixOutputs_1;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_5 = view__resp_plaInput_1[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_6 = view__resp_plaInput_1[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_8 = view__resp_plaInput_1[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_5 = view__resp_plaInput_1[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_7 = view__resp_plaInput_1[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_9 = view__resp_plaInput_1[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_5 = view__resp_invInputs_1[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_6 = view__resp_invInputs_1[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_7 = view__resp_invInputs_1[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_5 = view__resp_invInputs_1[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_6 = view__resp_invInputs_1[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_7 = view__resp_invInputs_1[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_2 = view__resp_invInputs_1[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_3 = view__resp_invInputs_1[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_5 = {view__resp_andMatrixOutputs_andMatrixInput_2_5, view__resp_andMatrixOutputs_andMatrixInput_3_5};
  wire [1:0]  view__resp_andMatrixOutputs_hi_5 = {view__resp_andMatrixOutputs_andMatrixInput_0_5, view__resp_andMatrixOutputs_andMatrixInput_1_5};
  wire        view__resp_andMatrixOutputs_4_2_1 = &{view__resp_andMatrixOutputs_hi_5, view__resp_andMatrixOutputs_lo_5};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_6 = view__resp_plaInput_1[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_7 = view__resp_plaInput_1[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_6 = {view__resp_andMatrixOutputs_andMatrixInput_2_6, view__resp_andMatrixOutputs_andMatrixInput_3_6};
  wire [1:0]  view__resp_andMatrixOutputs_hi_6 = {view__resp_andMatrixOutputs_andMatrixInput_0_6, view__resp_andMatrixOutputs_andMatrixInput_1_6};
  wire        view__resp_andMatrixOutputs_1_2_1 = &{view__resp_andMatrixOutputs_hi_6, view__resp_andMatrixOutputs_lo_6};
  wire [1:0]  view__resp_andMatrixOutputs_lo_7 = {view__resp_andMatrixOutputs_andMatrixInput_2_7, view__resp_andMatrixOutputs_andMatrixInput_3_7};
  wire [1:0]  view__resp_andMatrixOutputs_hi_7 = {view__resp_andMatrixOutputs_andMatrixInput_0_7, view__resp_andMatrixOutputs_andMatrixInput_1_7};
  wire        view__resp_andMatrixOutputs_3_2_1 = &{view__resp_andMatrixOutputs_hi_7, view__resp_andMatrixOutputs_lo_7};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_8 = view__resp_invInputs_1[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_8 = view__resp_invInputs_1[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_9 = view__resp_invInputs_1[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_8 = view__resp_plaInput_1[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_9 = view__resp_plaInput_1[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_8 = {view__resp_andMatrixOutputs_andMatrixInput_3_8, view__resp_andMatrixOutputs_andMatrixInput_4_2};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_2 = {view__resp_andMatrixOutputs_andMatrixInput_0_8, view__resp_andMatrixOutputs_andMatrixInput_1_8};
  wire [2:0]  view__resp_andMatrixOutputs_hi_8 = {view__resp_andMatrixOutputs_hi_hi_2, view__resp_andMatrixOutputs_andMatrixInput_2_8};
  wire        view__resp_andMatrixOutputs_0_2_1 = &{view__resp_andMatrixOutputs_hi_8, view__resp_andMatrixOutputs_lo_8};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_9 = view__resp_invInputs_1[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_9 = {view__resp_andMatrixOutputs_andMatrixInput_3_9, view__resp_andMatrixOutputs_andMatrixInput_4_3};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_3 = {view__resp_andMatrixOutputs_andMatrixInput_0_9, view__resp_andMatrixOutputs_andMatrixInput_1_9};
  wire [2:0]  view__resp_andMatrixOutputs_hi_9 = {view__resp_andMatrixOutputs_hi_hi_3, view__resp_andMatrixOutputs_andMatrixInput_2_9};
  wire        view__resp_andMatrixOutputs_2_2_1 = &{view__resp_andMatrixOutputs_hi_9, view__resp_andMatrixOutputs_lo_9};
  wire [1:0]  view__resp_orMatrixOutputs_lo_1 = {view__resp_andMatrixOutputs_0_2_1, view__resp_andMatrixOutputs_2_2_1};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_1 = {view__resp_andMatrixOutputs_4_2_1, view__resp_andMatrixOutputs_1_2_1};
  wire [2:0]  view__resp_orMatrixOutputs_hi_1 = {view__resp_orMatrixOutputs_hi_hi_1, view__resp_andMatrixOutputs_3_2_1};
  wire        view__resp_orMatrixOutputs_1 = |{view__resp_orMatrixOutputs_hi_1, view__resp_orMatrixOutputs_lo_1};
  assign view__resp_invMatrixOutputs_1 = view__resp_orMatrixOutputs_1;
  wire        view__resp_plaOutput_1 = view__resp_invMatrixOutputs_1;
  assign view__resp_plaInput_1 = {1'h0, req_opcode[1:0], req_src_0[1], req_opcode[2] ^ req_src_1[1]};
  wire [4:0]  view__resp_plaInput_2;
  wire [4:0]  view__resp_invInputs_2 = ~view__resp_plaInput_2;
  wire        view__resp_invMatrixOutputs_2;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_10 = view__resp_plaInput_2[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_11 = view__resp_plaInput_2[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_13 = view__resp_plaInput_2[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_10 = view__resp_plaInput_2[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_12 = view__resp_plaInput_2[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_14 = view__resp_plaInput_2[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_10 = view__resp_invInputs_2[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_11 = view__resp_invInputs_2[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_12 = view__resp_invInputs_2[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_10 = view__resp_invInputs_2[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_11 = view__resp_invInputs_2[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_12 = view__resp_invInputs_2[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_4 = view__resp_invInputs_2[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_5 = view__resp_invInputs_2[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_10 = {view__resp_andMatrixOutputs_andMatrixInput_2_10, view__resp_andMatrixOutputs_andMatrixInput_3_10};
  wire [1:0]  view__resp_andMatrixOutputs_hi_10 = {view__resp_andMatrixOutputs_andMatrixInput_0_10, view__resp_andMatrixOutputs_andMatrixInput_1_10};
  wire        view__resp_andMatrixOutputs_4_2_2 = &{view__resp_andMatrixOutputs_hi_10, view__resp_andMatrixOutputs_lo_10};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_11 = view__resp_plaInput_2[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_12 = view__resp_plaInput_2[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_11 = {view__resp_andMatrixOutputs_andMatrixInput_2_11, view__resp_andMatrixOutputs_andMatrixInput_3_11};
  wire [1:0]  view__resp_andMatrixOutputs_hi_11 = {view__resp_andMatrixOutputs_andMatrixInput_0_11, view__resp_andMatrixOutputs_andMatrixInput_1_11};
  wire        view__resp_andMatrixOutputs_1_2_2 = &{view__resp_andMatrixOutputs_hi_11, view__resp_andMatrixOutputs_lo_11};
  wire [1:0]  view__resp_andMatrixOutputs_lo_12 = {view__resp_andMatrixOutputs_andMatrixInput_2_12, view__resp_andMatrixOutputs_andMatrixInput_3_12};
  wire [1:0]  view__resp_andMatrixOutputs_hi_12 = {view__resp_andMatrixOutputs_andMatrixInput_0_12, view__resp_andMatrixOutputs_andMatrixInput_1_12};
  wire        view__resp_andMatrixOutputs_3_2_2 = &{view__resp_andMatrixOutputs_hi_12, view__resp_andMatrixOutputs_lo_12};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_13 = view__resp_invInputs_2[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_13 = view__resp_invInputs_2[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_14 = view__resp_invInputs_2[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_13 = view__resp_plaInput_2[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_14 = view__resp_plaInput_2[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_13 = {view__resp_andMatrixOutputs_andMatrixInput_3_13, view__resp_andMatrixOutputs_andMatrixInput_4_4};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_4 = {view__resp_andMatrixOutputs_andMatrixInput_0_13, view__resp_andMatrixOutputs_andMatrixInput_1_13};
  wire [2:0]  view__resp_andMatrixOutputs_hi_13 = {view__resp_andMatrixOutputs_hi_hi_4, view__resp_andMatrixOutputs_andMatrixInput_2_13};
  wire        view__resp_andMatrixOutputs_0_2_2 = &{view__resp_andMatrixOutputs_hi_13, view__resp_andMatrixOutputs_lo_13};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_14 = view__resp_invInputs_2[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_14 = {view__resp_andMatrixOutputs_andMatrixInput_3_14, view__resp_andMatrixOutputs_andMatrixInput_4_5};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_5 = {view__resp_andMatrixOutputs_andMatrixInput_0_14, view__resp_andMatrixOutputs_andMatrixInput_1_14};
  wire [2:0]  view__resp_andMatrixOutputs_hi_14 = {view__resp_andMatrixOutputs_hi_hi_5, view__resp_andMatrixOutputs_andMatrixInput_2_14};
  wire        view__resp_andMatrixOutputs_2_2_2 = &{view__resp_andMatrixOutputs_hi_14, view__resp_andMatrixOutputs_lo_14};
  wire [1:0]  view__resp_orMatrixOutputs_lo_2 = {view__resp_andMatrixOutputs_0_2_2, view__resp_andMatrixOutputs_2_2_2};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_2 = {view__resp_andMatrixOutputs_4_2_2, view__resp_andMatrixOutputs_1_2_2};
  wire [2:0]  view__resp_orMatrixOutputs_hi_2 = {view__resp_orMatrixOutputs_hi_hi_2, view__resp_andMatrixOutputs_3_2_2};
  wire        view__resp_orMatrixOutputs_2 = |{view__resp_orMatrixOutputs_hi_2, view__resp_orMatrixOutputs_lo_2};
  assign view__resp_invMatrixOutputs_2 = view__resp_orMatrixOutputs_2;
  wire        view__resp_plaOutput_2 = view__resp_invMatrixOutputs_2;
  assign view__resp_plaInput_2 = {1'h0, req_opcode[1:0], req_src_0[2], req_opcode[2] ^ req_src_1[2]};
  wire [4:0]  view__resp_plaInput_3;
  wire [4:0]  view__resp_invInputs_3 = ~view__resp_plaInput_3;
  wire        view__resp_invMatrixOutputs_3;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_15 = view__resp_plaInput_3[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_16 = view__resp_plaInput_3[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_18 = view__resp_plaInput_3[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_15 = view__resp_plaInput_3[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_17 = view__resp_plaInput_3[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_19 = view__resp_plaInput_3[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_15 = view__resp_invInputs_3[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_16 = view__resp_invInputs_3[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_17 = view__resp_invInputs_3[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_15 = view__resp_invInputs_3[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_16 = view__resp_invInputs_3[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_17 = view__resp_invInputs_3[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_6 = view__resp_invInputs_3[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_7 = view__resp_invInputs_3[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_15 = {view__resp_andMatrixOutputs_andMatrixInput_2_15, view__resp_andMatrixOutputs_andMatrixInput_3_15};
  wire [1:0]  view__resp_andMatrixOutputs_hi_15 = {view__resp_andMatrixOutputs_andMatrixInput_0_15, view__resp_andMatrixOutputs_andMatrixInput_1_15};
  wire        view__resp_andMatrixOutputs_4_2_3 = &{view__resp_andMatrixOutputs_hi_15, view__resp_andMatrixOutputs_lo_15};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_16 = view__resp_plaInput_3[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_17 = view__resp_plaInput_3[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_16 = {view__resp_andMatrixOutputs_andMatrixInput_2_16, view__resp_andMatrixOutputs_andMatrixInput_3_16};
  wire [1:0]  view__resp_andMatrixOutputs_hi_16 = {view__resp_andMatrixOutputs_andMatrixInput_0_16, view__resp_andMatrixOutputs_andMatrixInput_1_16};
  wire        view__resp_andMatrixOutputs_1_2_3 = &{view__resp_andMatrixOutputs_hi_16, view__resp_andMatrixOutputs_lo_16};
  wire [1:0]  view__resp_andMatrixOutputs_lo_17 = {view__resp_andMatrixOutputs_andMatrixInput_2_17, view__resp_andMatrixOutputs_andMatrixInput_3_17};
  wire [1:0]  view__resp_andMatrixOutputs_hi_17 = {view__resp_andMatrixOutputs_andMatrixInput_0_17, view__resp_andMatrixOutputs_andMatrixInput_1_17};
  wire        view__resp_andMatrixOutputs_3_2_3 = &{view__resp_andMatrixOutputs_hi_17, view__resp_andMatrixOutputs_lo_17};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_18 = view__resp_invInputs_3[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_18 = view__resp_invInputs_3[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_19 = view__resp_invInputs_3[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_18 = view__resp_plaInput_3[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_19 = view__resp_plaInput_3[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_18 = {view__resp_andMatrixOutputs_andMatrixInput_3_18, view__resp_andMatrixOutputs_andMatrixInput_4_6};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_6 = {view__resp_andMatrixOutputs_andMatrixInput_0_18, view__resp_andMatrixOutputs_andMatrixInput_1_18};
  wire [2:0]  view__resp_andMatrixOutputs_hi_18 = {view__resp_andMatrixOutputs_hi_hi_6, view__resp_andMatrixOutputs_andMatrixInput_2_18};
  wire        view__resp_andMatrixOutputs_0_2_3 = &{view__resp_andMatrixOutputs_hi_18, view__resp_andMatrixOutputs_lo_18};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_19 = view__resp_invInputs_3[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_19 = {view__resp_andMatrixOutputs_andMatrixInput_3_19, view__resp_andMatrixOutputs_andMatrixInput_4_7};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_7 = {view__resp_andMatrixOutputs_andMatrixInput_0_19, view__resp_andMatrixOutputs_andMatrixInput_1_19};
  wire [2:0]  view__resp_andMatrixOutputs_hi_19 = {view__resp_andMatrixOutputs_hi_hi_7, view__resp_andMatrixOutputs_andMatrixInput_2_19};
  wire        view__resp_andMatrixOutputs_2_2_3 = &{view__resp_andMatrixOutputs_hi_19, view__resp_andMatrixOutputs_lo_19};
  wire [1:0]  view__resp_orMatrixOutputs_lo_3 = {view__resp_andMatrixOutputs_0_2_3, view__resp_andMatrixOutputs_2_2_3};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_3 = {view__resp_andMatrixOutputs_4_2_3, view__resp_andMatrixOutputs_1_2_3};
  wire [2:0]  view__resp_orMatrixOutputs_hi_3 = {view__resp_orMatrixOutputs_hi_hi_3, view__resp_andMatrixOutputs_3_2_3};
  wire        view__resp_orMatrixOutputs_3 = |{view__resp_orMatrixOutputs_hi_3, view__resp_orMatrixOutputs_lo_3};
  assign view__resp_invMatrixOutputs_3 = view__resp_orMatrixOutputs_3;
  wire        view__resp_plaOutput_3 = view__resp_invMatrixOutputs_3;
  assign view__resp_plaInput_3 = {1'h0, req_opcode[1:0], req_src_0[3], req_opcode[2] ^ req_src_1[3]};
  wire [4:0]  view__resp_plaInput_4;
  wire [4:0]  view__resp_invInputs_4 = ~view__resp_plaInput_4;
  wire        view__resp_invMatrixOutputs_4;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_20 = view__resp_plaInput_4[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_21 = view__resp_plaInput_4[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_23 = view__resp_plaInput_4[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_20 = view__resp_plaInput_4[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_22 = view__resp_plaInput_4[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_24 = view__resp_plaInput_4[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_20 = view__resp_invInputs_4[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_21 = view__resp_invInputs_4[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_22 = view__resp_invInputs_4[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_20 = view__resp_invInputs_4[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_21 = view__resp_invInputs_4[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_22 = view__resp_invInputs_4[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_8 = view__resp_invInputs_4[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_9 = view__resp_invInputs_4[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_20 = {view__resp_andMatrixOutputs_andMatrixInput_2_20, view__resp_andMatrixOutputs_andMatrixInput_3_20};
  wire [1:0]  view__resp_andMatrixOutputs_hi_20 = {view__resp_andMatrixOutputs_andMatrixInput_0_20, view__resp_andMatrixOutputs_andMatrixInput_1_20};
  wire        view__resp_andMatrixOutputs_4_2_4 = &{view__resp_andMatrixOutputs_hi_20, view__resp_andMatrixOutputs_lo_20};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_21 = view__resp_plaInput_4[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_22 = view__resp_plaInput_4[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_21 = {view__resp_andMatrixOutputs_andMatrixInput_2_21, view__resp_andMatrixOutputs_andMatrixInput_3_21};
  wire [1:0]  view__resp_andMatrixOutputs_hi_21 = {view__resp_andMatrixOutputs_andMatrixInput_0_21, view__resp_andMatrixOutputs_andMatrixInput_1_21};
  wire        view__resp_andMatrixOutputs_1_2_4 = &{view__resp_andMatrixOutputs_hi_21, view__resp_andMatrixOutputs_lo_21};
  wire [1:0]  view__resp_andMatrixOutputs_lo_22 = {view__resp_andMatrixOutputs_andMatrixInput_2_22, view__resp_andMatrixOutputs_andMatrixInput_3_22};
  wire [1:0]  view__resp_andMatrixOutputs_hi_22 = {view__resp_andMatrixOutputs_andMatrixInput_0_22, view__resp_andMatrixOutputs_andMatrixInput_1_22};
  wire        view__resp_andMatrixOutputs_3_2_4 = &{view__resp_andMatrixOutputs_hi_22, view__resp_andMatrixOutputs_lo_22};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_23 = view__resp_invInputs_4[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_23 = view__resp_invInputs_4[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_24 = view__resp_invInputs_4[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_23 = view__resp_plaInput_4[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_24 = view__resp_plaInput_4[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_23 = {view__resp_andMatrixOutputs_andMatrixInput_3_23, view__resp_andMatrixOutputs_andMatrixInput_4_8};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_8 = {view__resp_andMatrixOutputs_andMatrixInput_0_23, view__resp_andMatrixOutputs_andMatrixInput_1_23};
  wire [2:0]  view__resp_andMatrixOutputs_hi_23 = {view__resp_andMatrixOutputs_hi_hi_8, view__resp_andMatrixOutputs_andMatrixInput_2_23};
  wire        view__resp_andMatrixOutputs_0_2_4 = &{view__resp_andMatrixOutputs_hi_23, view__resp_andMatrixOutputs_lo_23};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_24 = view__resp_invInputs_4[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_24 = {view__resp_andMatrixOutputs_andMatrixInput_3_24, view__resp_andMatrixOutputs_andMatrixInput_4_9};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_9 = {view__resp_andMatrixOutputs_andMatrixInput_0_24, view__resp_andMatrixOutputs_andMatrixInput_1_24};
  wire [2:0]  view__resp_andMatrixOutputs_hi_24 = {view__resp_andMatrixOutputs_hi_hi_9, view__resp_andMatrixOutputs_andMatrixInput_2_24};
  wire        view__resp_andMatrixOutputs_2_2_4 = &{view__resp_andMatrixOutputs_hi_24, view__resp_andMatrixOutputs_lo_24};
  wire [1:0]  view__resp_orMatrixOutputs_lo_4 = {view__resp_andMatrixOutputs_0_2_4, view__resp_andMatrixOutputs_2_2_4};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_4 = {view__resp_andMatrixOutputs_4_2_4, view__resp_andMatrixOutputs_1_2_4};
  wire [2:0]  view__resp_orMatrixOutputs_hi_4 = {view__resp_orMatrixOutputs_hi_hi_4, view__resp_andMatrixOutputs_3_2_4};
  wire        view__resp_orMatrixOutputs_4 = |{view__resp_orMatrixOutputs_hi_4, view__resp_orMatrixOutputs_lo_4};
  assign view__resp_invMatrixOutputs_4 = view__resp_orMatrixOutputs_4;
  wire        view__resp_plaOutput_4 = view__resp_invMatrixOutputs_4;
  assign view__resp_plaInput_4 = {1'h0, req_opcode[1:0], req_src_0[4], req_opcode[2] ^ req_src_1[4]};
  wire [4:0]  view__resp_plaInput_5;
  wire [4:0]  view__resp_invInputs_5 = ~view__resp_plaInput_5;
  wire        view__resp_invMatrixOutputs_5;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_25 = view__resp_plaInput_5[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_26 = view__resp_plaInput_5[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_28 = view__resp_plaInput_5[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_25 = view__resp_plaInput_5[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_27 = view__resp_plaInput_5[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_29 = view__resp_plaInput_5[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_25 = view__resp_invInputs_5[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_26 = view__resp_invInputs_5[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_27 = view__resp_invInputs_5[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_25 = view__resp_invInputs_5[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_26 = view__resp_invInputs_5[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_27 = view__resp_invInputs_5[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_10 = view__resp_invInputs_5[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_11 = view__resp_invInputs_5[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_25 = {view__resp_andMatrixOutputs_andMatrixInput_2_25, view__resp_andMatrixOutputs_andMatrixInput_3_25};
  wire [1:0]  view__resp_andMatrixOutputs_hi_25 = {view__resp_andMatrixOutputs_andMatrixInput_0_25, view__resp_andMatrixOutputs_andMatrixInput_1_25};
  wire        view__resp_andMatrixOutputs_4_2_5 = &{view__resp_andMatrixOutputs_hi_25, view__resp_andMatrixOutputs_lo_25};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_26 = view__resp_plaInput_5[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_27 = view__resp_plaInput_5[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_26 = {view__resp_andMatrixOutputs_andMatrixInput_2_26, view__resp_andMatrixOutputs_andMatrixInput_3_26};
  wire [1:0]  view__resp_andMatrixOutputs_hi_26 = {view__resp_andMatrixOutputs_andMatrixInput_0_26, view__resp_andMatrixOutputs_andMatrixInput_1_26};
  wire        view__resp_andMatrixOutputs_1_2_5 = &{view__resp_andMatrixOutputs_hi_26, view__resp_andMatrixOutputs_lo_26};
  wire [1:0]  view__resp_andMatrixOutputs_lo_27 = {view__resp_andMatrixOutputs_andMatrixInput_2_27, view__resp_andMatrixOutputs_andMatrixInput_3_27};
  wire [1:0]  view__resp_andMatrixOutputs_hi_27 = {view__resp_andMatrixOutputs_andMatrixInput_0_27, view__resp_andMatrixOutputs_andMatrixInput_1_27};
  wire        view__resp_andMatrixOutputs_3_2_5 = &{view__resp_andMatrixOutputs_hi_27, view__resp_andMatrixOutputs_lo_27};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_28 = view__resp_invInputs_5[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_28 = view__resp_invInputs_5[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_29 = view__resp_invInputs_5[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_28 = view__resp_plaInput_5[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_29 = view__resp_plaInput_5[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_28 = {view__resp_andMatrixOutputs_andMatrixInput_3_28, view__resp_andMatrixOutputs_andMatrixInput_4_10};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_10 = {view__resp_andMatrixOutputs_andMatrixInput_0_28, view__resp_andMatrixOutputs_andMatrixInput_1_28};
  wire [2:0]  view__resp_andMatrixOutputs_hi_28 = {view__resp_andMatrixOutputs_hi_hi_10, view__resp_andMatrixOutputs_andMatrixInput_2_28};
  wire        view__resp_andMatrixOutputs_0_2_5 = &{view__resp_andMatrixOutputs_hi_28, view__resp_andMatrixOutputs_lo_28};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_29 = view__resp_invInputs_5[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_29 = {view__resp_andMatrixOutputs_andMatrixInput_3_29, view__resp_andMatrixOutputs_andMatrixInput_4_11};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_11 = {view__resp_andMatrixOutputs_andMatrixInput_0_29, view__resp_andMatrixOutputs_andMatrixInput_1_29};
  wire [2:0]  view__resp_andMatrixOutputs_hi_29 = {view__resp_andMatrixOutputs_hi_hi_11, view__resp_andMatrixOutputs_andMatrixInput_2_29};
  wire        view__resp_andMatrixOutputs_2_2_5 = &{view__resp_andMatrixOutputs_hi_29, view__resp_andMatrixOutputs_lo_29};
  wire [1:0]  view__resp_orMatrixOutputs_lo_5 = {view__resp_andMatrixOutputs_0_2_5, view__resp_andMatrixOutputs_2_2_5};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_5 = {view__resp_andMatrixOutputs_4_2_5, view__resp_andMatrixOutputs_1_2_5};
  wire [2:0]  view__resp_orMatrixOutputs_hi_5 = {view__resp_orMatrixOutputs_hi_hi_5, view__resp_andMatrixOutputs_3_2_5};
  wire        view__resp_orMatrixOutputs_5 = |{view__resp_orMatrixOutputs_hi_5, view__resp_orMatrixOutputs_lo_5};
  assign view__resp_invMatrixOutputs_5 = view__resp_orMatrixOutputs_5;
  wire        view__resp_plaOutput_5 = view__resp_invMatrixOutputs_5;
  assign view__resp_plaInput_5 = {1'h0, req_opcode[1:0], req_src_0[5], req_opcode[2] ^ req_src_1[5]};
  wire [4:0]  view__resp_plaInput_6;
  wire [4:0]  view__resp_invInputs_6 = ~view__resp_plaInput_6;
  wire        view__resp_invMatrixOutputs_6;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_30 = view__resp_plaInput_6[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_31 = view__resp_plaInput_6[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_33 = view__resp_plaInput_6[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_30 = view__resp_plaInput_6[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_32 = view__resp_plaInput_6[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_34 = view__resp_plaInput_6[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_30 = view__resp_invInputs_6[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_31 = view__resp_invInputs_6[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_32 = view__resp_invInputs_6[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_30 = view__resp_invInputs_6[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_31 = view__resp_invInputs_6[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_32 = view__resp_invInputs_6[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_12 = view__resp_invInputs_6[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_13 = view__resp_invInputs_6[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_30 = {view__resp_andMatrixOutputs_andMatrixInput_2_30, view__resp_andMatrixOutputs_andMatrixInput_3_30};
  wire [1:0]  view__resp_andMatrixOutputs_hi_30 = {view__resp_andMatrixOutputs_andMatrixInput_0_30, view__resp_andMatrixOutputs_andMatrixInput_1_30};
  wire        view__resp_andMatrixOutputs_4_2_6 = &{view__resp_andMatrixOutputs_hi_30, view__resp_andMatrixOutputs_lo_30};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_31 = view__resp_plaInput_6[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_32 = view__resp_plaInput_6[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_31 = {view__resp_andMatrixOutputs_andMatrixInput_2_31, view__resp_andMatrixOutputs_andMatrixInput_3_31};
  wire [1:0]  view__resp_andMatrixOutputs_hi_31 = {view__resp_andMatrixOutputs_andMatrixInput_0_31, view__resp_andMatrixOutputs_andMatrixInput_1_31};
  wire        view__resp_andMatrixOutputs_1_2_6 = &{view__resp_andMatrixOutputs_hi_31, view__resp_andMatrixOutputs_lo_31};
  wire [1:0]  view__resp_andMatrixOutputs_lo_32 = {view__resp_andMatrixOutputs_andMatrixInput_2_32, view__resp_andMatrixOutputs_andMatrixInput_3_32};
  wire [1:0]  view__resp_andMatrixOutputs_hi_32 = {view__resp_andMatrixOutputs_andMatrixInput_0_32, view__resp_andMatrixOutputs_andMatrixInput_1_32};
  wire        view__resp_andMatrixOutputs_3_2_6 = &{view__resp_andMatrixOutputs_hi_32, view__resp_andMatrixOutputs_lo_32};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_33 = view__resp_invInputs_6[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_33 = view__resp_invInputs_6[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_34 = view__resp_invInputs_6[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_33 = view__resp_plaInput_6[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_34 = view__resp_plaInput_6[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_33 = {view__resp_andMatrixOutputs_andMatrixInput_3_33, view__resp_andMatrixOutputs_andMatrixInput_4_12};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_12 = {view__resp_andMatrixOutputs_andMatrixInput_0_33, view__resp_andMatrixOutputs_andMatrixInput_1_33};
  wire [2:0]  view__resp_andMatrixOutputs_hi_33 = {view__resp_andMatrixOutputs_hi_hi_12, view__resp_andMatrixOutputs_andMatrixInput_2_33};
  wire        view__resp_andMatrixOutputs_0_2_6 = &{view__resp_andMatrixOutputs_hi_33, view__resp_andMatrixOutputs_lo_33};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_34 = view__resp_invInputs_6[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_34 = {view__resp_andMatrixOutputs_andMatrixInput_3_34, view__resp_andMatrixOutputs_andMatrixInput_4_13};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_13 = {view__resp_andMatrixOutputs_andMatrixInput_0_34, view__resp_andMatrixOutputs_andMatrixInput_1_34};
  wire [2:0]  view__resp_andMatrixOutputs_hi_34 = {view__resp_andMatrixOutputs_hi_hi_13, view__resp_andMatrixOutputs_andMatrixInput_2_34};
  wire        view__resp_andMatrixOutputs_2_2_6 = &{view__resp_andMatrixOutputs_hi_34, view__resp_andMatrixOutputs_lo_34};
  wire [1:0]  view__resp_orMatrixOutputs_lo_6 = {view__resp_andMatrixOutputs_0_2_6, view__resp_andMatrixOutputs_2_2_6};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_6 = {view__resp_andMatrixOutputs_4_2_6, view__resp_andMatrixOutputs_1_2_6};
  wire [2:0]  view__resp_orMatrixOutputs_hi_6 = {view__resp_orMatrixOutputs_hi_hi_6, view__resp_andMatrixOutputs_3_2_6};
  wire        view__resp_orMatrixOutputs_6 = |{view__resp_orMatrixOutputs_hi_6, view__resp_orMatrixOutputs_lo_6};
  assign view__resp_invMatrixOutputs_6 = view__resp_orMatrixOutputs_6;
  wire        view__resp_plaOutput_6 = view__resp_invMatrixOutputs_6;
  assign view__resp_plaInput_6 = {1'h0, req_opcode[1:0], req_src_0[6], req_opcode[2] ^ req_src_1[6]};
  wire [4:0]  view__resp_plaInput_7;
  wire [4:0]  view__resp_invInputs_7 = ~view__resp_plaInput_7;
  wire        view__resp_invMatrixOutputs_7;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_35 = view__resp_plaInput_7[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_36 = view__resp_plaInput_7[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_38 = view__resp_plaInput_7[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_35 = view__resp_plaInput_7[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_37 = view__resp_plaInput_7[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_39 = view__resp_plaInput_7[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_35 = view__resp_invInputs_7[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_36 = view__resp_invInputs_7[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_37 = view__resp_invInputs_7[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_35 = view__resp_invInputs_7[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_36 = view__resp_invInputs_7[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_37 = view__resp_invInputs_7[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_14 = view__resp_invInputs_7[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_15 = view__resp_invInputs_7[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_35 = {view__resp_andMatrixOutputs_andMatrixInput_2_35, view__resp_andMatrixOutputs_andMatrixInput_3_35};
  wire [1:0]  view__resp_andMatrixOutputs_hi_35 = {view__resp_andMatrixOutputs_andMatrixInput_0_35, view__resp_andMatrixOutputs_andMatrixInput_1_35};
  wire        view__resp_andMatrixOutputs_4_2_7 = &{view__resp_andMatrixOutputs_hi_35, view__resp_andMatrixOutputs_lo_35};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_36 = view__resp_plaInput_7[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_37 = view__resp_plaInput_7[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_36 = {view__resp_andMatrixOutputs_andMatrixInput_2_36, view__resp_andMatrixOutputs_andMatrixInput_3_36};
  wire [1:0]  view__resp_andMatrixOutputs_hi_36 = {view__resp_andMatrixOutputs_andMatrixInput_0_36, view__resp_andMatrixOutputs_andMatrixInput_1_36};
  wire        view__resp_andMatrixOutputs_1_2_7 = &{view__resp_andMatrixOutputs_hi_36, view__resp_andMatrixOutputs_lo_36};
  wire [1:0]  view__resp_andMatrixOutputs_lo_37 = {view__resp_andMatrixOutputs_andMatrixInput_2_37, view__resp_andMatrixOutputs_andMatrixInput_3_37};
  wire [1:0]  view__resp_andMatrixOutputs_hi_37 = {view__resp_andMatrixOutputs_andMatrixInput_0_37, view__resp_andMatrixOutputs_andMatrixInput_1_37};
  wire        view__resp_andMatrixOutputs_3_2_7 = &{view__resp_andMatrixOutputs_hi_37, view__resp_andMatrixOutputs_lo_37};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_38 = view__resp_invInputs_7[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_38 = view__resp_invInputs_7[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_39 = view__resp_invInputs_7[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_38 = view__resp_plaInput_7[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_39 = view__resp_plaInput_7[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_38 = {view__resp_andMatrixOutputs_andMatrixInput_3_38, view__resp_andMatrixOutputs_andMatrixInput_4_14};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_14 = {view__resp_andMatrixOutputs_andMatrixInput_0_38, view__resp_andMatrixOutputs_andMatrixInput_1_38};
  wire [2:0]  view__resp_andMatrixOutputs_hi_38 = {view__resp_andMatrixOutputs_hi_hi_14, view__resp_andMatrixOutputs_andMatrixInput_2_38};
  wire        view__resp_andMatrixOutputs_0_2_7 = &{view__resp_andMatrixOutputs_hi_38, view__resp_andMatrixOutputs_lo_38};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_39 = view__resp_invInputs_7[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_39 = {view__resp_andMatrixOutputs_andMatrixInput_3_39, view__resp_andMatrixOutputs_andMatrixInput_4_15};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_15 = {view__resp_andMatrixOutputs_andMatrixInput_0_39, view__resp_andMatrixOutputs_andMatrixInput_1_39};
  wire [2:0]  view__resp_andMatrixOutputs_hi_39 = {view__resp_andMatrixOutputs_hi_hi_15, view__resp_andMatrixOutputs_andMatrixInput_2_39};
  wire        view__resp_andMatrixOutputs_2_2_7 = &{view__resp_andMatrixOutputs_hi_39, view__resp_andMatrixOutputs_lo_39};
  wire [1:0]  view__resp_orMatrixOutputs_lo_7 = {view__resp_andMatrixOutputs_0_2_7, view__resp_andMatrixOutputs_2_2_7};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_7 = {view__resp_andMatrixOutputs_4_2_7, view__resp_andMatrixOutputs_1_2_7};
  wire [2:0]  view__resp_orMatrixOutputs_hi_7 = {view__resp_orMatrixOutputs_hi_hi_7, view__resp_andMatrixOutputs_3_2_7};
  wire        view__resp_orMatrixOutputs_7 = |{view__resp_orMatrixOutputs_hi_7, view__resp_orMatrixOutputs_lo_7};
  assign view__resp_invMatrixOutputs_7 = view__resp_orMatrixOutputs_7;
  wire        view__resp_plaOutput_7 = view__resp_invMatrixOutputs_7;
  assign view__resp_plaInput_7 = {1'h0, req_opcode[1:0], req_src_0[7], req_opcode[2] ^ req_src_1[7]};
  wire [4:0]  view__resp_plaInput_8;
  wire [4:0]  view__resp_invInputs_8 = ~view__resp_plaInput_8;
  wire        view__resp_invMatrixOutputs_8;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_40 = view__resp_plaInput_8[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_41 = view__resp_plaInput_8[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_43 = view__resp_plaInput_8[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_40 = view__resp_plaInput_8[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_42 = view__resp_plaInput_8[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_44 = view__resp_plaInput_8[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_40 = view__resp_invInputs_8[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_41 = view__resp_invInputs_8[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_42 = view__resp_invInputs_8[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_40 = view__resp_invInputs_8[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_41 = view__resp_invInputs_8[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_42 = view__resp_invInputs_8[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_16 = view__resp_invInputs_8[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_17 = view__resp_invInputs_8[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_40 = {view__resp_andMatrixOutputs_andMatrixInput_2_40, view__resp_andMatrixOutputs_andMatrixInput_3_40};
  wire [1:0]  view__resp_andMatrixOutputs_hi_40 = {view__resp_andMatrixOutputs_andMatrixInput_0_40, view__resp_andMatrixOutputs_andMatrixInput_1_40};
  wire        view__resp_andMatrixOutputs_4_2_8 = &{view__resp_andMatrixOutputs_hi_40, view__resp_andMatrixOutputs_lo_40};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_41 = view__resp_plaInput_8[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_42 = view__resp_plaInput_8[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_41 = {view__resp_andMatrixOutputs_andMatrixInput_2_41, view__resp_andMatrixOutputs_andMatrixInput_3_41};
  wire [1:0]  view__resp_andMatrixOutputs_hi_41 = {view__resp_andMatrixOutputs_andMatrixInput_0_41, view__resp_andMatrixOutputs_andMatrixInput_1_41};
  wire        view__resp_andMatrixOutputs_1_2_8 = &{view__resp_andMatrixOutputs_hi_41, view__resp_andMatrixOutputs_lo_41};
  wire [1:0]  view__resp_andMatrixOutputs_lo_42 = {view__resp_andMatrixOutputs_andMatrixInput_2_42, view__resp_andMatrixOutputs_andMatrixInput_3_42};
  wire [1:0]  view__resp_andMatrixOutputs_hi_42 = {view__resp_andMatrixOutputs_andMatrixInput_0_42, view__resp_andMatrixOutputs_andMatrixInput_1_42};
  wire        view__resp_andMatrixOutputs_3_2_8 = &{view__resp_andMatrixOutputs_hi_42, view__resp_andMatrixOutputs_lo_42};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_43 = view__resp_invInputs_8[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_43 = view__resp_invInputs_8[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_44 = view__resp_invInputs_8[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_43 = view__resp_plaInput_8[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_44 = view__resp_plaInput_8[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_43 = {view__resp_andMatrixOutputs_andMatrixInput_3_43, view__resp_andMatrixOutputs_andMatrixInput_4_16};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_16 = {view__resp_andMatrixOutputs_andMatrixInput_0_43, view__resp_andMatrixOutputs_andMatrixInput_1_43};
  wire [2:0]  view__resp_andMatrixOutputs_hi_43 = {view__resp_andMatrixOutputs_hi_hi_16, view__resp_andMatrixOutputs_andMatrixInput_2_43};
  wire        view__resp_andMatrixOutputs_0_2_8 = &{view__resp_andMatrixOutputs_hi_43, view__resp_andMatrixOutputs_lo_43};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_44 = view__resp_invInputs_8[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_44 = {view__resp_andMatrixOutputs_andMatrixInput_3_44, view__resp_andMatrixOutputs_andMatrixInput_4_17};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_17 = {view__resp_andMatrixOutputs_andMatrixInput_0_44, view__resp_andMatrixOutputs_andMatrixInput_1_44};
  wire [2:0]  view__resp_andMatrixOutputs_hi_44 = {view__resp_andMatrixOutputs_hi_hi_17, view__resp_andMatrixOutputs_andMatrixInput_2_44};
  wire        view__resp_andMatrixOutputs_2_2_8 = &{view__resp_andMatrixOutputs_hi_44, view__resp_andMatrixOutputs_lo_44};
  wire [1:0]  view__resp_orMatrixOutputs_lo_8 = {view__resp_andMatrixOutputs_0_2_8, view__resp_andMatrixOutputs_2_2_8};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_8 = {view__resp_andMatrixOutputs_4_2_8, view__resp_andMatrixOutputs_1_2_8};
  wire [2:0]  view__resp_orMatrixOutputs_hi_8 = {view__resp_orMatrixOutputs_hi_hi_8, view__resp_andMatrixOutputs_3_2_8};
  wire        view__resp_orMatrixOutputs_8 = |{view__resp_orMatrixOutputs_hi_8, view__resp_orMatrixOutputs_lo_8};
  assign view__resp_invMatrixOutputs_8 = view__resp_orMatrixOutputs_8;
  wire        view__resp_plaOutput_8 = view__resp_invMatrixOutputs_8;
  assign view__resp_plaInput_8 = {1'h0, req_opcode[1:0], req_src_0[8], req_opcode[2] ^ req_src_1[8]};
  wire [4:0]  view__resp_plaInput_9;
  wire [4:0]  view__resp_invInputs_9 = ~view__resp_plaInput_9;
  wire        view__resp_invMatrixOutputs_9;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_45 = view__resp_plaInput_9[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_46 = view__resp_plaInput_9[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_48 = view__resp_plaInput_9[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_45 = view__resp_plaInput_9[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_47 = view__resp_plaInput_9[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_49 = view__resp_plaInput_9[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_45 = view__resp_invInputs_9[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_46 = view__resp_invInputs_9[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_47 = view__resp_invInputs_9[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_45 = view__resp_invInputs_9[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_46 = view__resp_invInputs_9[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_47 = view__resp_invInputs_9[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_18 = view__resp_invInputs_9[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_19 = view__resp_invInputs_9[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_45 = {view__resp_andMatrixOutputs_andMatrixInput_2_45, view__resp_andMatrixOutputs_andMatrixInput_3_45};
  wire [1:0]  view__resp_andMatrixOutputs_hi_45 = {view__resp_andMatrixOutputs_andMatrixInput_0_45, view__resp_andMatrixOutputs_andMatrixInput_1_45};
  wire        view__resp_andMatrixOutputs_4_2_9 = &{view__resp_andMatrixOutputs_hi_45, view__resp_andMatrixOutputs_lo_45};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_46 = view__resp_plaInput_9[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_47 = view__resp_plaInput_9[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_46 = {view__resp_andMatrixOutputs_andMatrixInput_2_46, view__resp_andMatrixOutputs_andMatrixInput_3_46};
  wire [1:0]  view__resp_andMatrixOutputs_hi_46 = {view__resp_andMatrixOutputs_andMatrixInput_0_46, view__resp_andMatrixOutputs_andMatrixInput_1_46};
  wire        view__resp_andMatrixOutputs_1_2_9 = &{view__resp_andMatrixOutputs_hi_46, view__resp_andMatrixOutputs_lo_46};
  wire [1:0]  view__resp_andMatrixOutputs_lo_47 = {view__resp_andMatrixOutputs_andMatrixInput_2_47, view__resp_andMatrixOutputs_andMatrixInput_3_47};
  wire [1:0]  view__resp_andMatrixOutputs_hi_47 = {view__resp_andMatrixOutputs_andMatrixInput_0_47, view__resp_andMatrixOutputs_andMatrixInput_1_47};
  wire        view__resp_andMatrixOutputs_3_2_9 = &{view__resp_andMatrixOutputs_hi_47, view__resp_andMatrixOutputs_lo_47};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_48 = view__resp_invInputs_9[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_48 = view__resp_invInputs_9[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_49 = view__resp_invInputs_9[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_48 = view__resp_plaInput_9[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_49 = view__resp_plaInput_9[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_48 = {view__resp_andMatrixOutputs_andMatrixInput_3_48, view__resp_andMatrixOutputs_andMatrixInput_4_18};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_18 = {view__resp_andMatrixOutputs_andMatrixInput_0_48, view__resp_andMatrixOutputs_andMatrixInput_1_48};
  wire [2:0]  view__resp_andMatrixOutputs_hi_48 = {view__resp_andMatrixOutputs_hi_hi_18, view__resp_andMatrixOutputs_andMatrixInput_2_48};
  wire        view__resp_andMatrixOutputs_0_2_9 = &{view__resp_andMatrixOutputs_hi_48, view__resp_andMatrixOutputs_lo_48};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_49 = view__resp_invInputs_9[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_49 = {view__resp_andMatrixOutputs_andMatrixInput_3_49, view__resp_andMatrixOutputs_andMatrixInput_4_19};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_19 = {view__resp_andMatrixOutputs_andMatrixInput_0_49, view__resp_andMatrixOutputs_andMatrixInput_1_49};
  wire [2:0]  view__resp_andMatrixOutputs_hi_49 = {view__resp_andMatrixOutputs_hi_hi_19, view__resp_andMatrixOutputs_andMatrixInput_2_49};
  wire        view__resp_andMatrixOutputs_2_2_9 = &{view__resp_andMatrixOutputs_hi_49, view__resp_andMatrixOutputs_lo_49};
  wire [1:0]  view__resp_orMatrixOutputs_lo_9 = {view__resp_andMatrixOutputs_0_2_9, view__resp_andMatrixOutputs_2_2_9};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_9 = {view__resp_andMatrixOutputs_4_2_9, view__resp_andMatrixOutputs_1_2_9};
  wire [2:0]  view__resp_orMatrixOutputs_hi_9 = {view__resp_orMatrixOutputs_hi_hi_9, view__resp_andMatrixOutputs_3_2_9};
  wire        view__resp_orMatrixOutputs_9 = |{view__resp_orMatrixOutputs_hi_9, view__resp_orMatrixOutputs_lo_9};
  assign view__resp_invMatrixOutputs_9 = view__resp_orMatrixOutputs_9;
  wire        view__resp_plaOutput_9 = view__resp_invMatrixOutputs_9;
  assign view__resp_plaInput_9 = {1'h0, req_opcode[1:0], req_src_0[9], req_opcode[2] ^ req_src_1[9]};
  wire [4:0]  view__resp_plaInput_10;
  wire [4:0]  view__resp_invInputs_10 = ~view__resp_plaInput_10;
  wire        view__resp_invMatrixOutputs_10;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_50 = view__resp_plaInput_10[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_51 = view__resp_plaInput_10[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_53 = view__resp_plaInput_10[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_50 = view__resp_plaInput_10[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_52 = view__resp_plaInput_10[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_54 = view__resp_plaInput_10[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_50 = view__resp_invInputs_10[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_51 = view__resp_invInputs_10[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_52 = view__resp_invInputs_10[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_50 = view__resp_invInputs_10[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_51 = view__resp_invInputs_10[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_52 = view__resp_invInputs_10[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_20 = view__resp_invInputs_10[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_21 = view__resp_invInputs_10[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_50 = {view__resp_andMatrixOutputs_andMatrixInput_2_50, view__resp_andMatrixOutputs_andMatrixInput_3_50};
  wire [1:0]  view__resp_andMatrixOutputs_hi_50 = {view__resp_andMatrixOutputs_andMatrixInput_0_50, view__resp_andMatrixOutputs_andMatrixInput_1_50};
  wire        view__resp_andMatrixOutputs_4_2_10 = &{view__resp_andMatrixOutputs_hi_50, view__resp_andMatrixOutputs_lo_50};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_51 = view__resp_plaInput_10[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_52 = view__resp_plaInput_10[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_51 = {view__resp_andMatrixOutputs_andMatrixInput_2_51, view__resp_andMatrixOutputs_andMatrixInput_3_51};
  wire [1:0]  view__resp_andMatrixOutputs_hi_51 = {view__resp_andMatrixOutputs_andMatrixInput_0_51, view__resp_andMatrixOutputs_andMatrixInput_1_51};
  wire        view__resp_andMatrixOutputs_1_2_10 = &{view__resp_andMatrixOutputs_hi_51, view__resp_andMatrixOutputs_lo_51};
  wire [1:0]  view__resp_andMatrixOutputs_lo_52 = {view__resp_andMatrixOutputs_andMatrixInput_2_52, view__resp_andMatrixOutputs_andMatrixInput_3_52};
  wire [1:0]  view__resp_andMatrixOutputs_hi_52 = {view__resp_andMatrixOutputs_andMatrixInput_0_52, view__resp_andMatrixOutputs_andMatrixInput_1_52};
  wire        view__resp_andMatrixOutputs_3_2_10 = &{view__resp_andMatrixOutputs_hi_52, view__resp_andMatrixOutputs_lo_52};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_53 = view__resp_invInputs_10[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_53 = view__resp_invInputs_10[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_54 = view__resp_invInputs_10[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_53 = view__resp_plaInput_10[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_54 = view__resp_plaInput_10[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_53 = {view__resp_andMatrixOutputs_andMatrixInput_3_53, view__resp_andMatrixOutputs_andMatrixInput_4_20};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_20 = {view__resp_andMatrixOutputs_andMatrixInput_0_53, view__resp_andMatrixOutputs_andMatrixInput_1_53};
  wire [2:0]  view__resp_andMatrixOutputs_hi_53 = {view__resp_andMatrixOutputs_hi_hi_20, view__resp_andMatrixOutputs_andMatrixInput_2_53};
  wire        view__resp_andMatrixOutputs_0_2_10 = &{view__resp_andMatrixOutputs_hi_53, view__resp_andMatrixOutputs_lo_53};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_54 = view__resp_invInputs_10[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_54 = {view__resp_andMatrixOutputs_andMatrixInput_3_54, view__resp_andMatrixOutputs_andMatrixInput_4_21};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_21 = {view__resp_andMatrixOutputs_andMatrixInput_0_54, view__resp_andMatrixOutputs_andMatrixInput_1_54};
  wire [2:0]  view__resp_andMatrixOutputs_hi_54 = {view__resp_andMatrixOutputs_hi_hi_21, view__resp_andMatrixOutputs_andMatrixInput_2_54};
  wire        view__resp_andMatrixOutputs_2_2_10 = &{view__resp_andMatrixOutputs_hi_54, view__resp_andMatrixOutputs_lo_54};
  wire [1:0]  view__resp_orMatrixOutputs_lo_10 = {view__resp_andMatrixOutputs_0_2_10, view__resp_andMatrixOutputs_2_2_10};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_10 = {view__resp_andMatrixOutputs_4_2_10, view__resp_andMatrixOutputs_1_2_10};
  wire [2:0]  view__resp_orMatrixOutputs_hi_10 = {view__resp_orMatrixOutputs_hi_hi_10, view__resp_andMatrixOutputs_3_2_10};
  wire        view__resp_orMatrixOutputs_10 = |{view__resp_orMatrixOutputs_hi_10, view__resp_orMatrixOutputs_lo_10};
  assign view__resp_invMatrixOutputs_10 = view__resp_orMatrixOutputs_10;
  wire        view__resp_plaOutput_10 = view__resp_invMatrixOutputs_10;
  assign view__resp_plaInput_10 = {1'h0, req_opcode[1:0], req_src_0[10], req_opcode[2] ^ req_src_1[10]};
  wire [4:0]  view__resp_plaInput_11;
  wire [4:0]  view__resp_invInputs_11 = ~view__resp_plaInput_11;
  wire        view__resp_invMatrixOutputs_11;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_55 = view__resp_plaInput_11[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_56 = view__resp_plaInput_11[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_58 = view__resp_plaInput_11[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_55 = view__resp_plaInput_11[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_57 = view__resp_plaInput_11[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_59 = view__resp_plaInput_11[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_55 = view__resp_invInputs_11[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_56 = view__resp_invInputs_11[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_57 = view__resp_invInputs_11[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_55 = view__resp_invInputs_11[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_56 = view__resp_invInputs_11[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_57 = view__resp_invInputs_11[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_22 = view__resp_invInputs_11[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_23 = view__resp_invInputs_11[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_55 = {view__resp_andMatrixOutputs_andMatrixInput_2_55, view__resp_andMatrixOutputs_andMatrixInput_3_55};
  wire [1:0]  view__resp_andMatrixOutputs_hi_55 = {view__resp_andMatrixOutputs_andMatrixInput_0_55, view__resp_andMatrixOutputs_andMatrixInput_1_55};
  wire        view__resp_andMatrixOutputs_4_2_11 = &{view__resp_andMatrixOutputs_hi_55, view__resp_andMatrixOutputs_lo_55};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_56 = view__resp_plaInput_11[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_57 = view__resp_plaInput_11[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_56 = {view__resp_andMatrixOutputs_andMatrixInput_2_56, view__resp_andMatrixOutputs_andMatrixInput_3_56};
  wire [1:0]  view__resp_andMatrixOutputs_hi_56 = {view__resp_andMatrixOutputs_andMatrixInput_0_56, view__resp_andMatrixOutputs_andMatrixInput_1_56};
  wire        view__resp_andMatrixOutputs_1_2_11 = &{view__resp_andMatrixOutputs_hi_56, view__resp_andMatrixOutputs_lo_56};
  wire [1:0]  view__resp_andMatrixOutputs_lo_57 = {view__resp_andMatrixOutputs_andMatrixInput_2_57, view__resp_andMatrixOutputs_andMatrixInput_3_57};
  wire [1:0]  view__resp_andMatrixOutputs_hi_57 = {view__resp_andMatrixOutputs_andMatrixInput_0_57, view__resp_andMatrixOutputs_andMatrixInput_1_57};
  wire        view__resp_andMatrixOutputs_3_2_11 = &{view__resp_andMatrixOutputs_hi_57, view__resp_andMatrixOutputs_lo_57};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_58 = view__resp_invInputs_11[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_58 = view__resp_invInputs_11[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_59 = view__resp_invInputs_11[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_58 = view__resp_plaInput_11[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_59 = view__resp_plaInput_11[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_58 = {view__resp_andMatrixOutputs_andMatrixInput_3_58, view__resp_andMatrixOutputs_andMatrixInput_4_22};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_22 = {view__resp_andMatrixOutputs_andMatrixInput_0_58, view__resp_andMatrixOutputs_andMatrixInput_1_58};
  wire [2:0]  view__resp_andMatrixOutputs_hi_58 = {view__resp_andMatrixOutputs_hi_hi_22, view__resp_andMatrixOutputs_andMatrixInput_2_58};
  wire        view__resp_andMatrixOutputs_0_2_11 = &{view__resp_andMatrixOutputs_hi_58, view__resp_andMatrixOutputs_lo_58};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_59 = view__resp_invInputs_11[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_59 = {view__resp_andMatrixOutputs_andMatrixInput_3_59, view__resp_andMatrixOutputs_andMatrixInput_4_23};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_23 = {view__resp_andMatrixOutputs_andMatrixInput_0_59, view__resp_andMatrixOutputs_andMatrixInput_1_59};
  wire [2:0]  view__resp_andMatrixOutputs_hi_59 = {view__resp_andMatrixOutputs_hi_hi_23, view__resp_andMatrixOutputs_andMatrixInput_2_59};
  wire        view__resp_andMatrixOutputs_2_2_11 = &{view__resp_andMatrixOutputs_hi_59, view__resp_andMatrixOutputs_lo_59};
  wire [1:0]  view__resp_orMatrixOutputs_lo_11 = {view__resp_andMatrixOutputs_0_2_11, view__resp_andMatrixOutputs_2_2_11};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_11 = {view__resp_andMatrixOutputs_4_2_11, view__resp_andMatrixOutputs_1_2_11};
  wire [2:0]  view__resp_orMatrixOutputs_hi_11 = {view__resp_orMatrixOutputs_hi_hi_11, view__resp_andMatrixOutputs_3_2_11};
  wire        view__resp_orMatrixOutputs_11 = |{view__resp_orMatrixOutputs_hi_11, view__resp_orMatrixOutputs_lo_11};
  assign view__resp_invMatrixOutputs_11 = view__resp_orMatrixOutputs_11;
  wire        view__resp_plaOutput_11 = view__resp_invMatrixOutputs_11;
  assign view__resp_plaInput_11 = {1'h0, req_opcode[1:0], req_src_0[11], req_opcode[2] ^ req_src_1[11]};
  wire [4:0]  view__resp_plaInput_12;
  wire [4:0]  view__resp_invInputs_12 = ~view__resp_plaInput_12;
  wire        view__resp_invMatrixOutputs_12;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_60 = view__resp_plaInput_12[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_61 = view__resp_plaInput_12[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_63 = view__resp_plaInput_12[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_60 = view__resp_plaInput_12[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_62 = view__resp_plaInput_12[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_64 = view__resp_plaInput_12[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_60 = view__resp_invInputs_12[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_61 = view__resp_invInputs_12[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_62 = view__resp_invInputs_12[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_60 = view__resp_invInputs_12[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_61 = view__resp_invInputs_12[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_62 = view__resp_invInputs_12[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_24 = view__resp_invInputs_12[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_25 = view__resp_invInputs_12[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_60 = {view__resp_andMatrixOutputs_andMatrixInput_2_60, view__resp_andMatrixOutputs_andMatrixInput_3_60};
  wire [1:0]  view__resp_andMatrixOutputs_hi_60 = {view__resp_andMatrixOutputs_andMatrixInput_0_60, view__resp_andMatrixOutputs_andMatrixInput_1_60};
  wire        view__resp_andMatrixOutputs_4_2_12 = &{view__resp_andMatrixOutputs_hi_60, view__resp_andMatrixOutputs_lo_60};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_61 = view__resp_plaInput_12[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_62 = view__resp_plaInput_12[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_61 = {view__resp_andMatrixOutputs_andMatrixInput_2_61, view__resp_andMatrixOutputs_andMatrixInput_3_61};
  wire [1:0]  view__resp_andMatrixOutputs_hi_61 = {view__resp_andMatrixOutputs_andMatrixInput_0_61, view__resp_andMatrixOutputs_andMatrixInput_1_61};
  wire        view__resp_andMatrixOutputs_1_2_12 = &{view__resp_andMatrixOutputs_hi_61, view__resp_andMatrixOutputs_lo_61};
  wire [1:0]  view__resp_andMatrixOutputs_lo_62 = {view__resp_andMatrixOutputs_andMatrixInput_2_62, view__resp_andMatrixOutputs_andMatrixInput_3_62};
  wire [1:0]  view__resp_andMatrixOutputs_hi_62 = {view__resp_andMatrixOutputs_andMatrixInput_0_62, view__resp_andMatrixOutputs_andMatrixInput_1_62};
  wire        view__resp_andMatrixOutputs_3_2_12 = &{view__resp_andMatrixOutputs_hi_62, view__resp_andMatrixOutputs_lo_62};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_63 = view__resp_invInputs_12[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_63 = view__resp_invInputs_12[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_64 = view__resp_invInputs_12[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_63 = view__resp_plaInput_12[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_64 = view__resp_plaInput_12[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_63 = {view__resp_andMatrixOutputs_andMatrixInput_3_63, view__resp_andMatrixOutputs_andMatrixInput_4_24};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_24 = {view__resp_andMatrixOutputs_andMatrixInput_0_63, view__resp_andMatrixOutputs_andMatrixInput_1_63};
  wire [2:0]  view__resp_andMatrixOutputs_hi_63 = {view__resp_andMatrixOutputs_hi_hi_24, view__resp_andMatrixOutputs_andMatrixInput_2_63};
  wire        view__resp_andMatrixOutputs_0_2_12 = &{view__resp_andMatrixOutputs_hi_63, view__resp_andMatrixOutputs_lo_63};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_64 = view__resp_invInputs_12[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_64 = {view__resp_andMatrixOutputs_andMatrixInput_3_64, view__resp_andMatrixOutputs_andMatrixInput_4_25};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_25 = {view__resp_andMatrixOutputs_andMatrixInput_0_64, view__resp_andMatrixOutputs_andMatrixInput_1_64};
  wire [2:0]  view__resp_andMatrixOutputs_hi_64 = {view__resp_andMatrixOutputs_hi_hi_25, view__resp_andMatrixOutputs_andMatrixInput_2_64};
  wire        view__resp_andMatrixOutputs_2_2_12 = &{view__resp_andMatrixOutputs_hi_64, view__resp_andMatrixOutputs_lo_64};
  wire [1:0]  view__resp_orMatrixOutputs_lo_12 = {view__resp_andMatrixOutputs_0_2_12, view__resp_andMatrixOutputs_2_2_12};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_12 = {view__resp_andMatrixOutputs_4_2_12, view__resp_andMatrixOutputs_1_2_12};
  wire [2:0]  view__resp_orMatrixOutputs_hi_12 = {view__resp_orMatrixOutputs_hi_hi_12, view__resp_andMatrixOutputs_3_2_12};
  wire        view__resp_orMatrixOutputs_12 = |{view__resp_orMatrixOutputs_hi_12, view__resp_orMatrixOutputs_lo_12};
  assign view__resp_invMatrixOutputs_12 = view__resp_orMatrixOutputs_12;
  wire        view__resp_plaOutput_12 = view__resp_invMatrixOutputs_12;
  assign view__resp_plaInput_12 = {1'h0, req_opcode[1:0], req_src_0[12], req_opcode[2] ^ req_src_1[12]};
  wire [4:0]  view__resp_plaInput_13;
  wire [4:0]  view__resp_invInputs_13 = ~view__resp_plaInput_13;
  wire        view__resp_invMatrixOutputs_13;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_65 = view__resp_plaInput_13[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_66 = view__resp_plaInput_13[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_68 = view__resp_plaInput_13[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_65 = view__resp_plaInput_13[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_67 = view__resp_plaInput_13[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_69 = view__resp_plaInput_13[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_65 = view__resp_invInputs_13[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_66 = view__resp_invInputs_13[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_67 = view__resp_invInputs_13[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_65 = view__resp_invInputs_13[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_66 = view__resp_invInputs_13[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_67 = view__resp_invInputs_13[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_26 = view__resp_invInputs_13[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_27 = view__resp_invInputs_13[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_65 = {view__resp_andMatrixOutputs_andMatrixInput_2_65, view__resp_andMatrixOutputs_andMatrixInput_3_65};
  wire [1:0]  view__resp_andMatrixOutputs_hi_65 = {view__resp_andMatrixOutputs_andMatrixInput_0_65, view__resp_andMatrixOutputs_andMatrixInput_1_65};
  wire        view__resp_andMatrixOutputs_4_2_13 = &{view__resp_andMatrixOutputs_hi_65, view__resp_andMatrixOutputs_lo_65};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_66 = view__resp_plaInput_13[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_67 = view__resp_plaInput_13[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_66 = {view__resp_andMatrixOutputs_andMatrixInput_2_66, view__resp_andMatrixOutputs_andMatrixInput_3_66};
  wire [1:0]  view__resp_andMatrixOutputs_hi_66 = {view__resp_andMatrixOutputs_andMatrixInput_0_66, view__resp_andMatrixOutputs_andMatrixInput_1_66};
  wire        view__resp_andMatrixOutputs_1_2_13 = &{view__resp_andMatrixOutputs_hi_66, view__resp_andMatrixOutputs_lo_66};
  wire [1:0]  view__resp_andMatrixOutputs_lo_67 = {view__resp_andMatrixOutputs_andMatrixInput_2_67, view__resp_andMatrixOutputs_andMatrixInput_3_67};
  wire [1:0]  view__resp_andMatrixOutputs_hi_67 = {view__resp_andMatrixOutputs_andMatrixInput_0_67, view__resp_andMatrixOutputs_andMatrixInput_1_67};
  wire        view__resp_andMatrixOutputs_3_2_13 = &{view__resp_andMatrixOutputs_hi_67, view__resp_andMatrixOutputs_lo_67};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_68 = view__resp_invInputs_13[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_68 = view__resp_invInputs_13[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_69 = view__resp_invInputs_13[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_68 = view__resp_plaInput_13[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_69 = view__resp_plaInput_13[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_68 = {view__resp_andMatrixOutputs_andMatrixInput_3_68, view__resp_andMatrixOutputs_andMatrixInput_4_26};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_26 = {view__resp_andMatrixOutputs_andMatrixInput_0_68, view__resp_andMatrixOutputs_andMatrixInput_1_68};
  wire [2:0]  view__resp_andMatrixOutputs_hi_68 = {view__resp_andMatrixOutputs_hi_hi_26, view__resp_andMatrixOutputs_andMatrixInput_2_68};
  wire        view__resp_andMatrixOutputs_0_2_13 = &{view__resp_andMatrixOutputs_hi_68, view__resp_andMatrixOutputs_lo_68};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_69 = view__resp_invInputs_13[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_69 = {view__resp_andMatrixOutputs_andMatrixInput_3_69, view__resp_andMatrixOutputs_andMatrixInput_4_27};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_27 = {view__resp_andMatrixOutputs_andMatrixInput_0_69, view__resp_andMatrixOutputs_andMatrixInput_1_69};
  wire [2:0]  view__resp_andMatrixOutputs_hi_69 = {view__resp_andMatrixOutputs_hi_hi_27, view__resp_andMatrixOutputs_andMatrixInput_2_69};
  wire        view__resp_andMatrixOutputs_2_2_13 = &{view__resp_andMatrixOutputs_hi_69, view__resp_andMatrixOutputs_lo_69};
  wire [1:0]  view__resp_orMatrixOutputs_lo_13 = {view__resp_andMatrixOutputs_0_2_13, view__resp_andMatrixOutputs_2_2_13};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_13 = {view__resp_andMatrixOutputs_4_2_13, view__resp_andMatrixOutputs_1_2_13};
  wire [2:0]  view__resp_orMatrixOutputs_hi_13 = {view__resp_orMatrixOutputs_hi_hi_13, view__resp_andMatrixOutputs_3_2_13};
  wire        view__resp_orMatrixOutputs_13 = |{view__resp_orMatrixOutputs_hi_13, view__resp_orMatrixOutputs_lo_13};
  assign view__resp_invMatrixOutputs_13 = view__resp_orMatrixOutputs_13;
  wire        view__resp_plaOutput_13 = view__resp_invMatrixOutputs_13;
  assign view__resp_plaInput_13 = {1'h0, req_opcode[1:0], req_src_0[13], req_opcode[2] ^ req_src_1[13]};
  wire [4:0]  view__resp_plaInput_14;
  wire [4:0]  view__resp_invInputs_14 = ~view__resp_plaInput_14;
  wire        view__resp_invMatrixOutputs_14;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_70 = view__resp_plaInput_14[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_71 = view__resp_plaInput_14[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_73 = view__resp_plaInput_14[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_70 = view__resp_plaInput_14[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_72 = view__resp_plaInput_14[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_74 = view__resp_plaInput_14[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_70 = view__resp_invInputs_14[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_71 = view__resp_invInputs_14[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_72 = view__resp_invInputs_14[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_70 = view__resp_invInputs_14[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_71 = view__resp_invInputs_14[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_72 = view__resp_invInputs_14[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_28 = view__resp_invInputs_14[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_29 = view__resp_invInputs_14[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_70 = {view__resp_andMatrixOutputs_andMatrixInput_2_70, view__resp_andMatrixOutputs_andMatrixInput_3_70};
  wire [1:0]  view__resp_andMatrixOutputs_hi_70 = {view__resp_andMatrixOutputs_andMatrixInput_0_70, view__resp_andMatrixOutputs_andMatrixInput_1_70};
  wire        view__resp_andMatrixOutputs_4_2_14 = &{view__resp_andMatrixOutputs_hi_70, view__resp_andMatrixOutputs_lo_70};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_71 = view__resp_plaInput_14[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_72 = view__resp_plaInput_14[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_71 = {view__resp_andMatrixOutputs_andMatrixInput_2_71, view__resp_andMatrixOutputs_andMatrixInput_3_71};
  wire [1:0]  view__resp_andMatrixOutputs_hi_71 = {view__resp_andMatrixOutputs_andMatrixInput_0_71, view__resp_andMatrixOutputs_andMatrixInput_1_71};
  wire        view__resp_andMatrixOutputs_1_2_14 = &{view__resp_andMatrixOutputs_hi_71, view__resp_andMatrixOutputs_lo_71};
  wire [1:0]  view__resp_andMatrixOutputs_lo_72 = {view__resp_andMatrixOutputs_andMatrixInput_2_72, view__resp_andMatrixOutputs_andMatrixInput_3_72};
  wire [1:0]  view__resp_andMatrixOutputs_hi_72 = {view__resp_andMatrixOutputs_andMatrixInput_0_72, view__resp_andMatrixOutputs_andMatrixInput_1_72};
  wire        view__resp_andMatrixOutputs_3_2_14 = &{view__resp_andMatrixOutputs_hi_72, view__resp_andMatrixOutputs_lo_72};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_73 = view__resp_invInputs_14[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_73 = view__resp_invInputs_14[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_74 = view__resp_invInputs_14[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_73 = view__resp_plaInput_14[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_74 = view__resp_plaInput_14[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_73 = {view__resp_andMatrixOutputs_andMatrixInput_3_73, view__resp_andMatrixOutputs_andMatrixInput_4_28};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_28 = {view__resp_andMatrixOutputs_andMatrixInput_0_73, view__resp_andMatrixOutputs_andMatrixInput_1_73};
  wire [2:0]  view__resp_andMatrixOutputs_hi_73 = {view__resp_andMatrixOutputs_hi_hi_28, view__resp_andMatrixOutputs_andMatrixInput_2_73};
  wire        view__resp_andMatrixOutputs_0_2_14 = &{view__resp_andMatrixOutputs_hi_73, view__resp_andMatrixOutputs_lo_73};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_74 = view__resp_invInputs_14[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_74 = {view__resp_andMatrixOutputs_andMatrixInput_3_74, view__resp_andMatrixOutputs_andMatrixInput_4_29};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_29 = {view__resp_andMatrixOutputs_andMatrixInput_0_74, view__resp_andMatrixOutputs_andMatrixInput_1_74};
  wire [2:0]  view__resp_andMatrixOutputs_hi_74 = {view__resp_andMatrixOutputs_hi_hi_29, view__resp_andMatrixOutputs_andMatrixInput_2_74};
  wire        view__resp_andMatrixOutputs_2_2_14 = &{view__resp_andMatrixOutputs_hi_74, view__resp_andMatrixOutputs_lo_74};
  wire [1:0]  view__resp_orMatrixOutputs_lo_14 = {view__resp_andMatrixOutputs_0_2_14, view__resp_andMatrixOutputs_2_2_14};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_14 = {view__resp_andMatrixOutputs_4_2_14, view__resp_andMatrixOutputs_1_2_14};
  wire [2:0]  view__resp_orMatrixOutputs_hi_14 = {view__resp_orMatrixOutputs_hi_hi_14, view__resp_andMatrixOutputs_3_2_14};
  wire        view__resp_orMatrixOutputs_14 = |{view__resp_orMatrixOutputs_hi_14, view__resp_orMatrixOutputs_lo_14};
  assign view__resp_invMatrixOutputs_14 = view__resp_orMatrixOutputs_14;
  wire        view__resp_plaOutput_14 = view__resp_invMatrixOutputs_14;
  assign view__resp_plaInput_14 = {1'h0, req_opcode[1:0], req_src_0[14], req_opcode[2] ^ req_src_1[14]};
  wire [4:0]  view__resp_plaInput_15;
  wire [4:0]  view__resp_invInputs_15 = ~view__resp_plaInput_15;
  wire        view__resp_invMatrixOutputs_15;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_75 = view__resp_plaInput_15[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_76 = view__resp_plaInput_15[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_78 = view__resp_plaInput_15[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_75 = view__resp_plaInput_15[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_77 = view__resp_plaInput_15[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_79 = view__resp_plaInput_15[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_75 = view__resp_invInputs_15[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_76 = view__resp_invInputs_15[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_77 = view__resp_invInputs_15[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_75 = view__resp_invInputs_15[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_76 = view__resp_invInputs_15[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_77 = view__resp_invInputs_15[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_30 = view__resp_invInputs_15[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_31 = view__resp_invInputs_15[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_75 = {view__resp_andMatrixOutputs_andMatrixInput_2_75, view__resp_andMatrixOutputs_andMatrixInput_3_75};
  wire [1:0]  view__resp_andMatrixOutputs_hi_75 = {view__resp_andMatrixOutputs_andMatrixInput_0_75, view__resp_andMatrixOutputs_andMatrixInput_1_75};
  wire        view__resp_andMatrixOutputs_4_2_15 = &{view__resp_andMatrixOutputs_hi_75, view__resp_andMatrixOutputs_lo_75};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_76 = view__resp_plaInput_15[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_77 = view__resp_plaInput_15[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_76 = {view__resp_andMatrixOutputs_andMatrixInput_2_76, view__resp_andMatrixOutputs_andMatrixInput_3_76};
  wire [1:0]  view__resp_andMatrixOutputs_hi_76 = {view__resp_andMatrixOutputs_andMatrixInput_0_76, view__resp_andMatrixOutputs_andMatrixInput_1_76};
  wire        view__resp_andMatrixOutputs_1_2_15 = &{view__resp_andMatrixOutputs_hi_76, view__resp_andMatrixOutputs_lo_76};
  wire [1:0]  view__resp_andMatrixOutputs_lo_77 = {view__resp_andMatrixOutputs_andMatrixInput_2_77, view__resp_andMatrixOutputs_andMatrixInput_3_77};
  wire [1:0]  view__resp_andMatrixOutputs_hi_77 = {view__resp_andMatrixOutputs_andMatrixInput_0_77, view__resp_andMatrixOutputs_andMatrixInput_1_77};
  wire        view__resp_andMatrixOutputs_3_2_15 = &{view__resp_andMatrixOutputs_hi_77, view__resp_andMatrixOutputs_lo_77};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_78 = view__resp_invInputs_15[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_78 = view__resp_invInputs_15[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_79 = view__resp_invInputs_15[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_78 = view__resp_plaInput_15[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_79 = view__resp_plaInput_15[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_78 = {view__resp_andMatrixOutputs_andMatrixInput_3_78, view__resp_andMatrixOutputs_andMatrixInput_4_30};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_30 = {view__resp_andMatrixOutputs_andMatrixInput_0_78, view__resp_andMatrixOutputs_andMatrixInput_1_78};
  wire [2:0]  view__resp_andMatrixOutputs_hi_78 = {view__resp_andMatrixOutputs_hi_hi_30, view__resp_andMatrixOutputs_andMatrixInput_2_78};
  wire        view__resp_andMatrixOutputs_0_2_15 = &{view__resp_andMatrixOutputs_hi_78, view__resp_andMatrixOutputs_lo_78};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_79 = view__resp_invInputs_15[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_79 = {view__resp_andMatrixOutputs_andMatrixInput_3_79, view__resp_andMatrixOutputs_andMatrixInput_4_31};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_31 = {view__resp_andMatrixOutputs_andMatrixInput_0_79, view__resp_andMatrixOutputs_andMatrixInput_1_79};
  wire [2:0]  view__resp_andMatrixOutputs_hi_79 = {view__resp_andMatrixOutputs_hi_hi_31, view__resp_andMatrixOutputs_andMatrixInput_2_79};
  wire        view__resp_andMatrixOutputs_2_2_15 = &{view__resp_andMatrixOutputs_hi_79, view__resp_andMatrixOutputs_lo_79};
  wire [1:0]  view__resp_orMatrixOutputs_lo_15 = {view__resp_andMatrixOutputs_0_2_15, view__resp_andMatrixOutputs_2_2_15};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_15 = {view__resp_andMatrixOutputs_4_2_15, view__resp_andMatrixOutputs_1_2_15};
  wire [2:0]  view__resp_orMatrixOutputs_hi_15 = {view__resp_orMatrixOutputs_hi_hi_15, view__resp_andMatrixOutputs_3_2_15};
  wire        view__resp_orMatrixOutputs_15 = |{view__resp_orMatrixOutputs_hi_15, view__resp_orMatrixOutputs_lo_15};
  assign view__resp_invMatrixOutputs_15 = view__resp_orMatrixOutputs_15;
  wire        view__resp_plaOutput_15 = view__resp_invMatrixOutputs_15;
  assign view__resp_plaInput_15 = {1'h0, req_opcode[1:0], req_src_0[15], req_opcode[2] ^ req_src_1[15]};
  wire [4:0]  view__resp_plaInput_16;
  wire [4:0]  view__resp_invInputs_16 = ~view__resp_plaInput_16;
  wire        view__resp_invMatrixOutputs_16;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_80 = view__resp_plaInput_16[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_81 = view__resp_plaInput_16[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_83 = view__resp_plaInput_16[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_80 = view__resp_plaInput_16[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_82 = view__resp_plaInput_16[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_84 = view__resp_plaInput_16[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_80 = view__resp_invInputs_16[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_81 = view__resp_invInputs_16[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_82 = view__resp_invInputs_16[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_80 = view__resp_invInputs_16[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_81 = view__resp_invInputs_16[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_82 = view__resp_invInputs_16[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_32 = view__resp_invInputs_16[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_33 = view__resp_invInputs_16[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_80 = {view__resp_andMatrixOutputs_andMatrixInput_2_80, view__resp_andMatrixOutputs_andMatrixInput_3_80};
  wire [1:0]  view__resp_andMatrixOutputs_hi_80 = {view__resp_andMatrixOutputs_andMatrixInput_0_80, view__resp_andMatrixOutputs_andMatrixInput_1_80};
  wire        view__resp_andMatrixOutputs_4_2_16 = &{view__resp_andMatrixOutputs_hi_80, view__resp_andMatrixOutputs_lo_80};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_81 = view__resp_plaInput_16[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_82 = view__resp_plaInput_16[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_81 = {view__resp_andMatrixOutputs_andMatrixInput_2_81, view__resp_andMatrixOutputs_andMatrixInput_3_81};
  wire [1:0]  view__resp_andMatrixOutputs_hi_81 = {view__resp_andMatrixOutputs_andMatrixInput_0_81, view__resp_andMatrixOutputs_andMatrixInput_1_81};
  wire        view__resp_andMatrixOutputs_1_2_16 = &{view__resp_andMatrixOutputs_hi_81, view__resp_andMatrixOutputs_lo_81};
  wire [1:0]  view__resp_andMatrixOutputs_lo_82 = {view__resp_andMatrixOutputs_andMatrixInput_2_82, view__resp_andMatrixOutputs_andMatrixInput_3_82};
  wire [1:0]  view__resp_andMatrixOutputs_hi_82 = {view__resp_andMatrixOutputs_andMatrixInput_0_82, view__resp_andMatrixOutputs_andMatrixInput_1_82};
  wire        view__resp_andMatrixOutputs_3_2_16 = &{view__resp_andMatrixOutputs_hi_82, view__resp_andMatrixOutputs_lo_82};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_83 = view__resp_invInputs_16[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_83 = view__resp_invInputs_16[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_84 = view__resp_invInputs_16[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_83 = view__resp_plaInput_16[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_84 = view__resp_plaInput_16[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_83 = {view__resp_andMatrixOutputs_andMatrixInput_3_83, view__resp_andMatrixOutputs_andMatrixInput_4_32};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_32 = {view__resp_andMatrixOutputs_andMatrixInput_0_83, view__resp_andMatrixOutputs_andMatrixInput_1_83};
  wire [2:0]  view__resp_andMatrixOutputs_hi_83 = {view__resp_andMatrixOutputs_hi_hi_32, view__resp_andMatrixOutputs_andMatrixInput_2_83};
  wire        view__resp_andMatrixOutputs_0_2_16 = &{view__resp_andMatrixOutputs_hi_83, view__resp_andMatrixOutputs_lo_83};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_84 = view__resp_invInputs_16[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_84 = {view__resp_andMatrixOutputs_andMatrixInput_3_84, view__resp_andMatrixOutputs_andMatrixInput_4_33};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_33 = {view__resp_andMatrixOutputs_andMatrixInput_0_84, view__resp_andMatrixOutputs_andMatrixInput_1_84};
  wire [2:0]  view__resp_andMatrixOutputs_hi_84 = {view__resp_andMatrixOutputs_hi_hi_33, view__resp_andMatrixOutputs_andMatrixInput_2_84};
  wire        view__resp_andMatrixOutputs_2_2_16 = &{view__resp_andMatrixOutputs_hi_84, view__resp_andMatrixOutputs_lo_84};
  wire [1:0]  view__resp_orMatrixOutputs_lo_16 = {view__resp_andMatrixOutputs_0_2_16, view__resp_andMatrixOutputs_2_2_16};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_16 = {view__resp_andMatrixOutputs_4_2_16, view__resp_andMatrixOutputs_1_2_16};
  wire [2:0]  view__resp_orMatrixOutputs_hi_16 = {view__resp_orMatrixOutputs_hi_hi_16, view__resp_andMatrixOutputs_3_2_16};
  wire        view__resp_orMatrixOutputs_16 = |{view__resp_orMatrixOutputs_hi_16, view__resp_orMatrixOutputs_lo_16};
  assign view__resp_invMatrixOutputs_16 = view__resp_orMatrixOutputs_16;
  wire        view__resp_plaOutput_16 = view__resp_invMatrixOutputs_16;
  assign view__resp_plaInput_16 = {1'h0, req_opcode[1:0], req_src_0[16], req_opcode[2] ^ req_src_1[16]};
  wire [4:0]  view__resp_plaInput_17;
  wire [4:0]  view__resp_invInputs_17 = ~view__resp_plaInput_17;
  wire        view__resp_invMatrixOutputs_17;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_85 = view__resp_plaInput_17[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_86 = view__resp_plaInput_17[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_88 = view__resp_plaInput_17[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_85 = view__resp_plaInput_17[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_87 = view__resp_plaInput_17[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_89 = view__resp_plaInput_17[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_85 = view__resp_invInputs_17[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_86 = view__resp_invInputs_17[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_87 = view__resp_invInputs_17[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_85 = view__resp_invInputs_17[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_86 = view__resp_invInputs_17[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_87 = view__resp_invInputs_17[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_34 = view__resp_invInputs_17[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_35 = view__resp_invInputs_17[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_85 = {view__resp_andMatrixOutputs_andMatrixInput_2_85, view__resp_andMatrixOutputs_andMatrixInput_3_85};
  wire [1:0]  view__resp_andMatrixOutputs_hi_85 = {view__resp_andMatrixOutputs_andMatrixInput_0_85, view__resp_andMatrixOutputs_andMatrixInput_1_85};
  wire        view__resp_andMatrixOutputs_4_2_17 = &{view__resp_andMatrixOutputs_hi_85, view__resp_andMatrixOutputs_lo_85};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_86 = view__resp_plaInput_17[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_87 = view__resp_plaInput_17[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_86 = {view__resp_andMatrixOutputs_andMatrixInput_2_86, view__resp_andMatrixOutputs_andMatrixInput_3_86};
  wire [1:0]  view__resp_andMatrixOutputs_hi_86 = {view__resp_andMatrixOutputs_andMatrixInput_0_86, view__resp_andMatrixOutputs_andMatrixInput_1_86};
  wire        view__resp_andMatrixOutputs_1_2_17 = &{view__resp_andMatrixOutputs_hi_86, view__resp_andMatrixOutputs_lo_86};
  wire [1:0]  view__resp_andMatrixOutputs_lo_87 = {view__resp_andMatrixOutputs_andMatrixInput_2_87, view__resp_andMatrixOutputs_andMatrixInput_3_87};
  wire [1:0]  view__resp_andMatrixOutputs_hi_87 = {view__resp_andMatrixOutputs_andMatrixInput_0_87, view__resp_andMatrixOutputs_andMatrixInput_1_87};
  wire        view__resp_andMatrixOutputs_3_2_17 = &{view__resp_andMatrixOutputs_hi_87, view__resp_andMatrixOutputs_lo_87};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_88 = view__resp_invInputs_17[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_88 = view__resp_invInputs_17[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_89 = view__resp_invInputs_17[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_88 = view__resp_plaInput_17[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_89 = view__resp_plaInput_17[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_88 = {view__resp_andMatrixOutputs_andMatrixInput_3_88, view__resp_andMatrixOutputs_andMatrixInput_4_34};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_34 = {view__resp_andMatrixOutputs_andMatrixInput_0_88, view__resp_andMatrixOutputs_andMatrixInput_1_88};
  wire [2:0]  view__resp_andMatrixOutputs_hi_88 = {view__resp_andMatrixOutputs_hi_hi_34, view__resp_andMatrixOutputs_andMatrixInput_2_88};
  wire        view__resp_andMatrixOutputs_0_2_17 = &{view__resp_andMatrixOutputs_hi_88, view__resp_andMatrixOutputs_lo_88};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_89 = view__resp_invInputs_17[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_89 = {view__resp_andMatrixOutputs_andMatrixInput_3_89, view__resp_andMatrixOutputs_andMatrixInput_4_35};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_35 = {view__resp_andMatrixOutputs_andMatrixInput_0_89, view__resp_andMatrixOutputs_andMatrixInput_1_89};
  wire [2:0]  view__resp_andMatrixOutputs_hi_89 = {view__resp_andMatrixOutputs_hi_hi_35, view__resp_andMatrixOutputs_andMatrixInput_2_89};
  wire        view__resp_andMatrixOutputs_2_2_17 = &{view__resp_andMatrixOutputs_hi_89, view__resp_andMatrixOutputs_lo_89};
  wire [1:0]  view__resp_orMatrixOutputs_lo_17 = {view__resp_andMatrixOutputs_0_2_17, view__resp_andMatrixOutputs_2_2_17};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_17 = {view__resp_andMatrixOutputs_4_2_17, view__resp_andMatrixOutputs_1_2_17};
  wire [2:0]  view__resp_orMatrixOutputs_hi_17 = {view__resp_orMatrixOutputs_hi_hi_17, view__resp_andMatrixOutputs_3_2_17};
  wire        view__resp_orMatrixOutputs_17 = |{view__resp_orMatrixOutputs_hi_17, view__resp_orMatrixOutputs_lo_17};
  assign view__resp_invMatrixOutputs_17 = view__resp_orMatrixOutputs_17;
  wire        view__resp_plaOutput_17 = view__resp_invMatrixOutputs_17;
  assign view__resp_plaInput_17 = {1'h0, req_opcode[1:0], req_src_0[17], req_opcode[2] ^ req_src_1[17]};
  wire [4:0]  view__resp_plaInput_18;
  wire [4:0]  view__resp_invInputs_18 = ~view__resp_plaInput_18;
  wire        view__resp_invMatrixOutputs_18;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_90 = view__resp_plaInput_18[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_91 = view__resp_plaInput_18[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_93 = view__resp_plaInput_18[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_90 = view__resp_plaInput_18[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_92 = view__resp_plaInput_18[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_94 = view__resp_plaInput_18[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_90 = view__resp_invInputs_18[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_91 = view__resp_invInputs_18[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_92 = view__resp_invInputs_18[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_90 = view__resp_invInputs_18[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_91 = view__resp_invInputs_18[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_92 = view__resp_invInputs_18[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_36 = view__resp_invInputs_18[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_37 = view__resp_invInputs_18[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_90 = {view__resp_andMatrixOutputs_andMatrixInput_2_90, view__resp_andMatrixOutputs_andMatrixInput_3_90};
  wire [1:0]  view__resp_andMatrixOutputs_hi_90 = {view__resp_andMatrixOutputs_andMatrixInput_0_90, view__resp_andMatrixOutputs_andMatrixInput_1_90};
  wire        view__resp_andMatrixOutputs_4_2_18 = &{view__resp_andMatrixOutputs_hi_90, view__resp_andMatrixOutputs_lo_90};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_91 = view__resp_plaInput_18[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_92 = view__resp_plaInput_18[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_91 = {view__resp_andMatrixOutputs_andMatrixInput_2_91, view__resp_andMatrixOutputs_andMatrixInput_3_91};
  wire [1:0]  view__resp_andMatrixOutputs_hi_91 = {view__resp_andMatrixOutputs_andMatrixInput_0_91, view__resp_andMatrixOutputs_andMatrixInput_1_91};
  wire        view__resp_andMatrixOutputs_1_2_18 = &{view__resp_andMatrixOutputs_hi_91, view__resp_andMatrixOutputs_lo_91};
  wire [1:0]  view__resp_andMatrixOutputs_lo_92 = {view__resp_andMatrixOutputs_andMatrixInput_2_92, view__resp_andMatrixOutputs_andMatrixInput_3_92};
  wire [1:0]  view__resp_andMatrixOutputs_hi_92 = {view__resp_andMatrixOutputs_andMatrixInput_0_92, view__resp_andMatrixOutputs_andMatrixInput_1_92};
  wire        view__resp_andMatrixOutputs_3_2_18 = &{view__resp_andMatrixOutputs_hi_92, view__resp_andMatrixOutputs_lo_92};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_93 = view__resp_invInputs_18[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_93 = view__resp_invInputs_18[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_94 = view__resp_invInputs_18[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_93 = view__resp_plaInput_18[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_94 = view__resp_plaInput_18[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_93 = {view__resp_andMatrixOutputs_andMatrixInput_3_93, view__resp_andMatrixOutputs_andMatrixInput_4_36};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_36 = {view__resp_andMatrixOutputs_andMatrixInput_0_93, view__resp_andMatrixOutputs_andMatrixInput_1_93};
  wire [2:0]  view__resp_andMatrixOutputs_hi_93 = {view__resp_andMatrixOutputs_hi_hi_36, view__resp_andMatrixOutputs_andMatrixInput_2_93};
  wire        view__resp_andMatrixOutputs_0_2_18 = &{view__resp_andMatrixOutputs_hi_93, view__resp_andMatrixOutputs_lo_93};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_94 = view__resp_invInputs_18[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_94 = {view__resp_andMatrixOutputs_andMatrixInput_3_94, view__resp_andMatrixOutputs_andMatrixInput_4_37};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_37 = {view__resp_andMatrixOutputs_andMatrixInput_0_94, view__resp_andMatrixOutputs_andMatrixInput_1_94};
  wire [2:0]  view__resp_andMatrixOutputs_hi_94 = {view__resp_andMatrixOutputs_hi_hi_37, view__resp_andMatrixOutputs_andMatrixInput_2_94};
  wire        view__resp_andMatrixOutputs_2_2_18 = &{view__resp_andMatrixOutputs_hi_94, view__resp_andMatrixOutputs_lo_94};
  wire [1:0]  view__resp_orMatrixOutputs_lo_18 = {view__resp_andMatrixOutputs_0_2_18, view__resp_andMatrixOutputs_2_2_18};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_18 = {view__resp_andMatrixOutputs_4_2_18, view__resp_andMatrixOutputs_1_2_18};
  wire [2:0]  view__resp_orMatrixOutputs_hi_18 = {view__resp_orMatrixOutputs_hi_hi_18, view__resp_andMatrixOutputs_3_2_18};
  wire        view__resp_orMatrixOutputs_18 = |{view__resp_orMatrixOutputs_hi_18, view__resp_orMatrixOutputs_lo_18};
  assign view__resp_invMatrixOutputs_18 = view__resp_orMatrixOutputs_18;
  wire        view__resp_plaOutput_18 = view__resp_invMatrixOutputs_18;
  assign view__resp_plaInput_18 = {1'h0, req_opcode[1:0], req_src_0[18], req_opcode[2] ^ req_src_1[18]};
  wire [4:0]  view__resp_plaInput_19;
  wire [4:0]  view__resp_invInputs_19 = ~view__resp_plaInput_19;
  wire        view__resp_invMatrixOutputs_19;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_95 = view__resp_plaInput_19[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_96 = view__resp_plaInput_19[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_98 = view__resp_plaInput_19[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_95 = view__resp_plaInput_19[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_97 = view__resp_plaInput_19[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_99 = view__resp_plaInput_19[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_95 = view__resp_invInputs_19[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_96 = view__resp_invInputs_19[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_97 = view__resp_invInputs_19[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_95 = view__resp_invInputs_19[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_96 = view__resp_invInputs_19[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_97 = view__resp_invInputs_19[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_38 = view__resp_invInputs_19[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_39 = view__resp_invInputs_19[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_95 = {view__resp_andMatrixOutputs_andMatrixInput_2_95, view__resp_andMatrixOutputs_andMatrixInput_3_95};
  wire [1:0]  view__resp_andMatrixOutputs_hi_95 = {view__resp_andMatrixOutputs_andMatrixInput_0_95, view__resp_andMatrixOutputs_andMatrixInput_1_95};
  wire        view__resp_andMatrixOutputs_4_2_19 = &{view__resp_andMatrixOutputs_hi_95, view__resp_andMatrixOutputs_lo_95};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_96 = view__resp_plaInput_19[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_97 = view__resp_plaInput_19[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_96 = {view__resp_andMatrixOutputs_andMatrixInput_2_96, view__resp_andMatrixOutputs_andMatrixInput_3_96};
  wire [1:0]  view__resp_andMatrixOutputs_hi_96 = {view__resp_andMatrixOutputs_andMatrixInput_0_96, view__resp_andMatrixOutputs_andMatrixInput_1_96};
  wire        view__resp_andMatrixOutputs_1_2_19 = &{view__resp_andMatrixOutputs_hi_96, view__resp_andMatrixOutputs_lo_96};
  wire [1:0]  view__resp_andMatrixOutputs_lo_97 = {view__resp_andMatrixOutputs_andMatrixInput_2_97, view__resp_andMatrixOutputs_andMatrixInput_3_97};
  wire [1:0]  view__resp_andMatrixOutputs_hi_97 = {view__resp_andMatrixOutputs_andMatrixInput_0_97, view__resp_andMatrixOutputs_andMatrixInput_1_97};
  wire        view__resp_andMatrixOutputs_3_2_19 = &{view__resp_andMatrixOutputs_hi_97, view__resp_andMatrixOutputs_lo_97};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_98 = view__resp_invInputs_19[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_98 = view__resp_invInputs_19[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_99 = view__resp_invInputs_19[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_98 = view__resp_plaInput_19[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_99 = view__resp_plaInput_19[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_98 = {view__resp_andMatrixOutputs_andMatrixInput_3_98, view__resp_andMatrixOutputs_andMatrixInput_4_38};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_38 = {view__resp_andMatrixOutputs_andMatrixInput_0_98, view__resp_andMatrixOutputs_andMatrixInput_1_98};
  wire [2:0]  view__resp_andMatrixOutputs_hi_98 = {view__resp_andMatrixOutputs_hi_hi_38, view__resp_andMatrixOutputs_andMatrixInput_2_98};
  wire        view__resp_andMatrixOutputs_0_2_19 = &{view__resp_andMatrixOutputs_hi_98, view__resp_andMatrixOutputs_lo_98};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_99 = view__resp_invInputs_19[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_99 = {view__resp_andMatrixOutputs_andMatrixInput_3_99, view__resp_andMatrixOutputs_andMatrixInput_4_39};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_39 = {view__resp_andMatrixOutputs_andMatrixInput_0_99, view__resp_andMatrixOutputs_andMatrixInput_1_99};
  wire [2:0]  view__resp_andMatrixOutputs_hi_99 = {view__resp_andMatrixOutputs_hi_hi_39, view__resp_andMatrixOutputs_andMatrixInput_2_99};
  wire        view__resp_andMatrixOutputs_2_2_19 = &{view__resp_andMatrixOutputs_hi_99, view__resp_andMatrixOutputs_lo_99};
  wire [1:0]  view__resp_orMatrixOutputs_lo_19 = {view__resp_andMatrixOutputs_0_2_19, view__resp_andMatrixOutputs_2_2_19};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_19 = {view__resp_andMatrixOutputs_4_2_19, view__resp_andMatrixOutputs_1_2_19};
  wire [2:0]  view__resp_orMatrixOutputs_hi_19 = {view__resp_orMatrixOutputs_hi_hi_19, view__resp_andMatrixOutputs_3_2_19};
  wire        view__resp_orMatrixOutputs_19 = |{view__resp_orMatrixOutputs_hi_19, view__resp_orMatrixOutputs_lo_19};
  assign view__resp_invMatrixOutputs_19 = view__resp_orMatrixOutputs_19;
  wire        view__resp_plaOutput_19 = view__resp_invMatrixOutputs_19;
  assign view__resp_plaInput_19 = {1'h0, req_opcode[1:0], req_src_0[19], req_opcode[2] ^ req_src_1[19]};
  wire [4:0]  view__resp_plaInput_20;
  wire [4:0]  view__resp_invInputs_20 = ~view__resp_plaInput_20;
  wire        view__resp_invMatrixOutputs_20;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_100 = view__resp_plaInput_20[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_101 = view__resp_plaInput_20[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_103 = view__resp_plaInput_20[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_100 = view__resp_plaInput_20[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_102 = view__resp_plaInput_20[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_104 = view__resp_plaInput_20[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_100 = view__resp_invInputs_20[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_101 = view__resp_invInputs_20[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_102 = view__resp_invInputs_20[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_100 = view__resp_invInputs_20[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_101 = view__resp_invInputs_20[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_102 = view__resp_invInputs_20[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_40 = view__resp_invInputs_20[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_41 = view__resp_invInputs_20[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_100 = {view__resp_andMatrixOutputs_andMatrixInput_2_100, view__resp_andMatrixOutputs_andMatrixInput_3_100};
  wire [1:0]  view__resp_andMatrixOutputs_hi_100 = {view__resp_andMatrixOutputs_andMatrixInput_0_100, view__resp_andMatrixOutputs_andMatrixInput_1_100};
  wire        view__resp_andMatrixOutputs_4_2_20 = &{view__resp_andMatrixOutputs_hi_100, view__resp_andMatrixOutputs_lo_100};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_101 = view__resp_plaInput_20[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_102 = view__resp_plaInput_20[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_101 = {view__resp_andMatrixOutputs_andMatrixInput_2_101, view__resp_andMatrixOutputs_andMatrixInput_3_101};
  wire [1:0]  view__resp_andMatrixOutputs_hi_101 = {view__resp_andMatrixOutputs_andMatrixInput_0_101, view__resp_andMatrixOutputs_andMatrixInput_1_101};
  wire        view__resp_andMatrixOutputs_1_2_20 = &{view__resp_andMatrixOutputs_hi_101, view__resp_andMatrixOutputs_lo_101};
  wire [1:0]  view__resp_andMatrixOutputs_lo_102 = {view__resp_andMatrixOutputs_andMatrixInput_2_102, view__resp_andMatrixOutputs_andMatrixInput_3_102};
  wire [1:0]  view__resp_andMatrixOutputs_hi_102 = {view__resp_andMatrixOutputs_andMatrixInput_0_102, view__resp_andMatrixOutputs_andMatrixInput_1_102};
  wire        view__resp_andMatrixOutputs_3_2_20 = &{view__resp_andMatrixOutputs_hi_102, view__resp_andMatrixOutputs_lo_102};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_103 = view__resp_invInputs_20[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_103 = view__resp_invInputs_20[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_104 = view__resp_invInputs_20[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_103 = view__resp_plaInput_20[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_104 = view__resp_plaInput_20[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_103 = {view__resp_andMatrixOutputs_andMatrixInput_3_103, view__resp_andMatrixOutputs_andMatrixInput_4_40};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_40 = {view__resp_andMatrixOutputs_andMatrixInput_0_103, view__resp_andMatrixOutputs_andMatrixInput_1_103};
  wire [2:0]  view__resp_andMatrixOutputs_hi_103 = {view__resp_andMatrixOutputs_hi_hi_40, view__resp_andMatrixOutputs_andMatrixInput_2_103};
  wire        view__resp_andMatrixOutputs_0_2_20 = &{view__resp_andMatrixOutputs_hi_103, view__resp_andMatrixOutputs_lo_103};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_104 = view__resp_invInputs_20[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_104 = {view__resp_andMatrixOutputs_andMatrixInput_3_104, view__resp_andMatrixOutputs_andMatrixInput_4_41};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_41 = {view__resp_andMatrixOutputs_andMatrixInput_0_104, view__resp_andMatrixOutputs_andMatrixInput_1_104};
  wire [2:0]  view__resp_andMatrixOutputs_hi_104 = {view__resp_andMatrixOutputs_hi_hi_41, view__resp_andMatrixOutputs_andMatrixInput_2_104};
  wire        view__resp_andMatrixOutputs_2_2_20 = &{view__resp_andMatrixOutputs_hi_104, view__resp_andMatrixOutputs_lo_104};
  wire [1:0]  view__resp_orMatrixOutputs_lo_20 = {view__resp_andMatrixOutputs_0_2_20, view__resp_andMatrixOutputs_2_2_20};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_20 = {view__resp_andMatrixOutputs_4_2_20, view__resp_andMatrixOutputs_1_2_20};
  wire [2:0]  view__resp_orMatrixOutputs_hi_20 = {view__resp_orMatrixOutputs_hi_hi_20, view__resp_andMatrixOutputs_3_2_20};
  wire        view__resp_orMatrixOutputs_20 = |{view__resp_orMatrixOutputs_hi_20, view__resp_orMatrixOutputs_lo_20};
  assign view__resp_invMatrixOutputs_20 = view__resp_orMatrixOutputs_20;
  wire        view__resp_plaOutput_20 = view__resp_invMatrixOutputs_20;
  assign view__resp_plaInput_20 = {1'h0, req_opcode[1:0], req_src_0[20], req_opcode[2] ^ req_src_1[20]};
  wire [4:0]  view__resp_plaInput_21;
  wire [4:0]  view__resp_invInputs_21 = ~view__resp_plaInput_21;
  wire        view__resp_invMatrixOutputs_21;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_105 = view__resp_plaInput_21[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_106 = view__resp_plaInput_21[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_108 = view__resp_plaInput_21[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_105 = view__resp_plaInput_21[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_107 = view__resp_plaInput_21[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_109 = view__resp_plaInput_21[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_105 = view__resp_invInputs_21[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_106 = view__resp_invInputs_21[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_107 = view__resp_invInputs_21[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_105 = view__resp_invInputs_21[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_106 = view__resp_invInputs_21[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_107 = view__resp_invInputs_21[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_42 = view__resp_invInputs_21[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_43 = view__resp_invInputs_21[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_105 = {view__resp_andMatrixOutputs_andMatrixInput_2_105, view__resp_andMatrixOutputs_andMatrixInput_3_105};
  wire [1:0]  view__resp_andMatrixOutputs_hi_105 = {view__resp_andMatrixOutputs_andMatrixInput_0_105, view__resp_andMatrixOutputs_andMatrixInput_1_105};
  wire        view__resp_andMatrixOutputs_4_2_21 = &{view__resp_andMatrixOutputs_hi_105, view__resp_andMatrixOutputs_lo_105};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_106 = view__resp_plaInput_21[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_107 = view__resp_plaInput_21[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_106 = {view__resp_andMatrixOutputs_andMatrixInput_2_106, view__resp_andMatrixOutputs_andMatrixInput_3_106};
  wire [1:0]  view__resp_andMatrixOutputs_hi_106 = {view__resp_andMatrixOutputs_andMatrixInput_0_106, view__resp_andMatrixOutputs_andMatrixInput_1_106};
  wire        view__resp_andMatrixOutputs_1_2_21 = &{view__resp_andMatrixOutputs_hi_106, view__resp_andMatrixOutputs_lo_106};
  wire [1:0]  view__resp_andMatrixOutputs_lo_107 = {view__resp_andMatrixOutputs_andMatrixInput_2_107, view__resp_andMatrixOutputs_andMatrixInput_3_107};
  wire [1:0]  view__resp_andMatrixOutputs_hi_107 = {view__resp_andMatrixOutputs_andMatrixInput_0_107, view__resp_andMatrixOutputs_andMatrixInput_1_107};
  wire        view__resp_andMatrixOutputs_3_2_21 = &{view__resp_andMatrixOutputs_hi_107, view__resp_andMatrixOutputs_lo_107};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_108 = view__resp_invInputs_21[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_108 = view__resp_invInputs_21[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_109 = view__resp_invInputs_21[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_108 = view__resp_plaInput_21[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_109 = view__resp_plaInput_21[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_108 = {view__resp_andMatrixOutputs_andMatrixInput_3_108, view__resp_andMatrixOutputs_andMatrixInput_4_42};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_42 = {view__resp_andMatrixOutputs_andMatrixInput_0_108, view__resp_andMatrixOutputs_andMatrixInput_1_108};
  wire [2:0]  view__resp_andMatrixOutputs_hi_108 = {view__resp_andMatrixOutputs_hi_hi_42, view__resp_andMatrixOutputs_andMatrixInput_2_108};
  wire        view__resp_andMatrixOutputs_0_2_21 = &{view__resp_andMatrixOutputs_hi_108, view__resp_andMatrixOutputs_lo_108};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_109 = view__resp_invInputs_21[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_109 = {view__resp_andMatrixOutputs_andMatrixInput_3_109, view__resp_andMatrixOutputs_andMatrixInput_4_43};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_43 = {view__resp_andMatrixOutputs_andMatrixInput_0_109, view__resp_andMatrixOutputs_andMatrixInput_1_109};
  wire [2:0]  view__resp_andMatrixOutputs_hi_109 = {view__resp_andMatrixOutputs_hi_hi_43, view__resp_andMatrixOutputs_andMatrixInput_2_109};
  wire        view__resp_andMatrixOutputs_2_2_21 = &{view__resp_andMatrixOutputs_hi_109, view__resp_andMatrixOutputs_lo_109};
  wire [1:0]  view__resp_orMatrixOutputs_lo_21 = {view__resp_andMatrixOutputs_0_2_21, view__resp_andMatrixOutputs_2_2_21};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_21 = {view__resp_andMatrixOutputs_4_2_21, view__resp_andMatrixOutputs_1_2_21};
  wire [2:0]  view__resp_orMatrixOutputs_hi_21 = {view__resp_orMatrixOutputs_hi_hi_21, view__resp_andMatrixOutputs_3_2_21};
  wire        view__resp_orMatrixOutputs_21 = |{view__resp_orMatrixOutputs_hi_21, view__resp_orMatrixOutputs_lo_21};
  assign view__resp_invMatrixOutputs_21 = view__resp_orMatrixOutputs_21;
  wire        view__resp_plaOutput_21 = view__resp_invMatrixOutputs_21;
  assign view__resp_plaInput_21 = {1'h0, req_opcode[1:0], req_src_0[21], req_opcode[2] ^ req_src_1[21]};
  wire [4:0]  view__resp_plaInput_22;
  wire [4:0]  view__resp_invInputs_22 = ~view__resp_plaInput_22;
  wire        view__resp_invMatrixOutputs_22;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_110 = view__resp_plaInput_22[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_111 = view__resp_plaInput_22[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_113 = view__resp_plaInput_22[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_110 = view__resp_plaInput_22[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_112 = view__resp_plaInput_22[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_114 = view__resp_plaInput_22[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_110 = view__resp_invInputs_22[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_111 = view__resp_invInputs_22[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_112 = view__resp_invInputs_22[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_110 = view__resp_invInputs_22[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_111 = view__resp_invInputs_22[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_112 = view__resp_invInputs_22[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_44 = view__resp_invInputs_22[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_45 = view__resp_invInputs_22[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_110 = {view__resp_andMatrixOutputs_andMatrixInput_2_110, view__resp_andMatrixOutputs_andMatrixInput_3_110};
  wire [1:0]  view__resp_andMatrixOutputs_hi_110 = {view__resp_andMatrixOutputs_andMatrixInput_0_110, view__resp_andMatrixOutputs_andMatrixInput_1_110};
  wire        view__resp_andMatrixOutputs_4_2_22 = &{view__resp_andMatrixOutputs_hi_110, view__resp_andMatrixOutputs_lo_110};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_111 = view__resp_plaInput_22[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_112 = view__resp_plaInput_22[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_111 = {view__resp_andMatrixOutputs_andMatrixInput_2_111, view__resp_andMatrixOutputs_andMatrixInput_3_111};
  wire [1:0]  view__resp_andMatrixOutputs_hi_111 = {view__resp_andMatrixOutputs_andMatrixInput_0_111, view__resp_andMatrixOutputs_andMatrixInput_1_111};
  wire        view__resp_andMatrixOutputs_1_2_22 = &{view__resp_andMatrixOutputs_hi_111, view__resp_andMatrixOutputs_lo_111};
  wire [1:0]  view__resp_andMatrixOutputs_lo_112 = {view__resp_andMatrixOutputs_andMatrixInput_2_112, view__resp_andMatrixOutputs_andMatrixInput_3_112};
  wire [1:0]  view__resp_andMatrixOutputs_hi_112 = {view__resp_andMatrixOutputs_andMatrixInput_0_112, view__resp_andMatrixOutputs_andMatrixInput_1_112};
  wire        view__resp_andMatrixOutputs_3_2_22 = &{view__resp_andMatrixOutputs_hi_112, view__resp_andMatrixOutputs_lo_112};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_113 = view__resp_invInputs_22[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_113 = view__resp_invInputs_22[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_114 = view__resp_invInputs_22[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_113 = view__resp_plaInput_22[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_114 = view__resp_plaInput_22[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_113 = {view__resp_andMatrixOutputs_andMatrixInput_3_113, view__resp_andMatrixOutputs_andMatrixInput_4_44};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_44 = {view__resp_andMatrixOutputs_andMatrixInput_0_113, view__resp_andMatrixOutputs_andMatrixInput_1_113};
  wire [2:0]  view__resp_andMatrixOutputs_hi_113 = {view__resp_andMatrixOutputs_hi_hi_44, view__resp_andMatrixOutputs_andMatrixInput_2_113};
  wire        view__resp_andMatrixOutputs_0_2_22 = &{view__resp_andMatrixOutputs_hi_113, view__resp_andMatrixOutputs_lo_113};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_114 = view__resp_invInputs_22[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_114 = {view__resp_andMatrixOutputs_andMatrixInput_3_114, view__resp_andMatrixOutputs_andMatrixInput_4_45};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_45 = {view__resp_andMatrixOutputs_andMatrixInput_0_114, view__resp_andMatrixOutputs_andMatrixInput_1_114};
  wire [2:0]  view__resp_andMatrixOutputs_hi_114 = {view__resp_andMatrixOutputs_hi_hi_45, view__resp_andMatrixOutputs_andMatrixInput_2_114};
  wire        view__resp_andMatrixOutputs_2_2_22 = &{view__resp_andMatrixOutputs_hi_114, view__resp_andMatrixOutputs_lo_114};
  wire [1:0]  view__resp_orMatrixOutputs_lo_22 = {view__resp_andMatrixOutputs_0_2_22, view__resp_andMatrixOutputs_2_2_22};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_22 = {view__resp_andMatrixOutputs_4_2_22, view__resp_andMatrixOutputs_1_2_22};
  wire [2:0]  view__resp_orMatrixOutputs_hi_22 = {view__resp_orMatrixOutputs_hi_hi_22, view__resp_andMatrixOutputs_3_2_22};
  wire        view__resp_orMatrixOutputs_22 = |{view__resp_orMatrixOutputs_hi_22, view__resp_orMatrixOutputs_lo_22};
  assign view__resp_invMatrixOutputs_22 = view__resp_orMatrixOutputs_22;
  wire        view__resp_plaOutput_22 = view__resp_invMatrixOutputs_22;
  assign view__resp_plaInput_22 = {1'h0, req_opcode[1:0], req_src_0[22], req_opcode[2] ^ req_src_1[22]};
  wire [4:0]  view__resp_plaInput_23;
  wire [4:0]  view__resp_invInputs_23 = ~view__resp_plaInput_23;
  wire        view__resp_invMatrixOutputs_23;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_115 = view__resp_plaInput_23[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_116 = view__resp_plaInput_23[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_118 = view__resp_plaInput_23[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_115 = view__resp_plaInput_23[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_117 = view__resp_plaInput_23[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_119 = view__resp_plaInput_23[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_115 = view__resp_invInputs_23[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_116 = view__resp_invInputs_23[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_117 = view__resp_invInputs_23[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_115 = view__resp_invInputs_23[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_116 = view__resp_invInputs_23[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_117 = view__resp_invInputs_23[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_46 = view__resp_invInputs_23[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_47 = view__resp_invInputs_23[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_115 = {view__resp_andMatrixOutputs_andMatrixInput_2_115, view__resp_andMatrixOutputs_andMatrixInput_3_115};
  wire [1:0]  view__resp_andMatrixOutputs_hi_115 = {view__resp_andMatrixOutputs_andMatrixInput_0_115, view__resp_andMatrixOutputs_andMatrixInput_1_115};
  wire        view__resp_andMatrixOutputs_4_2_23 = &{view__resp_andMatrixOutputs_hi_115, view__resp_andMatrixOutputs_lo_115};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_116 = view__resp_plaInput_23[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_117 = view__resp_plaInput_23[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_116 = {view__resp_andMatrixOutputs_andMatrixInput_2_116, view__resp_andMatrixOutputs_andMatrixInput_3_116};
  wire [1:0]  view__resp_andMatrixOutputs_hi_116 = {view__resp_andMatrixOutputs_andMatrixInput_0_116, view__resp_andMatrixOutputs_andMatrixInput_1_116};
  wire        view__resp_andMatrixOutputs_1_2_23 = &{view__resp_andMatrixOutputs_hi_116, view__resp_andMatrixOutputs_lo_116};
  wire [1:0]  view__resp_andMatrixOutputs_lo_117 = {view__resp_andMatrixOutputs_andMatrixInput_2_117, view__resp_andMatrixOutputs_andMatrixInput_3_117};
  wire [1:0]  view__resp_andMatrixOutputs_hi_117 = {view__resp_andMatrixOutputs_andMatrixInput_0_117, view__resp_andMatrixOutputs_andMatrixInput_1_117};
  wire        view__resp_andMatrixOutputs_3_2_23 = &{view__resp_andMatrixOutputs_hi_117, view__resp_andMatrixOutputs_lo_117};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_118 = view__resp_invInputs_23[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_118 = view__resp_invInputs_23[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_119 = view__resp_invInputs_23[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_118 = view__resp_plaInput_23[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_119 = view__resp_plaInput_23[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_118 = {view__resp_andMatrixOutputs_andMatrixInput_3_118, view__resp_andMatrixOutputs_andMatrixInput_4_46};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_46 = {view__resp_andMatrixOutputs_andMatrixInput_0_118, view__resp_andMatrixOutputs_andMatrixInput_1_118};
  wire [2:0]  view__resp_andMatrixOutputs_hi_118 = {view__resp_andMatrixOutputs_hi_hi_46, view__resp_andMatrixOutputs_andMatrixInput_2_118};
  wire        view__resp_andMatrixOutputs_0_2_23 = &{view__resp_andMatrixOutputs_hi_118, view__resp_andMatrixOutputs_lo_118};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_119 = view__resp_invInputs_23[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_119 = {view__resp_andMatrixOutputs_andMatrixInput_3_119, view__resp_andMatrixOutputs_andMatrixInput_4_47};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_47 = {view__resp_andMatrixOutputs_andMatrixInput_0_119, view__resp_andMatrixOutputs_andMatrixInput_1_119};
  wire [2:0]  view__resp_andMatrixOutputs_hi_119 = {view__resp_andMatrixOutputs_hi_hi_47, view__resp_andMatrixOutputs_andMatrixInput_2_119};
  wire        view__resp_andMatrixOutputs_2_2_23 = &{view__resp_andMatrixOutputs_hi_119, view__resp_andMatrixOutputs_lo_119};
  wire [1:0]  view__resp_orMatrixOutputs_lo_23 = {view__resp_andMatrixOutputs_0_2_23, view__resp_andMatrixOutputs_2_2_23};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_23 = {view__resp_andMatrixOutputs_4_2_23, view__resp_andMatrixOutputs_1_2_23};
  wire [2:0]  view__resp_orMatrixOutputs_hi_23 = {view__resp_orMatrixOutputs_hi_hi_23, view__resp_andMatrixOutputs_3_2_23};
  wire        view__resp_orMatrixOutputs_23 = |{view__resp_orMatrixOutputs_hi_23, view__resp_orMatrixOutputs_lo_23};
  assign view__resp_invMatrixOutputs_23 = view__resp_orMatrixOutputs_23;
  wire        view__resp_plaOutput_23 = view__resp_invMatrixOutputs_23;
  assign view__resp_plaInput_23 = {1'h0, req_opcode[1:0], req_src_0[23], req_opcode[2] ^ req_src_1[23]};
  wire [4:0]  view__resp_plaInput_24;
  wire [4:0]  view__resp_invInputs_24 = ~view__resp_plaInput_24;
  wire        view__resp_invMatrixOutputs_24;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_120 = view__resp_plaInput_24[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_121 = view__resp_plaInput_24[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_123 = view__resp_plaInput_24[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_120 = view__resp_plaInput_24[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_122 = view__resp_plaInput_24[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_124 = view__resp_plaInput_24[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_120 = view__resp_invInputs_24[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_121 = view__resp_invInputs_24[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_122 = view__resp_invInputs_24[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_120 = view__resp_invInputs_24[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_121 = view__resp_invInputs_24[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_122 = view__resp_invInputs_24[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_48 = view__resp_invInputs_24[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_49 = view__resp_invInputs_24[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_120 = {view__resp_andMatrixOutputs_andMatrixInput_2_120, view__resp_andMatrixOutputs_andMatrixInput_3_120};
  wire [1:0]  view__resp_andMatrixOutputs_hi_120 = {view__resp_andMatrixOutputs_andMatrixInput_0_120, view__resp_andMatrixOutputs_andMatrixInput_1_120};
  wire        view__resp_andMatrixOutputs_4_2_24 = &{view__resp_andMatrixOutputs_hi_120, view__resp_andMatrixOutputs_lo_120};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_121 = view__resp_plaInput_24[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_122 = view__resp_plaInput_24[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_121 = {view__resp_andMatrixOutputs_andMatrixInput_2_121, view__resp_andMatrixOutputs_andMatrixInput_3_121};
  wire [1:0]  view__resp_andMatrixOutputs_hi_121 = {view__resp_andMatrixOutputs_andMatrixInput_0_121, view__resp_andMatrixOutputs_andMatrixInput_1_121};
  wire        view__resp_andMatrixOutputs_1_2_24 = &{view__resp_andMatrixOutputs_hi_121, view__resp_andMatrixOutputs_lo_121};
  wire [1:0]  view__resp_andMatrixOutputs_lo_122 = {view__resp_andMatrixOutputs_andMatrixInput_2_122, view__resp_andMatrixOutputs_andMatrixInput_3_122};
  wire [1:0]  view__resp_andMatrixOutputs_hi_122 = {view__resp_andMatrixOutputs_andMatrixInput_0_122, view__resp_andMatrixOutputs_andMatrixInput_1_122};
  wire        view__resp_andMatrixOutputs_3_2_24 = &{view__resp_andMatrixOutputs_hi_122, view__resp_andMatrixOutputs_lo_122};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_123 = view__resp_invInputs_24[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_123 = view__resp_invInputs_24[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_124 = view__resp_invInputs_24[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_123 = view__resp_plaInput_24[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_124 = view__resp_plaInput_24[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_123 = {view__resp_andMatrixOutputs_andMatrixInput_3_123, view__resp_andMatrixOutputs_andMatrixInput_4_48};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_48 = {view__resp_andMatrixOutputs_andMatrixInput_0_123, view__resp_andMatrixOutputs_andMatrixInput_1_123};
  wire [2:0]  view__resp_andMatrixOutputs_hi_123 = {view__resp_andMatrixOutputs_hi_hi_48, view__resp_andMatrixOutputs_andMatrixInput_2_123};
  wire        view__resp_andMatrixOutputs_0_2_24 = &{view__resp_andMatrixOutputs_hi_123, view__resp_andMatrixOutputs_lo_123};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_124 = view__resp_invInputs_24[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_124 = {view__resp_andMatrixOutputs_andMatrixInput_3_124, view__resp_andMatrixOutputs_andMatrixInput_4_49};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_49 = {view__resp_andMatrixOutputs_andMatrixInput_0_124, view__resp_andMatrixOutputs_andMatrixInput_1_124};
  wire [2:0]  view__resp_andMatrixOutputs_hi_124 = {view__resp_andMatrixOutputs_hi_hi_49, view__resp_andMatrixOutputs_andMatrixInput_2_124};
  wire        view__resp_andMatrixOutputs_2_2_24 = &{view__resp_andMatrixOutputs_hi_124, view__resp_andMatrixOutputs_lo_124};
  wire [1:0]  view__resp_orMatrixOutputs_lo_24 = {view__resp_andMatrixOutputs_0_2_24, view__resp_andMatrixOutputs_2_2_24};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_24 = {view__resp_andMatrixOutputs_4_2_24, view__resp_andMatrixOutputs_1_2_24};
  wire [2:0]  view__resp_orMatrixOutputs_hi_24 = {view__resp_orMatrixOutputs_hi_hi_24, view__resp_andMatrixOutputs_3_2_24};
  wire        view__resp_orMatrixOutputs_24 = |{view__resp_orMatrixOutputs_hi_24, view__resp_orMatrixOutputs_lo_24};
  assign view__resp_invMatrixOutputs_24 = view__resp_orMatrixOutputs_24;
  wire        view__resp_plaOutput_24 = view__resp_invMatrixOutputs_24;
  assign view__resp_plaInput_24 = {1'h0, req_opcode[1:0], req_src_0[24], req_opcode[2] ^ req_src_1[24]};
  wire [4:0]  view__resp_plaInput_25;
  wire [4:0]  view__resp_invInputs_25 = ~view__resp_plaInput_25;
  wire        view__resp_invMatrixOutputs_25;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_125 = view__resp_plaInput_25[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_126 = view__resp_plaInput_25[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_128 = view__resp_plaInput_25[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_125 = view__resp_plaInput_25[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_127 = view__resp_plaInput_25[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_129 = view__resp_plaInput_25[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_125 = view__resp_invInputs_25[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_126 = view__resp_invInputs_25[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_127 = view__resp_invInputs_25[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_125 = view__resp_invInputs_25[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_126 = view__resp_invInputs_25[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_127 = view__resp_invInputs_25[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_50 = view__resp_invInputs_25[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_51 = view__resp_invInputs_25[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_125 = {view__resp_andMatrixOutputs_andMatrixInput_2_125, view__resp_andMatrixOutputs_andMatrixInput_3_125};
  wire [1:0]  view__resp_andMatrixOutputs_hi_125 = {view__resp_andMatrixOutputs_andMatrixInput_0_125, view__resp_andMatrixOutputs_andMatrixInput_1_125};
  wire        view__resp_andMatrixOutputs_4_2_25 = &{view__resp_andMatrixOutputs_hi_125, view__resp_andMatrixOutputs_lo_125};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_126 = view__resp_plaInput_25[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_127 = view__resp_plaInput_25[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_126 = {view__resp_andMatrixOutputs_andMatrixInput_2_126, view__resp_andMatrixOutputs_andMatrixInput_3_126};
  wire [1:0]  view__resp_andMatrixOutputs_hi_126 = {view__resp_andMatrixOutputs_andMatrixInput_0_126, view__resp_andMatrixOutputs_andMatrixInput_1_126};
  wire        view__resp_andMatrixOutputs_1_2_25 = &{view__resp_andMatrixOutputs_hi_126, view__resp_andMatrixOutputs_lo_126};
  wire [1:0]  view__resp_andMatrixOutputs_lo_127 = {view__resp_andMatrixOutputs_andMatrixInput_2_127, view__resp_andMatrixOutputs_andMatrixInput_3_127};
  wire [1:0]  view__resp_andMatrixOutputs_hi_127 = {view__resp_andMatrixOutputs_andMatrixInput_0_127, view__resp_andMatrixOutputs_andMatrixInput_1_127};
  wire        view__resp_andMatrixOutputs_3_2_25 = &{view__resp_andMatrixOutputs_hi_127, view__resp_andMatrixOutputs_lo_127};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_128 = view__resp_invInputs_25[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_128 = view__resp_invInputs_25[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_129 = view__resp_invInputs_25[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_128 = view__resp_plaInput_25[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_129 = view__resp_plaInput_25[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_128 = {view__resp_andMatrixOutputs_andMatrixInput_3_128, view__resp_andMatrixOutputs_andMatrixInput_4_50};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_50 = {view__resp_andMatrixOutputs_andMatrixInput_0_128, view__resp_andMatrixOutputs_andMatrixInput_1_128};
  wire [2:0]  view__resp_andMatrixOutputs_hi_128 = {view__resp_andMatrixOutputs_hi_hi_50, view__resp_andMatrixOutputs_andMatrixInput_2_128};
  wire        view__resp_andMatrixOutputs_0_2_25 = &{view__resp_andMatrixOutputs_hi_128, view__resp_andMatrixOutputs_lo_128};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_129 = view__resp_invInputs_25[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_129 = {view__resp_andMatrixOutputs_andMatrixInput_3_129, view__resp_andMatrixOutputs_andMatrixInput_4_51};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_51 = {view__resp_andMatrixOutputs_andMatrixInput_0_129, view__resp_andMatrixOutputs_andMatrixInput_1_129};
  wire [2:0]  view__resp_andMatrixOutputs_hi_129 = {view__resp_andMatrixOutputs_hi_hi_51, view__resp_andMatrixOutputs_andMatrixInput_2_129};
  wire        view__resp_andMatrixOutputs_2_2_25 = &{view__resp_andMatrixOutputs_hi_129, view__resp_andMatrixOutputs_lo_129};
  wire [1:0]  view__resp_orMatrixOutputs_lo_25 = {view__resp_andMatrixOutputs_0_2_25, view__resp_andMatrixOutputs_2_2_25};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_25 = {view__resp_andMatrixOutputs_4_2_25, view__resp_andMatrixOutputs_1_2_25};
  wire [2:0]  view__resp_orMatrixOutputs_hi_25 = {view__resp_orMatrixOutputs_hi_hi_25, view__resp_andMatrixOutputs_3_2_25};
  wire        view__resp_orMatrixOutputs_25 = |{view__resp_orMatrixOutputs_hi_25, view__resp_orMatrixOutputs_lo_25};
  assign view__resp_invMatrixOutputs_25 = view__resp_orMatrixOutputs_25;
  wire        view__resp_plaOutput_25 = view__resp_invMatrixOutputs_25;
  assign view__resp_plaInput_25 = {1'h0, req_opcode[1:0], req_src_0[25], req_opcode[2] ^ req_src_1[25]};
  wire [4:0]  view__resp_plaInput_26;
  wire [4:0]  view__resp_invInputs_26 = ~view__resp_plaInput_26;
  wire        view__resp_invMatrixOutputs_26;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_130 = view__resp_plaInput_26[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_131 = view__resp_plaInput_26[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_133 = view__resp_plaInput_26[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_130 = view__resp_plaInput_26[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_132 = view__resp_plaInput_26[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_134 = view__resp_plaInput_26[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_130 = view__resp_invInputs_26[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_131 = view__resp_invInputs_26[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_132 = view__resp_invInputs_26[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_130 = view__resp_invInputs_26[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_131 = view__resp_invInputs_26[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_132 = view__resp_invInputs_26[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_52 = view__resp_invInputs_26[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_53 = view__resp_invInputs_26[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_130 = {view__resp_andMatrixOutputs_andMatrixInput_2_130, view__resp_andMatrixOutputs_andMatrixInput_3_130};
  wire [1:0]  view__resp_andMatrixOutputs_hi_130 = {view__resp_andMatrixOutputs_andMatrixInput_0_130, view__resp_andMatrixOutputs_andMatrixInput_1_130};
  wire        view__resp_andMatrixOutputs_4_2_26 = &{view__resp_andMatrixOutputs_hi_130, view__resp_andMatrixOutputs_lo_130};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_131 = view__resp_plaInput_26[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_132 = view__resp_plaInput_26[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_131 = {view__resp_andMatrixOutputs_andMatrixInput_2_131, view__resp_andMatrixOutputs_andMatrixInput_3_131};
  wire [1:0]  view__resp_andMatrixOutputs_hi_131 = {view__resp_andMatrixOutputs_andMatrixInput_0_131, view__resp_andMatrixOutputs_andMatrixInput_1_131};
  wire        view__resp_andMatrixOutputs_1_2_26 = &{view__resp_andMatrixOutputs_hi_131, view__resp_andMatrixOutputs_lo_131};
  wire [1:0]  view__resp_andMatrixOutputs_lo_132 = {view__resp_andMatrixOutputs_andMatrixInput_2_132, view__resp_andMatrixOutputs_andMatrixInput_3_132};
  wire [1:0]  view__resp_andMatrixOutputs_hi_132 = {view__resp_andMatrixOutputs_andMatrixInput_0_132, view__resp_andMatrixOutputs_andMatrixInput_1_132};
  wire        view__resp_andMatrixOutputs_3_2_26 = &{view__resp_andMatrixOutputs_hi_132, view__resp_andMatrixOutputs_lo_132};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_133 = view__resp_invInputs_26[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_133 = view__resp_invInputs_26[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_134 = view__resp_invInputs_26[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_133 = view__resp_plaInput_26[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_134 = view__resp_plaInput_26[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_133 = {view__resp_andMatrixOutputs_andMatrixInput_3_133, view__resp_andMatrixOutputs_andMatrixInput_4_52};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_52 = {view__resp_andMatrixOutputs_andMatrixInput_0_133, view__resp_andMatrixOutputs_andMatrixInput_1_133};
  wire [2:0]  view__resp_andMatrixOutputs_hi_133 = {view__resp_andMatrixOutputs_hi_hi_52, view__resp_andMatrixOutputs_andMatrixInput_2_133};
  wire        view__resp_andMatrixOutputs_0_2_26 = &{view__resp_andMatrixOutputs_hi_133, view__resp_andMatrixOutputs_lo_133};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_134 = view__resp_invInputs_26[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_134 = {view__resp_andMatrixOutputs_andMatrixInput_3_134, view__resp_andMatrixOutputs_andMatrixInput_4_53};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_53 = {view__resp_andMatrixOutputs_andMatrixInput_0_134, view__resp_andMatrixOutputs_andMatrixInput_1_134};
  wire [2:0]  view__resp_andMatrixOutputs_hi_134 = {view__resp_andMatrixOutputs_hi_hi_53, view__resp_andMatrixOutputs_andMatrixInput_2_134};
  wire        view__resp_andMatrixOutputs_2_2_26 = &{view__resp_andMatrixOutputs_hi_134, view__resp_andMatrixOutputs_lo_134};
  wire [1:0]  view__resp_orMatrixOutputs_lo_26 = {view__resp_andMatrixOutputs_0_2_26, view__resp_andMatrixOutputs_2_2_26};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_26 = {view__resp_andMatrixOutputs_4_2_26, view__resp_andMatrixOutputs_1_2_26};
  wire [2:0]  view__resp_orMatrixOutputs_hi_26 = {view__resp_orMatrixOutputs_hi_hi_26, view__resp_andMatrixOutputs_3_2_26};
  wire        view__resp_orMatrixOutputs_26 = |{view__resp_orMatrixOutputs_hi_26, view__resp_orMatrixOutputs_lo_26};
  assign view__resp_invMatrixOutputs_26 = view__resp_orMatrixOutputs_26;
  wire        view__resp_plaOutput_26 = view__resp_invMatrixOutputs_26;
  assign view__resp_plaInput_26 = {1'h0, req_opcode[1:0], req_src_0[26], req_opcode[2] ^ req_src_1[26]};
  wire [4:0]  view__resp_plaInput_27;
  wire [4:0]  view__resp_invInputs_27 = ~view__resp_plaInput_27;
  wire        view__resp_invMatrixOutputs_27;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_135 = view__resp_plaInput_27[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_136 = view__resp_plaInput_27[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_138 = view__resp_plaInput_27[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_135 = view__resp_plaInput_27[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_137 = view__resp_plaInput_27[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_139 = view__resp_plaInput_27[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_135 = view__resp_invInputs_27[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_136 = view__resp_invInputs_27[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_137 = view__resp_invInputs_27[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_135 = view__resp_invInputs_27[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_136 = view__resp_invInputs_27[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_137 = view__resp_invInputs_27[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_54 = view__resp_invInputs_27[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_55 = view__resp_invInputs_27[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_135 = {view__resp_andMatrixOutputs_andMatrixInput_2_135, view__resp_andMatrixOutputs_andMatrixInput_3_135};
  wire [1:0]  view__resp_andMatrixOutputs_hi_135 = {view__resp_andMatrixOutputs_andMatrixInput_0_135, view__resp_andMatrixOutputs_andMatrixInput_1_135};
  wire        view__resp_andMatrixOutputs_4_2_27 = &{view__resp_andMatrixOutputs_hi_135, view__resp_andMatrixOutputs_lo_135};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_136 = view__resp_plaInput_27[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_137 = view__resp_plaInput_27[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_136 = {view__resp_andMatrixOutputs_andMatrixInput_2_136, view__resp_andMatrixOutputs_andMatrixInput_3_136};
  wire [1:0]  view__resp_andMatrixOutputs_hi_136 = {view__resp_andMatrixOutputs_andMatrixInput_0_136, view__resp_andMatrixOutputs_andMatrixInput_1_136};
  wire        view__resp_andMatrixOutputs_1_2_27 = &{view__resp_andMatrixOutputs_hi_136, view__resp_andMatrixOutputs_lo_136};
  wire [1:0]  view__resp_andMatrixOutputs_lo_137 = {view__resp_andMatrixOutputs_andMatrixInput_2_137, view__resp_andMatrixOutputs_andMatrixInput_3_137};
  wire [1:0]  view__resp_andMatrixOutputs_hi_137 = {view__resp_andMatrixOutputs_andMatrixInput_0_137, view__resp_andMatrixOutputs_andMatrixInput_1_137};
  wire        view__resp_andMatrixOutputs_3_2_27 = &{view__resp_andMatrixOutputs_hi_137, view__resp_andMatrixOutputs_lo_137};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_138 = view__resp_invInputs_27[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_138 = view__resp_invInputs_27[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_139 = view__resp_invInputs_27[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_138 = view__resp_plaInput_27[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_139 = view__resp_plaInput_27[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_138 = {view__resp_andMatrixOutputs_andMatrixInput_3_138, view__resp_andMatrixOutputs_andMatrixInput_4_54};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_54 = {view__resp_andMatrixOutputs_andMatrixInput_0_138, view__resp_andMatrixOutputs_andMatrixInput_1_138};
  wire [2:0]  view__resp_andMatrixOutputs_hi_138 = {view__resp_andMatrixOutputs_hi_hi_54, view__resp_andMatrixOutputs_andMatrixInput_2_138};
  wire        view__resp_andMatrixOutputs_0_2_27 = &{view__resp_andMatrixOutputs_hi_138, view__resp_andMatrixOutputs_lo_138};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_139 = view__resp_invInputs_27[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_139 = {view__resp_andMatrixOutputs_andMatrixInput_3_139, view__resp_andMatrixOutputs_andMatrixInput_4_55};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_55 = {view__resp_andMatrixOutputs_andMatrixInput_0_139, view__resp_andMatrixOutputs_andMatrixInput_1_139};
  wire [2:0]  view__resp_andMatrixOutputs_hi_139 = {view__resp_andMatrixOutputs_hi_hi_55, view__resp_andMatrixOutputs_andMatrixInput_2_139};
  wire        view__resp_andMatrixOutputs_2_2_27 = &{view__resp_andMatrixOutputs_hi_139, view__resp_andMatrixOutputs_lo_139};
  wire [1:0]  view__resp_orMatrixOutputs_lo_27 = {view__resp_andMatrixOutputs_0_2_27, view__resp_andMatrixOutputs_2_2_27};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_27 = {view__resp_andMatrixOutputs_4_2_27, view__resp_andMatrixOutputs_1_2_27};
  wire [2:0]  view__resp_orMatrixOutputs_hi_27 = {view__resp_orMatrixOutputs_hi_hi_27, view__resp_andMatrixOutputs_3_2_27};
  wire        view__resp_orMatrixOutputs_27 = |{view__resp_orMatrixOutputs_hi_27, view__resp_orMatrixOutputs_lo_27};
  assign view__resp_invMatrixOutputs_27 = view__resp_orMatrixOutputs_27;
  wire        view__resp_plaOutput_27 = view__resp_invMatrixOutputs_27;
  assign view__resp_plaInput_27 = {1'h0, req_opcode[1:0], req_src_0[27], req_opcode[2] ^ req_src_1[27]};
  wire [4:0]  view__resp_plaInput_28;
  wire [4:0]  view__resp_invInputs_28 = ~view__resp_plaInput_28;
  wire        view__resp_invMatrixOutputs_28;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_140 = view__resp_plaInput_28[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_141 = view__resp_plaInput_28[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_143 = view__resp_plaInput_28[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_140 = view__resp_plaInput_28[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_142 = view__resp_plaInput_28[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_144 = view__resp_plaInput_28[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_140 = view__resp_invInputs_28[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_141 = view__resp_invInputs_28[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_142 = view__resp_invInputs_28[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_140 = view__resp_invInputs_28[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_141 = view__resp_invInputs_28[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_142 = view__resp_invInputs_28[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_56 = view__resp_invInputs_28[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_57 = view__resp_invInputs_28[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_140 = {view__resp_andMatrixOutputs_andMatrixInput_2_140, view__resp_andMatrixOutputs_andMatrixInput_3_140};
  wire [1:0]  view__resp_andMatrixOutputs_hi_140 = {view__resp_andMatrixOutputs_andMatrixInput_0_140, view__resp_andMatrixOutputs_andMatrixInput_1_140};
  wire        view__resp_andMatrixOutputs_4_2_28 = &{view__resp_andMatrixOutputs_hi_140, view__resp_andMatrixOutputs_lo_140};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_141 = view__resp_plaInput_28[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_142 = view__resp_plaInput_28[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_141 = {view__resp_andMatrixOutputs_andMatrixInput_2_141, view__resp_andMatrixOutputs_andMatrixInput_3_141};
  wire [1:0]  view__resp_andMatrixOutputs_hi_141 = {view__resp_andMatrixOutputs_andMatrixInput_0_141, view__resp_andMatrixOutputs_andMatrixInput_1_141};
  wire        view__resp_andMatrixOutputs_1_2_28 = &{view__resp_andMatrixOutputs_hi_141, view__resp_andMatrixOutputs_lo_141};
  wire [1:0]  view__resp_andMatrixOutputs_lo_142 = {view__resp_andMatrixOutputs_andMatrixInput_2_142, view__resp_andMatrixOutputs_andMatrixInput_3_142};
  wire [1:0]  view__resp_andMatrixOutputs_hi_142 = {view__resp_andMatrixOutputs_andMatrixInput_0_142, view__resp_andMatrixOutputs_andMatrixInput_1_142};
  wire        view__resp_andMatrixOutputs_3_2_28 = &{view__resp_andMatrixOutputs_hi_142, view__resp_andMatrixOutputs_lo_142};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_143 = view__resp_invInputs_28[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_143 = view__resp_invInputs_28[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_144 = view__resp_invInputs_28[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_143 = view__resp_plaInput_28[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_144 = view__resp_plaInput_28[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_143 = {view__resp_andMatrixOutputs_andMatrixInput_3_143, view__resp_andMatrixOutputs_andMatrixInput_4_56};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_56 = {view__resp_andMatrixOutputs_andMatrixInput_0_143, view__resp_andMatrixOutputs_andMatrixInput_1_143};
  wire [2:0]  view__resp_andMatrixOutputs_hi_143 = {view__resp_andMatrixOutputs_hi_hi_56, view__resp_andMatrixOutputs_andMatrixInput_2_143};
  wire        view__resp_andMatrixOutputs_0_2_28 = &{view__resp_andMatrixOutputs_hi_143, view__resp_andMatrixOutputs_lo_143};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_144 = view__resp_invInputs_28[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_144 = {view__resp_andMatrixOutputs_andMatrixInput_3_144, view__resp_andMatrixOutputs_andMatrixInput_4_57};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_57 = {view__resp_andMatrixOutputs_andMatrixInput_0_144, view__resp_andMatrixOutputs_andMatrixInput_1_144};
  wire [2:0]  view__resp_andMatrixOutputs_hi_144 = {view__resp_andMatrixOutputs_hi_hi_57, view__resp_andMatrixOutputs_andMatrixInput_2_144};
  wire        view__resp_andMatrixOutputs_2_2_28 = &{view__resp_andMatrixOutputs_hi_144, view__resp_andMatrixOutputs_lo_144};
  wire [1:0]  view__resp_orMatrixOutputs_lo_28 = {view__resp_andMatrixOutputs_0_2_28, view__resp_andMatrixOutputs_2_2_28};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_28 = {view__resp_andMatrixOutputs_4_2_28, view__resp_andMatrixOutputs_1_2_28};
  wire [2:0]  view__resp_orMatrixOutputs_hi_28 = {view__resp_orMatrixOutputs_hi_hi_28, view__resp_andMatrixOutputs_3_2_28};
  wire        view__resp_orMatrixOutputs_28 = |{view__resp_orMatrixOutputs_hi_28, view__resp_orMatrixOutputs_lo_28};
  assign view__resp_invMatrixOutputs_28 = view__resp_orMatrixOutputs_28;
  wire        view__resp_plaOutput_28 = view__resp_invMatrixOutputs_28;
  assign view__resp_plaInput_28 = {1'h0, req_opcode[1:0], req_src_0[28], req_opcode[2] ^ req_src_1[28]};
  wire [4:0]  view__resp_plaInput_29;
  wire [4:0]  view__resp_invInputs_29 = ~view__resp_plaInput_29;
  wire        view__resp_invMatrixOutputs_29;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_145 = view__resp_plaInput_29[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_146 = view__resp_plaInput_29[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_148 = view__resp_plaInput_29[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_145 = view__resp_plaInput_29[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_147 = view__resp_plaInput_29[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_149 = view__resp_plaInput_29[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_145 = view__resp_invInputs_29[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_146 = view__resp_invInputs_29[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_147 = view__resp_invInputs_29[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_145 = view__resp_invInputs_29[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_146 = view__resp_invInputs_29[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_147 = view__resp_invInputs_29[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_58 = view__resp_invInputs_29[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_59 = view__resp_invInputs_29[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_145 = {view__resp_andMatrixOutputs_andMatrixInput_2_145, view__resp_andMatrixOutputs_andMatrixInput_3_145};
  wire [1:0]  view__resp_andMatrixOutputs_hi_145 = {view__resp_andMatrixOutputs_andMatrixInput_0_145, view__resp_andMatrixOutputs_andMatrixInput_1_145};
  wire        view__resp_andMatrixOutputs_4_2_29 = &{view__resp_andMatrixOutputs_hi_145, view__resp_andMatrixOutputs_lo_145};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_146 = view__resp_plaInput_29[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_147 = view__resp_plaInput_29[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_146 = {view__resp_andMatrixOutputs_andMatrixInput_2_146, view__resp_andMatrixOutputs_andMatrixInput_3_146};
  wire [1:0]  view__resp_andMatrixOutputs_hi_146 = {view__resp_andMatrixOutputs_andMatrixInput_0_146, view__resp_andMatrixOutputs_andMatrixInput_1_146};
  wire        view__resp_andMatrixOutputs_1_2_29 = &{view__resp_andMatrixOutputs_hi_146, view__resp_andMatrixOutputs_lo_146};
  wire [1:0]  view__resp_andMatrixOutputs_lo_147 = {view__resp_andMatrixOutputs_andMatrixInput_2_147, view__resp_andMatrixOutputs_andMatrixInput_3_147};
  wire [1:0]  view__resp_andMatrixOutputs_hi_147 = {view__resp_andMatrixOutputs_andMatrixInput_0_147, view__resp_andMatrixOutputs_andMatrixInput_1_147};
  wire        view__resp_andMatrixOutputs_3_2_29 = &{view__resp_andMatrixOutputs_hi_147, view__resp_andMatrixOutputs_lo_147};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_148 = view__resp_invInputs_29[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_148 = view__resp_invInputs_29[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_149 = view__resp_invInputs_29[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_148 = view__resp_plaInput_29[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_149 = view__resp_plaInput_29[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_148 = {view__resp_andMatrixOutputs_andMatrixInput_3_148, view__resp_andMatrixOutputs_andMatrixInput_4_58};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_58 = {view__resp_andMatrixOutputs_andMatrixInput_0_148, view__resp_andMatrixOutputs_andMatrixInput_1_148};
  wire [2:0]  view__resp_andMatrixOutputs_hi_148 = {view__resp_andMatrixOutputs_hi_hi_58, view__resp_andMatrixOutputs_andMatrixInput_2_148};
  wire        view__resp_andMatrixOutputs_0_2_29 = &{view__resp_andMatrixOutputs_hi_148, view__resp_andMatrixOutputs_lo_148};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_149 = view__resp_invInputs_29[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_149 = {view__resp_andMatrixOutputs_andMatrixInput_3_149, view__resp_andMatrixOutputs_andMatrixInput_4_59};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_59 = {view__resp_andMatrixOutputs_andMatrixInput_0_149, view__resp_andMatrixOutputs_andMatrixInput_1_149};
  wire [2:0]  view__resp_andMatrixOutputs_hi_149 = {view__resp_andMatrixOutputs_hi_hi_59, view__resp_andMatrixOutputs_andMatrixInput_2_149};
  wire        view__resp_andMatrixOutputs_2_2_29 = &{view__resp_andMatrixOutputs_hi_149, view__resp_andMatrixOutputs_lo_149};
  wire [1:0]  view__resp_orMatrixOutputs_lo_29 = {view__resp_andMatrixOutputs_0_2_29, view__resp_andMatrixOutputs_2_2_29};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_29 = {view__resp_andMatrixOutputs_4_2_29, view__resp_andMatrixOutputs_1_2_29};
  wire [2:0]  view__resp_orMatrixOutputs_hi_29 = {view__resp_orMatrixOutputs_hi_hi_29, view__resp_andMatrixOutputs_3_2_29};
  wire        view__resp_orMatrixOutputs_29 = |{view__resp_orMatrixOutputs_hi_29, view__resp_orMatrixOutputs_lo_29};
  assign view__resp_invMatrixOutputs_29 = view__resp_orMatrixOutputs_29;
  wire        view__resp_plaOutput_29 = view__resp_invMatrixOutputs_29;
  assign view__resp_plaInput_29 = {1'h0, req_opcode[1:0], req_src_0[29], req_opcode[2] ^ req_src_1[29]};
  wire [4:0]  view__resp_plaInput_30;
  wire [4:0]  view__resp_invInputs_30 = ~view__resp_plaInput_30;
  wire        view__resp_invMatrixOutputs_30;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_150 = view__resp_plaInput_30[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_151 = view__resp_plaInput_30[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_153 = view__resp_plaInput_30[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_150 = view__resp_plaInput_30[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_152 = view__resp_plaInput_30[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_154 = view__resp_plaInput_30[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_150 = view__resp_invInputs_30[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_151 = view__resp_invInputs_30[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_152 = view__resp_invInputs_30[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_150 = view__resp_invInputs_30[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_151 = view__resp_invInputs_30[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_152 = view__resp_invInputs_30[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_60 = view__resp_invInputs_30[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_61 = view__resp_invInputs_30[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_150 = {view__resp_andMatrixOutputs_andMatrixInput_2_150, view__resp_andMatrixOutputs_andMatrixInput_3_150};
  wire [1:0]  view__resp_andMatrixOutputs_hi_150 = {view__resp_andMatrixOutputs_andMatrixInput_0_150, view__resp_andMatrixOutputs_andMatrixInput_1_150};
  wire        view__resp_andMatrixOutputs_4_2_30 = &{view__resp_andMatrixOutputs_hi_150, view__resp_andMatrixOutputs_lo_150};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_151 = view__resp_plaInput_30[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_152 = view__resp_plaInput_30[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_151 = {view__resp_andMatrixOutputs_andMatrixInput_2_151, view__resp_andMatrixOutputs_andMatrixInput_3_151};
  wire [1:0]  view__resp_andMatrixOutputs_hi_151 = {view__resp_andMatrixOutputs_andMatrixInput_0_151, view__resp_andMatrixOutputs_andMatrixInput_1_151};
  wire        view__resp_andMatrixOutputs_1_2_30 = &{view__resp_andMatrixOutputs_hi_151, view__resp_andMatrixOutputs_lo_151};
  wire [1:0]  view__resp_andMatrixOutputs_lo_152 = {view__resp_andMatrixOutputs_andMatrixInput_2_152, view__resp_andMatrixOutputs_andMatrixInput_3_152};
  wire [1:0]  view__resp_andMatrixOutputs_hi_152 = {view__resp_andMatrixOutputs_andMatrixInput_0_152, view__resp_andMatrixOutputs_andMatrixInput_1_152};
  wire        view__resp_andMatrixOutputs_3_2_30 = &{view__resp_andMatrixOutputs_hi_152, view__resp_andMatrixOutputs_lo_152};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_153 = view__resp_invInputs_30[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_153 = view__resp_invInputs_30[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_154 = view__resp_invInputs_30[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_153 = view__resp_plaInput_30[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_154 = view__resp_plaInput_30[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_153 = {view__resp_andMatrixOutputs_andMatrixInput_3_153, view__resp_andMatrixOutputs_andMatrixInput_4_60};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_60 = {view__resp_andMatrixOutputs_andMatrixInput_0_153, view__resp_andMatrixOutputs_andMatrixInput_1_153};
  wire [2:0]  view__resp_andMatrixOutputs_hi_153 = {view__resp_andMatrixOutputs_hi_hi_60, view__resp_andMatrixOutputs_andMatrixInput_2_153};
  wire        view__resp_andMatrixOutputs_0_2_30 = &{view__resp_andMatrixOutputs_hi_153, view__resp_andMatrixOutputs_lo_153};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_154 = view__resp_invInputs_30[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_154 = {view__resp_andMatrixOutputs_andMatrixInput_3_154, view__resp_andMatrixOutputs_andMatrixInput_4_61};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_61 = {view__resp_andMatrixOutputs_andMatrixInput_0_154, view__resp_andMatrixOutputs_andMatrixInput_1_154};
  wire [2:0]  view__resp_andMatrixOutputs_hi_154 = {view__resp_andMatrixOutputs_hi_hi_61, view__resp_andMatrixOutputs_andMatrixInput_2_154};
  wire        view__resp_andMatrixOutputs_2_2_30 = &{view__resp_andMatrixOutputs_hi_154, view__resp_andMatrixOutputs_lo_154};
  wire [1:0]  view__resp_orMatrixOutputs_lo_30 = {view__resp_andMatrixOutputs_0_2_30, view__resp_andMatrixOutputs_2_2_30};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_30 = {view__resp_andMatrixOutputs_4_2_30, view__resp_andMatrixOutputs_1_2_30};
  wire [2:0]  view__resp_orMatrixOutputs_hi_30 = {view__resp_orMatrixOutputs_hi_hi_30, view__resp_andMatrixOutputs_3_2_30};
  wire        view__resp_orMatrixOutputs_30 = |{view__resp_orMatrixOutputs_hi_30, view__resp_orMatrixOutputs_lo_30};
  assign view__resp_invMatrixOutputs_30 = view__resp_orMatrixOutputs_30;
  wire        view__resp_plaOutput_30 = view__resp_invMatrixOutputs_30;
  assign view__resp_plaInput_30 = {1'h0, req_opcode[1:0], req_src_0[30], req_opcode[2] ^ req_src_1[30]};
  wire [4:0]  view__resp_plaInput_31;
  wire [4:0]  view__resp_invInputs_31 = ~view__resp_plaInput_31;
  wire        view__resp_invMatrixOutputs_31;
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_155 = view__resp_plaInput_31[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_156 = view__resp_plaInput_31[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_158 = view__resp_plaInput_31[0];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_155 = view__resp_plaInput_31[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_157 = view__resp_plaInput_31[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_159 = view__resp_plaInput_31[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_155 = view__resp_invInputs_31[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_156 = view__resp_invInputs_31[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_157 = view__resp_invInputs_31[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_155 = view__resp_invInputs_31[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_156 = view__resp_invInputs_31[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_157 = view__resp_invInputs_31[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_62 = view__resp_invInputs_31[4];
  wire        view__resp_andMatrixOutputs_andMatrixInput_4_63 = view__resp_invInputs_31[4];
  wire [1:0]  view__resp_andMatrixOutputs_lo_155 = {view__resp_andMatrixOutputs_andMatrixInput_2_155, view__resp_andMatrixOutputs_andMatrixInput_3_155};
  wire [1:0]  view__resp_andMatrixOutputs_hi_155 = {view__resp_andMatrixOutputs_andMatrixInput_0_155, view__resp_andMatrixOutputs_andMatrixInput_1_155};
  wire        view__resp_andMatrixOutputs_4_2_31 = &{view__resp_andMatrixOutputs_hi_155, view__resp_andMatrixOutputs_lo_155};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_156 = view__resp_plaInput_31[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_157 = view__resp_plaInput_31[2];
  wire [1:0]  view__resp_andMatrixOutputs_lo_156 = {view__resp_andMatrixOutputs_andMatrixInput_2_156, view__resp_andMatrixOutputs_andMatrixInput_3_156};
  wire [1:0]  view__resp_andMatrixOutputs_hi_156 = {view__resp_andMatrixOutputs_andMatrixInput_0_156, view__resp_andMatrixOutputs_andMatrixInput_1_156};
  wire        view__resp_andMatrixOutputs_1_2_31 = &{view__resp_andMatrixOutputs_hi_156, view__resp_andMatrixOutputs_lo_156};
  wire [1:0]  view__resp_andMatrixOutputs_lo_157 = {view__resp_andMatrixOutputs_andMatrixInput_2_157, view__resp_andMatrixOutputs_andMatrixInput_3_157};
  wire [1:0]  view__resp_andMatrixOutputs_hi_157 = {view__resp_andMatrixOutputs_andMatrixInput_0_157, view__resp_andMatrixOutputs_andMatrixInput_1_157};
  wire        view__resp_andMatrixOutputs_3_2_31 = &{view__resp_andMatrixOutputs_hi_157, view__resp_andMatrixOutputs_lo_157};
  wire        view__resp_andMatrixOutputs_andMatrixInput_1_158 = view__resp_invInputs_31[1];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_158 = view__resp_invInputs_31[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_2_159 = view__resp_invInputs_31[2];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_158 = view__resp_plaInput_31[3];
  wire        view__resp_andMatrixOutputs_andMatrixInput_3_159 = view__resp_plaInput_31[3];
  wire [1:0]  view__resp_andMatrixOutputs_lo_158 = {view__resp_andMatrixOutputs_andMatrixInput_3_158, view__resp_andMatrixOutputs_andMatrixInput_4_62};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_62 = {view__resp_andMatrixOutputs_andMatrixInput_0_158, view__resp_andMatrixOutputs_andMatrixInput_1_158};
  wire [2:0]  view__resp_andMatrixOutputs_hi_158 = {view__resp_andMatrixOutputs_hi_hi_62, view__resp_andMatrixOutputs_andMatrixInput_2_158};
  wire        view__resp_andMatrixOutputs_0_2_31 = &{view__resp_andMatrixOutputs_hi_158, view__resp_andMatrixOutputs_lo_158};
  wire        view__resp_andMatrixOutputs_andMatrixInput_0_159 = view__resp_invInputs_31[0];
  wire [1:0]  view__resp_andMatrixOutputs_lo_159 = {view__resp_andMatrixOutputs_andMatrixInput_3_159, view__resp_andMatrixOutputs_andMatrixInput_4_63};
  wire [1:0]  view__resp_andMatrixOutputs_hi_hi_63 = {view__resp_andMatrixOutputs_andMatrixInput_0_159, view__resp_andMatrixOutputs_andMatrixInput_1_159};
  wire [2:0]  view__resp_andMatrixOutputs_hi_159 = {view__resp_andMatrixOutputs_hi_hi_63, view__resp_andMatrixOutputs_andMatrixInput_2_159};
  wire        view__resp_andMatrixOutputs_2_2_31 = &{view__resp_andMatrixOutputs_hi_159, view__resp_andMatrixOutputs_lo_159};
  wire [1:0]  view__resp_orMatrixOutputs_lo_31 = {view__resp_andMatrixOutputs_0_2_31, view__resp_andMatrixOutputs_2_2_31};
  wire [1:0]  view__resp_orMatrixOutputs_hi_hi_31 = {view__resp_andMatrixOutputs_4_2_31, view__resp_andMatrixOutputs_1_2_31};
  wire [2:0]  view__resp_orMatrixOutputs_hi_31 = {view__resp_orMatrixOutputs_hi_hi_31, view__resp_andMatrixOutputs_3_2_31};
  wire        view__resp_orMatrixOutputs_31 = |{view__resp_orMatrixOutputs_hi_31, view__resp_orMatrixOutputs_lo_31};
  assign view__resp_invMatrixOutputs_31 = view__resp_orMatrixOutputs_31;
  wire        view__resp_plaOutput_31 = view__resp_invMatrixOutputs_31;
  assign view__resp_plaInput_31 = {1'h0, req_opcode[1:0], req_src_0[31], req_opcode[2] ^ req_src_1[31]};
  wire [1:0]  view__resp_lo_lo_lo_lo = {view__resp_plaOutput_1 ^ req_opcode[3], view__resp_plaOutput ^ req_opcode[3]};
  wire [1:0]  view__resp_lo_lo_lo_hi = {view__resp_plaOutput_3 ^ req_opcode[3], view__resp_plaOutput_2 ^ req_opcode[3]};
  wire [3:0]  view__resp_lo_lo_lo = {view__resp_lo_lo_lo_hi, view__resp_lo_lo_lo_lo};
  wire [1:0]  view__resp_lo_lo_hi_lo = {view__resp_plaOutput_5 ^ req_opcode[3], view__resp_plaOutput_4 ^ req_opcode[3]};
  wire [1:0]  view__resp_lo_lo_hi_hi = {view__resp_plaOutput_7 ^ req_opcode[3], view__resp_plaOutput_6 ^ req_opcode[3]};
  wire [3:0]  view__resp_lo_lo_hi = {view__resp_lo_lo_hi_hi, view__resp_lo_lo_hi_lo};
  wire [7:0]  view__resp_lo_lo = {view__resp_lo_lo_hi, view__resp_lo_lo_lo};
  wire [1:0]  view__resp_lo_hi_lo_lo = {view__resp_plaOutput_9 ^ req_opcode[3], view__resp_plaOutput_8 ^ req_opcode[3]};
  wire [1:0]  view__resp_lo_hi_lo_hi = {view__resp_plaOutput_11 ^ req_opcode[3], view__resp_plaOutput_10 ^ req_opcode[3]};
  wire [3:0]  view__resp_lo_hi_lo = {view__resp_lo_hi_lo_hi, view__resp_lo_hi_lo_lo};
  wire [1:0]  view__resp_lo_hi_hi_lo = {view__resp_plaOutput_13 ^ req_opcode[3], view__resp_plaOutput_12 ^ req_opcode[3]};
  wire [1:0]  view__resp_lo_hi_hi_hi = {view__resp_plaOutput_15 ^ req_opcode[3], view__resp_plaOutput_14 ^ req_opcode[3]};
  wire [3:0]  view__resp_lo_hi_hi = {view__resp_lo_hi_hi_hi, view__resp_lo_hi_hi_lo};
  wire [7:0]  view__resp_lo_hi = {view__resp_lo_hi_hi, view__resp_lo_hi_lo};
  wire [15:0] view__resp_lo = {view__resp_lo_hi, view__resp_lo_lo};
  wire [1:0]  view__resp_hi_lo_lo_lo = {view__resp_plaOutput_17 ^ req_opcode[3], view__resp_plaOutput_16 ^ req_opcode[3]};
  wire [1:0]  view__resp_hi_lo_lo_hi = {view__resp_plaOutput_19 ^ req_opcode[3], view__resp_plaOutput_18 ^ req_opcode[3]};
  wire [3:0]  view__resp_hi_lo_lo = {view__resp_hi_lo_lo_hi, view__resp_hi_lo_lo_lo};
  wire [1:0]  view__resp_hi_lo_hi_lo = {view__resp_plaOutput_21 ^ req_opcode[3], view__resp_plaOutput_20 ^ req_opcode[3]};
  wire [1:0]  view__resp_hi_lo_hi_hi = {view__resp_plaOutput_23 ^ req_opcode[3], view__resp_plaOutput_22 ^ req_opcode[3]};
  wire [3:0]  view__resp_hi_lo_hi = {view__resp_hi_lo_hi_hi, view__resp_hi_lo_hi_lo};
  wire [7:0]  view__resp_hi_lo = {view__resp_hi_lo_hi, view__resp_hi_lo_lo};
  wire [1:0]  view__resp_hi_hi_lo_lo = {view__resp_plaOutput_25 ^ req_opcode[3], view__resp_plaOutput_24 ^ req_opcode[3]};
  wire [1:0]  view__resp_hi_hi_lo_hi = {view__resp_plaOutput_27 ^ req_opcode[3], view__resp_plaOutput_26 ^ req_opcode[3]};
  wire [3:0]  view__resp_hi_hi_lo = {view__resp_hi_hi_lo_hi, view__resp_hi_hi_lo_lo};
  wire [1:0]  view__resp_hi_hi_hi_lo = {view__resp_plaOutput_29 ^ req_opcode[3], view__resp_plaOutput_28 ^ req_opcode[3]};
  wire [1:0]  view__resp_hi_hi_hi_hi = {view__resp_plaOutput_31 ^ req_opcode[3], view__resp_plaOutput_30 ^ req_opcode[3]};
  wire [3:0]  view__resp_hi_hi_hi = {view__resp_hi_hi_hi_hi, view__resp_hi_hi_hi_lo};
  wire [7:0]  view__resp_hi_hi = {view__resp_hi_hi_hi, view__resp_hi_hi_lo};
  wire [15:0] view__resp_hi = {view__resp_hi_hi, view__resp_hi_lo};
  assign resp = {view__resp_hi, view__resp_lo};
endmodule

