
// Include register initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for register randomization.

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_
module MaskUnit(
  input         clock,
                reset,
                instReq_valid,
  input  [2:0]  instReq_bits_instructionIndex,
  input         instReq_bits_decodeResult_specialSlot,
  input  [4:0]  instReq_bits_decodeResult_topUop,
  input         instReq_bits_decodeResult_popCount,
                instReq_bits_decodeResult_ffo,
                instReq_bits_decodeResult_average,
                instReq_bits_decodeResult_reverse,
                instReq_bits_decodeResult_dontNeedExecuteInLane,
                instReq_bits_decodeResult_scheduler,
                instReq_bits_decodeResult_sReadVD,
                instReq_bits_decodeResult_vtype,
                instReq_bits_decodeResult_sWrite,
                instReq_bits_decodeResult_crossRead,
                instReq_bits_decodeResult_crossWrite,
                instReq_bits_decodeResult_maskUnit,
                instReq_bits_decodeResult_special,
                instReq_bits_decodeResult_saturate,
                instReq_bits_decodeResult_vwmacc,
                instReq_bits_decodeResult_readOnly,
                instReq_bits_decodeResult_maskSource,
                instReq_bits_decodeResult_maskDestination,
                instReq_bits_decodeResult_maskLogic,
  input  [3:0]  instReq_bits_decodeResult_uop,
  input         instReq_bits_decodeResult_iota,
                instReq_bits_decodeResult_mv,
                instReq_bits_decodeResult_extend,
                instReq_bits_decodeResult_unOrderWrite,
                instReq_bits_decodeResult_compress,
                instReq_bits_decodeResult_gather16,
                instReq_bits_decodeResult_gather,
                instReq_bits_decodeResult_slid,
                instReq_bits_decodeResult_targetRd,
                instReq_bits_decodeResult_widenReduce,
                instReq_bits_decodeResult_red,
                instReq_bits_decodeResult_nr,
                instReq_bits_decodeResult_itype,
                instReq_bits_decodeResult_unsigned1,
                instReq_bits_decodeResult_unsigned0,
                instReq_bits_decodeResult_other,
                instReq_bits_decodeResult_multiCycle,
                instReq_bits_decodeResult_divider,
                instReq_bits_decodeResult_multiplier,
                instReq_bits_decodeResult_shift,
                instReq_bits_decodeResult_adder,
                instReq_bits_decodeResult_logic,
  input  [31:0] instReq_bits_readFromScala,
  input  [1:0]  instReq_bits_sew,
  input  [2:0]  instReq_bits_vlmul,
  input         instReq_bits_maskType,
  input  [2:0]  instReq_bits_vxrm,
  input  [4:0]  instReq_bits_vs2,
                instReq_bits_vs1,
                instReq_bits_vd,
  input  [13:0] instReq_bits_vl,
  input         exeReq_0_valid,
  input  [31:0] exeReq_0_bits_source1,
                exeReq_0_bits_source2,
  input  [2:0]  exeReq_0_bits_index,
  input         exeReq_0_bits_ffo,
                exeReq_1_valid,
  input  [31:0] exeReq_1_bits_source1,
                exeReq_1_bits_source2,
  input  [2:0]  exeReq_1_bits_index,
  input         exeReq_1_bits_ffo,
                exeReq_2_valid,
  input  [31:0] exeReq_2_bits_source1,
                exeReq_2_bits_source2,
  input  [2:0]  exeReq_2_bits_index,
  input         exeReq_2_bits_ffo,
                exeReq_3_valid,
  input  [31:0] exeReq_3_bits_source1,
                exeReq_3_bits_source2,
  input  [2:0]  exeReq_3_bits_index,
  input         exeReq_3_bits_ffo,
                exeResp_0_ready,
  output        exeResp_0_valid,
  output [4:0]  exeResp_0_bits_vd,
  output [5:0]  exeResp_0_bits_offset,
  output [3:0]  exeResp_0_bits_mask,
  output [31:0] exeResp_0_bits_data,
  output [2:0]  exeResp_0_bits_instructionIndex,
  input         exeResp_1_ready,
  output        exeResp_1_valid,
  output [4:0]  exeResp_1_bits_vd,
  output [5:0]  exeResp_1_bits_offset,
  output [3:0]  exeResp_1_bits_mask,
  output [31:0] exeResp_1_bits_data,
  output [2:0]  exeResp_1_bits_instructionIndex,
  input         exeResp_2_ready,
  output        exeResp_2_valid,
  output [4:0]  exeResp_2_bits_vd,
  output [5:0]  exeResp_2_bits_offset,
  output [3:0]  exeResp_2_bits_mask,
  output [31:0] exeResp_2_bits_data,
  output [2:0]  exeResp_2_bits_instructionIndex,
  input         exeResp_3_ready,
  output        exeResp_3_valid,
  output [4:0]  exeResp_3_bits_vd,
  output [5:0]  exeResp_3_bits_offset,
  output [3:0]  exeResp_3_bits_mask,
  output [31:0] exeResp_3_bits_data,
  output [2:0]  exeResp_3_bits_instructionIndex,
  input         writeRelease_0,
                writeRelease_1,
                writeRelease_2,
                writeRelease_3,
  output        tokenIO_0_maskRequestRelease,
                tokenIO_1_maskRequestRelease,
                tokenIO_2_maskRequestRelease,
                tokenIO_3_maskRequestRelease,
  input         readChannel_0_ready,
  output        readChannel_0_valid,
  output [4:0]  readChannel_0_bits_vs,
  output [5:0]  readChannel_0_bits_offset,
  output [2:0]  readChannel_0_bits_instructionIndex,
  input         readChannel_1_ready,
  output        readChannel_1_valid,
  output [4:0]  readChannel_1_bits_vs,
  output [5:0]  readChannel_1_bits_offset,
  output [2:0]  readChannel_1_bits_instructionIndex,
  input         readChannel_2_ready,
  output        readChannel_2_valid,
  output [4:0]  readChannel_2_bits_vs,
  output [5:0]  readChannel_2_bits_offset,
  output [2:0]  readChannel_2_bits_instructionIndex,
  input         readChannel_3_ready,
  output        readChannel_3_valid,
  output [4:0]  readChannel_3_bits_vs,
  output [5:0]  readChannel_3_bits_offset,
  output [2:0]  readChannel_3_bits_instructionIndex,
  input         readResult_0_valid,
  input  [31:0] readResult_0_bits,
  input         readResult_1_valid,
  input  [31:0] readResult_1_bits,
  input         readResult_2_valid,
  input  [31:0] readResult_2_bits,
  input         readResult_3_valid,
  input  [31:0] readResult_3_bits,
  output [7:0]  lastReport,
  output [31:0] laneMaskInput_0,
                laneMaskInput_1,
                laneMaskInput_2,
                laneMaskInput_3,
  input  [7:0]  laneMaskSelect_0,
                laneMaskSelect_1,
                laneMaskSelect_2,
                laneMaskSelect_3,
  input  [1:0]  laneMaskSewSelect_0,
                laneMaskSewSelect_1,
                laneMaskSewSelect_2,
                laneMaskSewSelect_3,
  input         v0UpdateVec_0_valid,
  input  [31:0] v0UpdateVec_0_bits_data,
  input  [5:0]  v0UpdateVec_0_bits_offset,
  input  [3:0]  v0UpdateVec_0_bits_mask,
  input         v0UpdateVec_1_valid,
  input  [31:0] v0UpdateVec_1_bits_data,
  input  [5:0]  v0UpdateVec_1_bits_offset,
  input  [3:0]  v0UpdateVec_1_bits_mask,
  input         v0UpdateVec_2_valid,
  input  [31:0] v0UpdateVec_2_bits_data,
  input  [5:0]  v0UpdateVec_2_bits_offset,
  input  [3:0]  v0UpdateVec_2_bits_mask,
  input         v0UpdateVec_3_valid,
  input  [31:0] v0UpdateVec_3_bits_data,
  input  [5:0]  v0UpdateVec_3_bits_offset,
  input  [3:0]  v0UpdateVec_3_bits_mask,
  output [31:0] writeRDData,
  input         gatherData_ready,
  output        gatherData_valid,
  output [31:0] gatherData_bits,
  input         gatherRead
);

  wire               readCrossBar_input_3_valid;
  wire               readCrossBar_input_2_valid;
  wire               readCrossBar_input_1_valid;
  wire               readCrossBar_input_0_valid;
  wire               _writeQueue_fifo_3_empty;
  wire               _writeQueue_fifo_3_full;
  wire               _writeQueue_fifo_3_error;
  wire [54:0]        _writeQueue_fifo_3_data_out;
  wire               _writeQueue_fifo_2_empty;
  wire               _writeQueue_fifo_2_full;
  wire               _writeQueue_fifo_2_error;
  wire [54:0]        _writeQueue_fifo_2_data_out;
  wire               _writeQueue_fifo_1_empty;
  wire               _writeQueue_fifo_1_full;
  wire               _writeQueue_fifo_1_error;
  wire [54:0]        _writeQueue_fifo_1_data_out;
  wire               _writeQueue_fifo_empty;
  wire               _writeQueue_fifo_full;
  wire               _writeQueue_fifo_error;
  wire [54:0]        _writeQueue_fifo_data_out;
  wire [127:0]       _extendUnit_out;
  wire               _reduceUnit_in_ready;
  wire               _reduceUnit_out_valid;
  wire [31:0]        _reduceUnit_out_bits_data;
  wire [3:0]         _reduceUnit_out_bits_mask;
  wire               _compressUnit_out_compressValid;
  wire [31:0]        _compressUnit_writeData;
  wire               _compressUnit_stageValid;
  wire               _readData_readDataQueue_fifo_3_empty;
  wire               _readData_readDataQueue_fifo_3_full;
  wire               _readData_readDataQueue_fifo_3_error;
  wire [31:0]        _readData_readDataQueue_fifo_3_data_out;
  wire               _readData_readDataQueue_fifo_2_empty;
  wire               _readData_readDataQueue_fifo_2_full;
  wire               _readData_readDataQueue_fifo_2_error;
  wire [31:0]        _readData_readDataQueue_fifo_2_data_out;
  wire               _readData_readDataQueue_fifo_1_empty;
  wire               _readData_readDataQueue_fifo_1_full;
  wire               _readData_readDataQueue_fifo_1_error;
  wire [31:0]        _readData_readDataQueue_fifo_1_data_out;
  wire               _readData_readDataQueue_fifo_empty;
  wire               _readData_readDataQueue_fifo_full;
  wire               _readData_readDataQueue_fifo_error;
  wire [31:0]        _readData_readDataQueue_fifo_data_out;
  wire               _readMessageQueue_fifo_3_empty;
  wire               _readMessageQueue_fifo_3_full;
  wire               _readMessageQueue_fifo_3_error;
  wire [5:0]         _readMessageQueue_fifo_3_data_out;
  wire               _readMessageQueue_fifo_2_empty;
  wire               _readMessageQueue_fifo_2_full;
  wire               _readMessageQueue_fifo_2_error;
  wire [5:0]         _readMessageQueue_fifo_2_data_out;
  wire               _readMessageQueue_fifo_1_empty;
  wire               _readMessageQueue_fifo_1_full;
  wire               _readMessageQueue_fifo_1_error;
  wire [5:0]         _readMessageQueue_fifo_1_data_out;
  wire               _readMessageQueue_fifo_empty;
  wire               _readMessageQueue_fifo_full;
  wire               _readMessageQueue_fifo_error;
  wire [5:0]         _readMessageQueue_fifo_data_out;
  wire               _reorderQueueVec_fifo_3_empty;
  wire               _reorderQueueVec_fifo_3_full;
  wire               _reorderQueueVec_fifo_3_error;
  wire [35:0]        _reorderQueueVec_fifo_3_data_out;
  wire               _reorderQueueVec_fifo_2_empty;
  wire               _reorderQueueVec_fifo_2_full;
  wire               _reorderQueueVec_fifo_2_error;
  wire [35:0]        _reorderQueueVec_fifo_2_data_out;
  wire               _reorderQueueVec_fifo_1_empty;
  wire               _reorderQueueVec_fifo_1_full;
  wire               _reorderQueueVec_fifo_1_error;
  wire [35:0]        _reorderQueueVec_fifo_1_data_out;
  wire               _reorderQueueVec_fifo_empty;
  wire               _reorderQueueVec_fifo_full;
  wire               _reorderQueueVec_fifo_error;
  wire [35:0]        _reorderQueueVec_fifo_data_out;
  wire               _compressUnitResultQueue_fifo_empty;
  wire               _compressUnitResultQueue_fifo_full;
  wire               _compressUnitResultQueue_fifo_error;
  wire [158:0]       _compressUnitResultQueue_fifo_data_out;
  wire               _readWaitQueue_fifo_empty;
  wire               _readWaitQueue_fifo_full;
  wire               _readWaitQueue_fifo_error;
  wire [24:0]        _readWaitQueue_fifo_data_out;
  wire               _readCrossBar_input_0_ready;
  wire               _readCrossBar_input_1_ready;
  wire               _readCrossBar_input_2_ready;
  wire               _readCrossBar_input_3_ready;
  wire               _readCrossBar_output_0_valid;
  wire [4:0]         _readCrossBar_output_0_bits_vs;
  wire [5:0]         _readCrossBar_output_0_bits_offset;
  wire [1:0]         _readCrossBar_output_0_bits_writeIndex;
  wire               _readCrossBar_output_1_valid;
  wire [4:0]         _readCrossBar_output_1_bits_vs;
  wire [5:0]         _readCrossBar_output_1_bits_offset;
  wire [1:0]         _readCrossBar_output_1_bits_writeIndex;
  wire               _readCrossBar_output_2_valid;
  wire [4:0]         _readCrossBar_output_2_bits_vs;
  wire [5:0]         _readCrossBar_output_2_bits_offset;
  wire [1:0]         _readCrossBar_output_2_bits_writeIndex;
  wire               _readCrossBar_output_3_valid;
  wire [4:0]         _readCrossBar_output_3_bits_vs;
  wire [5:0]         _readCrossBar_output_3_bits_offset;
  wire [1:0]         _readCrossBar_output_3_bits_writeIndex;
  wire               _accessCountQueue_fifo_empty;
  wire               _accessCountQueue_fifo_full;
  wire               _accessCountQueue_fifo_error;
  wire [11:0]        _accessCountQueue_fifo_data_out;
  wire               _slideAddressGen_indexDeq_valid;
  wire [3:0]         _slideAddressGen_indexDeq_bits_needRead;
  wire [3:0]         _slideAddressGen_indexDeq_bits_elementValid;
  wire [3:0]         _slideAddressGen_indexDeq_bits_replaceVs1;
  wire [23:0]        _slideAddressGen_indexDeq_bits_readOffset;
  wire [1:0]         _slideAddressGen_indexDeq_bits_accessLane_0;
  wire [1:0]         _slideAddressGen_indexDeq_bits_accessLane_1;
  wire [1:0]         _slideAddressGen_indexDeq_bits_accessLane_2;
  wire [1:0]         _slideAddressGen_indexDeq_bits_accessLane_3;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_0;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_1;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_2;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_3;
  wire [11:0]        _slideAddressGen_indexDeq_bits_executeGroup;
  wire [7:0]         _slideAddressGen_indexDeq_bits_readDataOffset;
  wire               _slideAddressGen_indexDeq_bits_last;
  wire [11:0]        _slideAddressGen_slideGroupOut;
  wire               _exeRequestQueue_queue_fifo_3_empty;
  wire               _exeRequestQueue_queue_fifo_3_full;
  wire               _exeRequestQueue_queue_fifo_3_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_3_data_out;
  wire               _exeRequestQueue_queue_fifo_2_empty;
  wire               _exeRequestQueue_queue_fifo_2_full;
  wire               _exeRequestQueue_queue_fifo_2_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_2_data_out;
  wire               _exeRequestQueue_queue_fifo_1_empty;
  wire               _exeRequestQueue_queue_fifo_1_full;
  wire               _exeRequestQueue_queue_fifo_1_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_1_data_out;
  wire               _exeRequestQueue_queue_fifo_empty;
  wire               _exeRequestQueue_queue_fifo_full;
  wire               _exeRequestQueue_queue_fifo_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_data_out;
  wire               _maskedWrite_in_0_ready;
  wire               _maskedWrite_in_1_ready;
  wire               _maskedWrite_in_2_ready;
  wire               _maskedWrite_in_3_ready;
  wire               _maskedWrite_out_0_valid;
  wire               _maskedWrite_out_0_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_0_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_0_bits_writeData_mask;
  wire [9:0]         _maskedWrite_out_0_bits_writeData_groupCounter;
  wire               _maskedWrite_out_1_valid;
  wire               _maskedWrite_out_1_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_1_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_1_bits_writeData_mask;
  wire [9:0]         _maskedWrite_out_1_bits_writeData_groupCounter;
  wire               _maskedWrite_out_2_valid;
  wire               _maskedWrite_out_2_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_2_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_2_bits_writeData_mask;
  wire [9:0]         _maskedWrite_out_2_bits_writeData_groupCounter;
  wire               _maskedWrite_out_3_valid;
  wire               _maskedWrite_out_3_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_3_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_3_bits_writeData_mask;
  wire [9:0]         _maskedWrite_out_3_bits_writeData_groupCounter;
  wire               _maskedWrite_readChannel_0_valid;
  wire [4:0]         _maskedWrite_readChannel_0_bits_vs;
  wire [5:0]         _maskedWrite_readChannel_0_bits_offset;
  wire               _maskedWrite_readChannel_1_valid;
  wire [4:0]         _maskedWrite_readChannel_1_bits_vs;
  wire [5:0]         _maskedWrite_readChannel_1_bits_offset;
  wire               _maskedWrite_readChannel_2_valid;
  wire [4:0]         _maskedWrite_readChannel_2_bits_vs;
  wire [5:0]         _maskedWrite_readChannel_2_bits_offset;
  wire               _maskedWrite_readChannel_3_valid;
  wire [4:0]         _maskedWrite_readChannel_3_bits_vs;
  wire [5:0]         _maskedWrite_readChannel_3_bits_offset;
  wire               _maskedWrite_stageClear;
  wire               writeQueue_3_almostFull;
  wire               writeQueue_3_almostEmpty;
  wire               writeQueue_2_almostFull;
  wire               writeQueue_2_almostEmpty;
  wire               writeQueue_1_almostFull;
  wire               writeQueue_1_almostEmpty;
  wire               writeQueue_0_almostFull;
  wire               writeQueue_0_almostEmpty;
  wire               readData_readDataQueue_3_almostFull;
  wire               readData_readDataQueue_3_almostEmpty;
  wire               readData_readDataQueue_2_almostFull;
  wire               readData_readDataQueue_2_almostEmpty;
  wire               readData_readDataQueue_1_almostFull;
  wire               readData_readDataQueue_1_almostEmpty;
  wire               readData_readDataQueue_almostFull;
  wire               readData_readDataQueue_almostEmpty;
  wire               readMessageQueue_3_almostFull;
  wire               readMessageQueue_3_almostEmpty;
  wire               readMessageQueue_2_almostFull;
  wire               readMessageQueue_2_almostEmpty;
  wire               readMessageQueue_1_almostFull;
  wire               readMessageQueue_1_almostEmpty;
  wire               readMessageQueue_almostFull;
  wire               readMessageQueue_almostEmpty;
  wire               reorderQueueVec_3_almostFull;
  wire               reorderQueueVec_3_almostEmpty;
  wire               reorderQueueVec_2_almostFull;
  wire               reorderQueueVec_2_almostEmpty;
  wire               reorderQueueVec_1_almostFull;
  wire               reorderQueueVec_1_almostEmpty;
  wire               reorderQueueVec_0_almostFull;
  wire               reorderQueueVec_0_almostEmpty;
  wire               compressUnitResultQueue_almostFull;
  wire               compressUnitResultQueue_almostEmpty;
  wire               readWaitQueue_almostFull;
  wire               readWaitQueue_almostEmpty;
  wire               accessCountQueue_almostFull;
  wire               accessCountQueue_almostEmpty;
  wire               exeRequestQueue_3_almostFull;
  wire               exeRequestQueue_3_almostEmpty;
  wire               exeRequestQueue_2_almostFull;
  wire               exeRequestQueue_2_almostEmpty;
  wire               exeRequestQueue_1_almostFull;
  wire               exeRequestQueue_1_almostEmpty;
  wire               exeRequestQueue_0_almostFull;
  wire               exeRequestQueue_0_almostEmpty;
  wire [31:0]        reorderQueueVec_3_deq_bits_data;
  wire [31:0]        reorderQueueVec_2_deq_bits_data;
  wire [31:0]        reorderQueueVec_1_deq_bits_data;
  wire [31:0]        reorderQueueVec_0_deq_bits_data;
  wire [2:0]         accessCountEnq_3;
  wire [2:0]         accessCountEnq_2;
  wire [2:0]         accessCountEnq_1;
  wire [2:0]         accessCountEnq_0;
  wire               exeResp_0_ready_0 = exeResp_0_ready;
  wire               exeResp_1_ready_0 = exeResp_1_ready;
  wire               exeResp_2_ready_0 = exeResp_2_ready;
  wire               exeResp_3_ready_0 = exeResp_3_ready;
  wire               readChannel_0_ready_0 = readChannel_0_ready;
  wire               readChannel_1_ready_0 = readChannel_1_ready;
  wire               readChannel_2_ready_0 = readChannel_2_ready;
  wire               readChannel_3_ready_0 = readChannel_3_ready;
  wire               gatherData_ready_0 = gatherData_ready;
  wire               exeRequestQueue_0_enq_valid = exeReq_0_valid;
  wire [31:0]        exeRequestQueue_0_enq_bits_source1 = exeReq_0_bits_source1;
  wire [31:0]        exeRequestQueue_0_enq_bits_source2 = exeReq_0_bits_source2;
  wire [2:0]         exeRequestQueue_0_enq_bits_index = exeReq_0_bits_index;
  wire               exeRequestQueue_0_enq_bits_ffo = exeReq_0_bits_ffo;
  wire               exeRequestQueue_1_enq_valid = exeReq_1_valid;
  wire [31:0]        exeRequestQueue_1_enq_bits_source1 = exeReq_1_bits_source1;
  wire [31:0]        exeRequestQueue_1_enq_bits_source2 = exeReq_1_bits_source2;
  wire [2:0]         exeRequestQueue_1_enq_bits_index = exeReq_1_bits_index;
  wire               exeRequestQueue_1_enq_bits_ffo = exeReq_1_bits_ffo;
  wire               exeRequestQueue_2_enq_valid = exeReq_2_valid;
  wire [31:0]        exeRequestQueue_2_enq_bits_source1 = exeReq_2_bits_source1;
  wire [31:0]        exeRequestQueue_2_enq_bits_source2 = exeReq_2_bits_source2;
  wire [2:0]         exeRequestQueue_2_enq_bits_index = exeReq_2_bits_index;
  wire               exeRequestQueue_2_enq_bits_ffo = exeReq_2_bits_ffo;
  wire               exeRequestQueue_3_enq_valid = exeReq_3_valid;
  wire [31:0]        exeRequestQueue_3_enq_bits_source1 = exeReq_3_bits_source1;
  wire [31:0]        exeRequestQueue_3_enq_bits_source2 = exeReq_3_bits_source2;
  wire [2:0]         exeRequestQueue_3_enq_bits_index = exeReq_3_bits_index;
  wire               exeRequestQueue_3_enq_bits_ffo = exeReq_3_bits_ffo;
  wire               reorderQueueVec_0_enq_valid = readResult_0_valid;
  wire               reorderQueueVec_1_enq_valid = readResult_1_valid;
  wire               reorderQueueVec_2_enq_valid = readResult_2_valid;
  wire               reorderQueueVec_3_enq_valid = readResult_3_valid;
  wire               readMessageQueue_deq_ready = readResult_0_valid;
  wire               readMessageQueue_1_deq_ready = readResult_1_valid;
  wire               readMessageQueue_2_deq_ready = readResult_2_valid;
  wire               readMessageQueue_3_deq_ready = readResult_3_valid;
  wire [7:0]         checkVec_checkResult_lo_14 = 8'hFF;
  wire [7:0]         checkVec_checkResult_hi_14 = 8'hFF;
  wire [15:0]        checkVec_2_0 = 16'hFFFF;
  wire [7:0]         checkVec_2_1 = 8'h0;
  wire [1:0]         readVS1Req_requestIndex = 2'h0;
  wire [1:0]         checkVec_checkResultVec_0_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_1_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_2_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_3_1_2 = 2'h0;
  wire [1:0]         selectExecuteReq_0_bits_requestIndex = 2'h0;
  wire [1:0]         selectExecuteReq_1_bits_requestIndex = 2'h1;
  wire [1:0]         selectExecuteReq_3_bits_requestIndex = 2'h3;
  wire [3:0]         checkVec_checkResult_lo_15 = 4'h0;
  wire [3:0]         checkVec_checkResult_hi_15 = 4'h0;
  wire [1:0]         readChannel_0_bits_readSource = 2'h2;
  wire [1:0]         readChannel_1_bits_readSource = 2'h2;
  wire [1:0]         readChannel_2_bits_readSource = 2'h2;
  wire [1:0]         readChannel_3_bits_readSource = 2'h2;
  wire [1:0]         selectExecuteReq_2_bits_requestIndex = 2'h2;
  wire               exeResp_0_bits_last = 1'h0;
  wire               exeResp_1_bits_last = 1'h0;
  wire               exeResp_2_bits_last = 1'h0;
  wire               exeResp_3_bits_last = 1'h0;
  wire               writeRequest_0_ffoByOther = 1'h0;
  wire               writeRequest_1_ffoByOther = 1'h0;
  wire               writeRequest_2_ffoByOther = 1'h0;
  wire               writeRequest_3_ffoByOther = 1'h0;
  wire               writeQueue_0_deq_ready = exeResp_0_ready_0;
  wire               writeQueue_0_deq_valid;
  wire [3:0]         writeQueue_0_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_0_deq_bits_writeData_data;
  wire               writeQueue_1_deq_ready = exeResp_1_ready_0;
  wire               writeQueue_1_deq_valid;
  wire [3:0]         writeQueue_1_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_1_deq_bits_writeData_data;
  wire               writeQueue_2_deq_ready = exeResp_2_ready_0;
  wire               writeQueue_2_deq_valid;
  wire [3:0]         writeQueue_2_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_2_deq_bits_writeData_data;
  wire               writeQueue_3_deq_ready = exeResp_3_ready_0;
  wire               writeQueue_3_deq_valid;
  wire [3:0]         writeQueue_3_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_3_deq_bits_writeData_data;
  wire               gatherResponse;
  reg  [31:0]        v0_0;
  reg  [31:0]        v0_1;
  reg  [31:0]        v0_2;
  reg  [31:0]        v0_3;
  reg  [31:0]        v0_4;
  reg  [31:0]        v0_5;
  reg  [31:0]        v0_6;
  reg  [31:0]        v0_7;
  reg  [31:0]        v0_8;
  reg  [31:0]        v0_9;
  reg  [31:0]        v0_10;
  reg  [31:0]        v0_11;
  reg  [31:0]        v0_12;
  reg  [31:0]        v0_13;
  reg  [31:0]        v0_14;
  reg  [31:0]        v0_15;
  reg  [31:0]        v0_16;
  reg  [31:0]        v0_17;
  reg  [31:0]        v0_18;
  reg  [31:0]        v0_19;
  reg  [31:0]        v0_20;
  reg  [31:0]        v0_21;
  reg  [31:0]        v0_22;
  reg  [31:0]        v0_23;
  reg  [31:0]        v0_24;
  reg  [31:0]        v0_25;
  reg  [31:0]        v0_26;
  reg  [31:0]        v0_27;
  reg  [31:0]        v0_28;
  reg  [31:0]        v0_29;
  reg  [31:0]        v0_30;
  reg  [31:0]        v0_31;
  reg  [31:0]        v0_32;
  reg  [31:0]        v0_33;
  reg  [31:0]        v0_34;
  reg  [31:0]        v0_35;
  reg  [31:0]        v0_36;
  reg  [31:0]        v0_37;
  reg  [31:0]        v0_38;
  reg  [31:0]        v0_39;
  reg  [31:0]        v0_40;
  reg  [31:0]        v0_41;
  reg  [31:0]        v0_42;
  reg  [31:0]        v0_43;
  reg  [31:0]        v0_44;
  reg  [31:0]        v0_45;
  reg  [31:0]        v0_46;
  reg  [31:0]        v0_47;
  reg  [31:0]        v0_48;
  reg  [31:0]        v0_49;
  reg  [31:0]        v0_50;
  reg  [31:0]        v0_51;
  reg  [31:0]        v0_52;
  reg  [31:0]        v0_53;
  reg  [31:0]        v0_54;
  reg  [31:0]        v0_55;
  reg  [31:0]        v0_56;
  reg  [31:0]        v0_57;
  reg  [31:0]        v0_58;
  reg  [31:0]        v0_59;
  reg  [31:0]        v0_60;
  reg  [31:0]        v0_61;
  reg  [31:0]        v0_62;
  reg  [31:0]        v0_63;
  reg  [31:0]        v0_64;
  reg  [31:0]        v0_65;
  reg  [31:0]        v0_66;
  reg  [31:0]        v0_67;
  reg  [31:0]        v0_68;
  reg  [31:0]        v0_69;
  reg  [31:0]        v0_70;
  reg  [31:0]        v0_71;
  reg  [31:0]        v0_72;
  reg  [31:0]        v0_73;
  reg  [31:0]        v0_74;
  reg  [31:0]        v0_75;
  reg  [31:0]        v0_76;
  reg  [31:0]        v0_77;
  reg  [31:0]        v0_78;
  reg  [31:0]        v0_79;
  reg  [31:0]        v0_80;
  reg  [31:0]        v0_81;
  reg  [31:0]        v0_82;
  reg  [31:0]        v0_83;
  reg  [31:0]        v0_84;
  reg  [31:0]        v0_85;
  reg  [31:0]        v0_86;
  reg  [31:0]        v0_87;
  reg  [31:0]        v0_88;
  reg  [31:0]        v0_89;
  reg  [31:0]        v0_90;
  reg  [31:0]        v0_91;
  reg  [31:0]        v0_92;
  reg  [31:0]        v0_93;
  reg  [31:0]        v0_94;
  reg  [31:0]        v0_95;
  reg  [31:0]        v0_96;
  reg  [31:0]        v0_97;
  reg  [31:0]        v0_98;
  reg  [31:0]        v0_99;
  reg  [31:0]        v0_100;
  reg  [31:0]        v0_101;
  reg  [31:0]        v0_102;
  reg  [31:0]        v0_103;
  reg  [31:0]        v0_104;
  reg  [31:0]        v0_105;
  reg  [31:0]        v0_106;
  reg  [31:0]        v0_107;
  reg  [31:0]        v0_108;
  reg  [31:0]        v0_109;
  reg  [31:0]        v0_110;
  reg  [31:0]        v0_111;
  reg  [31:0]        v0_112;
  reg  [31:0]        v0_113;
  reg  [31:0]        v0_114;
  reg  [31:0]        v0_115;
  reg  [31:0]        v0_116;
  reg  [31:0]        v0_117;
  reg  [31:0]        v0_118;
  reg  [31:0]        v0_119;
  reg  [31:0]        v0_120;
  reg  [31:0]        v0_121;
  reg  [31:0]        v0_122;
  reg  [31:0]        v0_123;
  reg  [31:0]        v0_124;
  reg  [31:0]        v0_125;
  reg  [31:0]        v0_126;
  reg  [31:0]        v0_127;
  reg  [31:0]        v0_128;
  reg  [31:0]        v0_129;
  reg  [31:0]        v0_130;
  reg  [31:0]        v0_131;
  reg  [31:0]        v0_132;
  reg  [31:0]        v0_133;
  reg  [31:0]        v0_134;
  reg  [31:0]        v0_135;
  reg  [31:0]        v0_136;
  reg  [31:0]        v0_137;
  reg  [31:0]        v0_138;
  reg  [31:0]        v0_139;
  reg  [31:0]        v0_140;
  reg  [31:0]        v0_141;
  reg  [31:0]        v0_142;
  reg  [31:0]        v0_143;
  reg  [31:0]        v0_144;
  reg  [31:0]        v0_145;
  reg  [31:0]        v0_146;
  reg  [31:0]        v0_147;
  reg  [31:0]        v0_148;
  reg  [31:0]        v0_149;
  reg  [31:0]        v0_150;
  reg  [31:0]        v0_151;
  reg  [31:0]        v0_152;
  reg  [31:0]        v0_153;
  reg  [31:0]        v0_154;
  reg  [31:0]        v0_155;
  reg  [31:0]        v0_156;
  reg  [31:0]        v0_157;
  reg  [31:0]        v0_158;
  reg  [31:0]        v0_159;
  reg  [31:0]        v0_160;
  reg  [31:0]        v0_161;
  reg  [31:0]        v0_162;
  reg  [31:0]        v0_163;
  reg  [31:0]        v0_164;
  reg  [31:0]        v0_165;
  reg  [31:0]        v0_166;
  reg  [31:0]        v0_167;
  reg  [31:0]        v0_168;
  reg  [31:0]        v0_169;
  reg  [31:0]        v0_170;
  reg  [31:0]        v0_171;
  reg  [31:0]        v0_172;
  reg  [31:0]        v0_173;
  reg  [31:0]        v0_174;
  reg  [31:0]        v0_175;
  reg  [31:0]        v0_176;
  reg  [31:0]        v0_177;
  reg  [31:0]        v0_178;
  reg  [31:0]        v0_179;
  reg  [31:0]        v0_180;
  reg  [31:0]        v0_181;
  reg  [31:0]        v0_182;
  reg  [31:0]        v0_183;
  reg  [31:0]        v0_184;
  reg  [31:0]        v0_185;
  reg  [31:0]        v0_186;
  reg  [31:0]        v0_187;
  reg  [31:0]        v0_188;
  reg  [31:0]        v0_189;
  reg  [31:0]        v0_190;
  reg  [31:0]        v0_191;
  reg  [31:0]        v0_192;
  reg  [31:0]        v0_193;
  reg  [31:0]        v0_194;
  reg  [31:0]        v0_195;
  reg  [31:0]        v0_196;
  reg  [31:0]        v0_197;
  reg  [31:0]        v0_198;
  reg  [31:0]        v0_199;
  reg  [31:0]        v0_200;
  reg  [31:0]        v0_201;
  reg  [31:0]        v0_202;
  reg  [31:0]        v0_203;
  reg  [31:0]        v0_204;
  reg  [31:0]        v0_205;
  reg  [31:0]        v0_206;
  reg  [31:0]        v0_207;
  reg  [31:0]        v0_208;
  reg  [31:0]        v0_209;
  reg  [31:0]        v0_210;
  reg  [31:0]        v0_211;
  reg  [31:0]        v0_212;
  reg  [31:0]        v0_213;
  reg  [31:0]        v0_214;
  reg  [31:0]        v0_215;
  reg  [31:0]        v0_216;
  reg  [31:0]        v0_217;
  reg  [31:0]        v0_218;
  reg  [31:0]        v0_219;
  reg  [31:0]        v0_220;
  reg  [31:0]        v0_221;
  reg  [31:0]        v0_222;
  reg  [31:0]        v0_223;
  reg  [31:0]        v0_224;
  reg  [31:0]        v0_225;
  reg  [31:0]        v0_226;
  reg  [31:0]        v0_227;
  reg  [31:0]        v0_228;
  reg  [31:0]        v0_229;
  reg  [31:0]        v0_230;
  reg  [31:0]        v0_231;
  reg  [31:0]        v0_232;
  reg  [31:0]        v0_233;
  reg  [31:0]        v0_234;
  reg  [31:0]        v0_235;
  reg  [31:0]        v0_236;
  reg  [31:0]        v0_237;
  reg  [31:0]        v0_238;
  reg  [31:0]        v0_239;
  reg  [31:0]        v0_240;
  reg  [31:0]        v0_241;
  reg  [31:0]        v0_242;
  reg  [31:0]        v0_243;
  reg  [31:0]        v0_244;
  reg  [31:0]        v0_245;
  reg  [31:0]        v0_246;
  reg  [31:0]        v0_247;
  reg  [31:0]        v0_248;
  reg  [31:0]        v0_249;
  reg  [31:0]        v0_250;
  reg  [31:0]        v0_251;
  reg  [31:0]        v0_252;
  reg  [31:0]        v0_253;
  reg  [31:0]        v0_254;
  reg  [31:0]        v0_255;
  wire [15:0]        maskExt_lo = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt = {maskExt_hi, maskExt_lo};
  wire [15:0]        maskExt_lo_1 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_1 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_1 = {maskExt_hi_1, maskExt_lo_1};
  wire [15:0]        maskExt_lo_2 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_2 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_2 = {maskExt_hi_2, maskExt_lo_2};
  wire [15:0]        maskExt_lo_3 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_3 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_3 = {maskExt_hi_3, maskExt_lo_3};
  wire [15:0]        maskExt_lo_4 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_4 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_4 = {maskExt_hi_4, maskExt_lo_4};
  wire [15:0]        maskExt_lo_5 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_5 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_5 = {maskExt_hi_5, maskExt_lo_5};
  wire [15:0]        maskExt_lo_6 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_6 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_6 = {maskExt_hi_6, maskExt_lo_6};
  wire [15:0]        maskExt_lo_7 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_7 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_7 = {maskExt_hi_7, maskExt_lo_7};
  wire [15:0]        maskExt_lo_8 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_8 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_8 = {maskExt_hi_8, maskExt_lo_8};
  wire [15:0]        maskExt_lo_9 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_9 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_9 = {maskExt_hi_9, maskExt_lo_9};
  wire [15:0]        maskExt_lo_10 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_10 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_10 = {maskExt_hi_10, maskExt_lo_10};
  wire [15:0]        maskExt_lo_11 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_11 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_11 = {maskExt_hi_11, maskExt_lo_11};
  wire [15:0]        maskExt_lo_12 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_12 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_12 = {maskExt_hi_12, maskExt_lo_12};
  wire [15:0]        maskExt_lo_13 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_13 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_13 = {maskExt_hi_13, maskExt_lo_13};
  wire [15:0]        maskExt_lo_14 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_14 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_14 = {maskExt_hi_14, maskExt_lo_14};
  wire [15:0]        maskExt_lo_15 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_15 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_15 = {maskExt_hi_15, maskExt_lo_15};
  wire [15:0]        maskExt_lo_16 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_16 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_16 = {maskExt_hi_16, maskExt_lo_16};
  wire [15:0]        maskExt_lo_17 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_17 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_17 = {maskExt_hi_17, maskExt_lo_17};
  wire [15:0]        maskExt_lo_18 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_18 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_18 = {maskExt_hi_18, maskExt_lo_18};
  wire [15:0]        maskExt_lo_19 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_19 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_19 = {maskExt_hi_19, maskExt_lo_19};
  wire [15:0]        maskExt_lo_20 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_20 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_20 = {maskExt_hi_20, maskExt_lo_20};
  wire [15:0]        maskExt_lo_21 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_21 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_21 = {maskExt_hi_21, maskExt_lo_21};
  wire [15:0]        maskExt_lo_22 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_22 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_22 = {maskExt_hi_22, maskExt_lo_22};
  wire [15:0]        maskExt_lo_23 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_23 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_23 = {maskExt_hi_23, maskExt_lo_23};
  wire [15:0]        maskExt_lo_24 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_24 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_24 = {maskExt_hi_24, maskExt_lo_24};
  wire [15:0]        maskExt_lo_25 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_25 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_25 = {maskExt_hi_25, maskExt_lo_25};
  wire [15:0]        maskExt_lo_26 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_26 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_26 = {maskExt_hi_26, maskExt_lo_26};
  wire [15:0]        maskExt_lo_27 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_27 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_27 = {maskExt_hi_27, maskExt_lo_27};
  wire [15:0]        maskExt_lo_28 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_28 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_28 = {maskExt_hi_28, maskExt_lo_28};
  wire [15:0]        maskExt_lo_29 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_29 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_29 = {maskExt_hi_29, maskExt_lo_29};
  wire [15:0]        maskExt_lo_30 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_30 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_30 = {maskExt_hi_30, maskExt_lo_30};
  wire [15:0]        maskExt_lo_31 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_31 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_31 = {maskExt_hi_31, maskExt_lo_31};
  wire [15:0]        maskExt_lo_32 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_32 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_32 = {maskExt_hi_32, maskExt_lo_32};
  wire [15:0]        maskExt_lo_33 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_33 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_33 = {maskExt_hi_33, maskExt_lo_33};
  wire [15:0]        maskExt_lo_34 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_34 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_34 = {maskExt_hi_34, maskExt_lo_34};
  wire [15:0]        maskExt_lo_35 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_35 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_35 = {maskExt_hi_35, maskExt_lo_35};
  wire [15:0]        maskExt_lo_36 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_36 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_36 = {maskExt_hi_36, maskExt_lo_36};
  wire [15:0]        maskExt_lo_37 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_37 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_37 = {maskExt_hi_37, maskExt_lo_37};
  wire [15:0]        maskExt_lo_38 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_38 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_38 = {maskExt_hi_38, maskExt_lo_38};
  wire [15:0]        maskExt_lo_39 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_39 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_39 = {maskExt_hi_39, maskExt_lo_39};
  wire [15:0]        maskExt_lo_40 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_40 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_40 = {maskExt_hi_40, maskExt_lo_40};
  wire [15:0]        maskExt_lo_41 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_41 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_41 = {maskExt_hi_41, maskExt_lo_41};
  wire [15:0]        maskExt_lo_42 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_42 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_42 = {maskExt_hi_42, maskExt_lo_42};
  wire [15:0]        maskExt_lo_43 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_43 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_43 = {maskExt_hi_43, maskExt_lo_43};
  wire [15:0]        maskExt_lo_44 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_44 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_44 = {maskExt_hi_44, maskExt_lo_44};
  wire [15:0]        maskExt_lo_45 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_45 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_45 = {maskExt_hi_45, maskExt_lo_45};
  wire [15:0]        maskExt_lo_46 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_46 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_46 = {maskExt_hi_46, maskExt_lo_46};
  wire [15:0]        maskExt_lo_47 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_47 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_47 = {maskExt_hi_47, maskExt_lo_47};
  wire [15:0]        maskExt_lo_48 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_48 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_48 = {maskExt_hi_48, maskExt_lo_48};
  wire [15:0]        maskExt_lo_49 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_49 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_49 = {maskExt_hi_49, maskExt_lo_49};
  wire [15:0]        maskExt_lo_50 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_50 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_50 = {maskExt_hi_50, maskExt_lo_50};
  wire [15:0]        maskExt_lo_51 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_51 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_51 = {maskExt_hi_51, maskExt_lo_51};
  wire [15:0]        maskExt_lo_52 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_52 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_52 = {maskExt_hi_52, maskExt_lo_52};
  wire [15:0]        maskExt_lo_53 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_53 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_53 = {maskExt_hi_53, maskExt_lo_53};
  wire [15:0]        maskExt_lo_54 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_54 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_54 = {maskExt_hi_54, maskExt_lo_54};
  wire [15:0]        maskExt_lo_55 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_55 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_55 = {maskExt_hi_55, maskExt_lo_55};
  wire [15:0]        maskExt_lo_56 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_56 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_56 = {maskExt_hi_56, maskExt_lo_56};
  wire [15:0]        maskExt_lo_57 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_57 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_57 = {maskExt_hi_57, maskExt_lo_57};
  wire [15:0]        maskExt_lo_58 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_58 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_58 = {maskExt_hi_58, maskExt_lo_58};
  wire [15:0]        maskExt_lo_59 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_59 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_59 = {maskExt_hi_59, maskExt_lo_59};
  wire [15:0]        maskExt_lo_60 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_60 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_60 = {maskExt_hi_60, maskExt_lo_60};
  wire [15:0]        maskExt_lo_61 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_61 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_61 = {maskExt_hi_61, maskExt_lo_61};
  wire [15:0]        maskExt_lo_62 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_62 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_62 = {maskExt_hi_62, maskExt_lo_62};
  wire [15:0]        maskExt_lo_63 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_63 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_63 = {maskExt_hi_63, maskExt_lo_63};
  wire [15:0]        maskExt_lo_64 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_64 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_64 = {maskExt_hi_64, maskExt_lo_64};
  wire [15:0]        maskExt_lo_65 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_65 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_65 = {maskExt_hi_65, maskExt_lo_65};
  wire [15:0]        maskExt_lo_66 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_66 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_66 = {maskExt_hi_66, maskExt_lo_66};
  wire [15:0]        maskExt_lo_67 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_67 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_67 = {maskExt_hi_67, maskExt_lo_67};
  wire [15:0]        maskExt_lo_68 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_68 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_68 = {maskExt_hi_68, maskExt_lo_68};
  wire [15:0]        maskExt_lo_69 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_69 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_69 = {maskExt_hi_69, maskExt_lo_69};
  wire [15:0]        maskExt_lo_70 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_70 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_70 = {maskExt_hi_70, maskExt_lo_70};
  wire [15:0]        maskExt_lo_71 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_71 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_71 = {maskExt_hi_71, maskExt_lo_71};
  wire [15:0]        maskExt_lo_72 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_72 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_72 = {maskExt_hi_72, maskExt_lo_72};
  wire [15:0]        maskExt_lo_73 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_73 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_73 = {maskExt_hi_73, maskExt_lo_73};
  wire [15:0]        maskExt_lo_74 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_74 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_74 = {maskExt_hi_74, maskExt_lo_74};
  wire [15:0]        maskExt_lo_75 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_75 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_75 = {maskExt_hi_75, maskExt_lo_75};
  wire [15:0]        maskExt_lo_76 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_76 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_76 = {maskExt_hi_76, maskExt_lo_76};
  wire [15:0]        maskExt_lo_77 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_77 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_77 = {maskExt_hi_77, maskExt_lo_77};
  wire [15:0]        maskExt_lo_78 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_78 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_78 = {maskExt_hi_78, maskExt_lo_78};
  wire [15:0]        maskExt_lo_79 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_79 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_79 = {maskExt_hi_79, maskExt_lo_79};
  wire [15:0]        maskExt_lo_80 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_80 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_80 = {maskExt_hi_80, maskExt_lo_80};
  wire [15:0]        maskExt_lo_81 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_81 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_81 = {maskExt_hi_81, maskExt_lo_81};
  wire [15:0]        maskExt_lo_82 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_82 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_82 = {maskExt_hi_82, maskExt_lo_82};
  wire [15:0]        maskExt_lo_83 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_83 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_83 = {maskExt_hi_83, maskExt_lo_83};
  wire [15:0]        maskExt_lo_84 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_84 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_84 = {maskExt_hi_84, maskExt_lo_84};
  wire [15:0]        maskExt_lo_85 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_85 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_85 = {maskExt_hi_85, maskExt_lo_85};
  wire [15:0]        maskExt_lo_86 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_86 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_86 = {maskExt_hi_86, maskExt_lo_86};
  wire [15:0]        maskExt_lo_87 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_87 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_87 = {maskExt_hi_87, maskExt_lo_87};
  wire [15:0]        maskExt_lo_88 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_88 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_88 = {maskExt_hi_88, maskExt_lo_88};
  wire [15:0]        maskExt_lo_89 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_89 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_89 = {maskExt_hi_89, maskExt_lo_89};
  wire [15:0]        maskExt_lo_90 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_90 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_90 = {maskExt_hi_90, maskExt_lo_90};
  wire [15:0]        maskExt_lo_91 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_91 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_91 = {maskExt_hi_91, maskExt_lo_91};
  wire [15:0]        maskExt_lo_92 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_92 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_92 = {maskExt_hi_92, maskExt_lo_92};
  wire [15:0]        maskExt_lo_93 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_93 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_93 = {maskExt_hi_93, maskExt_lo_93};
  wire [15:0]        maskExt_lo_94 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_94 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_94 = {maskExt_hi_94, maskExt_lo_94};
  wire [15:0]        maskExt_lo_95 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_95 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_95 = {maskExt_hi_95, maskExt_lo_95};
  wire [15:0]        maskExt_lo_96 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_96 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_96 = {maskExt_hi_96, maskExt_lo_96};
  wire [15:0]        maskExt_lo_97 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_97 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_97 = {maskExt_hi_97, maskExt_lo_97};
  wire [15:0]        maskExt_lo_98 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_98 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_98 = {maskExt_hi_98, maskExt_lo_98};
  wire [15:0]        maskExt_lo_99 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_99 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_99 = {maskExt_hi_99, maskExt_lo_99};
  wire [15:0]        maskExt_lo_100 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_100 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_100 = {maskExt_hi_100, maskExt_lo_100};
  wire [15:0]        maskExt_lo_101 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_101 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_101 = {maskExt_hi_101, maskExt_lo_101};
  wire [15:0]        maskExt_lo_102 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_102 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_102 = {maskExt_hi_102, maskExt_lo_102};
  wire [15:0]        maskExt_lo_103 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_103 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_103 = {maskExt_hi_103, maskExt_lo_103};
  wire [15:0]        maskExt_lo_104 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_104 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_104 = {maskExt_hi_104, maskExt_lo_104};
  wire [15:0]        maskExt_lo_105 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_105 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_105 = {maskExt_hi_105, maskExt_lo_105};
  wire [15:0]        maskExt_lo_106 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_106 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_106 = {maskExt_hi_106, maskExt_lo_106};
  wire [15:0]        maskExt_lo_107 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_107 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_107 = {maskExt_hi_107, maskExt_lo_107};
  wire [15:0]        maskExt_lo_108 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_108 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_108 = {maskExt_hi_108, maskExt_lo_108};
  wire [15:0]        maskExt_lo_109 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_109 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_109 = {maskExt_hi_109, maskExt_lo_109};
  wire [15:0]        maskExt_lo_110 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_110 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_110 = {maskExt_hi_110, maskExt_lo_110};
  wire [15:0]        maskExt_lo_111 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_111 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_111 = {maskExt_hi_111, maskExt_lo_111};
  wire [15:0]        maskExt_lo_112 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_112 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_112 = {maskExt_hi_112, maskExt_lo_112};
  wire [15:0]        maskExt_lo_113 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_113 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_113 = {maskExt_hi_113, maskExt_lo_113};
  wire [15:0]        maskExt_lo_114 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_114 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_114 = {maskExt_hi_114, maskExt_lo_114};
  wire [15:0]        maskExt_lo_115 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_115 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_115 = {maskExt_hi_115, maskExt_lo_115};
  wire [15:0]        maskExt_lo_116 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_116 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_116 = {maskExt_hi_116, maskExt_lo_116};
  wire [15:0]        maskExt_lo_117 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_117 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_117 = {maskExt_hi_117, maskExt_lo_117};
  wire [15:0]        maskExt_lo_118 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_118 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_118 = {maskExt_hi_118, maskExt_lo_118};
  wire [15:0]        maskExt_lo_119 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_119 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_119 = {maskExt_hi_119, maskExt_lo_119};
  wire [15:0]        maskExt_lo_120 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_120 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_120 = {maskExt_hi_120, maskExt_lo_120};
  wire [15:0]        maskExt_lo_121 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_121 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_121 = {maskExt_hi_121, maskExt_lo_121};
  wire [15:0]        maskExt_lo_122 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_122 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_122 = {maskExt_hi_122, maskExt_lo_122};
  wire [15:0]        maskExt_lo_123 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_123 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_123 = {maskExt_hi_123, maskExt_lo_123};
  wire [15:0]        maskExt_lo_124 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_124 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_124 = {maskExt_hi_124, maskExt_lo_124};
  wire [15:0]        maskExt_lo_125 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_125 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_125 = {maskExt_hi_125, maskExt_lo_125};
  wire [15:0]        maskExt_lo_126 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_126 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_126 = {maskExt_hi_126, maskExt_lo_126};
  wire [15:0]        maskExt_lo_127 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_127 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_127 = {maskExt_hi_127, maskExt_lo_127};
  wire [15:0]        maskExt_lo_128 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_128 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_128 = {maskExt_hi_128, maskExt_lo_128};
  wire [15:0]        maskExt_lo_129 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_129 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_129 = {maskExt_hi_129, maskExt_lo_129};
  wire [15:0]        maskExt_lo_130 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_130 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_130 = {maskExt_hi_130, maskExt_lo_130};
  wire [15:0]        maskExt_lo_131 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_131 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_131 = {maskExt_hi_131, maskExt_lo_131};
  wire [15:0]        maskExt_lo_132 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_132 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_132 = {maskExt_hi_132, maskExt_lo_132};
  wire [15:0]        maskExt_lo_133 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_133 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_133 = {maskExt_hi_133, maskExt_lo_133};
  wire [15:0]        maskExt_lo_134 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_134 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_134 = {maskExt_hi_134, maskExt_lo_134};
  wire [15:0]        maskExt_lo_135 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_135 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_135 = {maskExt_hi_135, maskExt_lo_135};
  wire [15:0]        maskExt_lo_136 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_136 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_136 = {maskExt_hi_136, maskExt_lo_136};
  wire [15:0]        maskExt_lo_137 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_137 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_137 = {maskExt_hi_137, maskExt_lo_137};
  wire [15:0]        maskExt_lo_138 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_138 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_138 = {maskExt_hi_138, maskExt_lo_138};
  wire [15:0]        maskExt_lo_139 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_139 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_139 = {maskExt_hi_139, maskExt_lo_139};
  wire [15:0]        maskExt_lo_140 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_140 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_140 = {maskExt_hi_140, maskExt_lo_140};
  wire [15:0]        maskExt_lo_141 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_141 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_141 = {maskExt_hi_141, maskExt_lo_141};
  wire [15:0]        maskExt_lo_142 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_142 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_142 = {maskExt_hi_142, maskExt_lo_142};
  wire [15:0]        maskExt_lo_143 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_143 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_143 = {maskExt_hi_143, maskExt_lo_143};
  wire [15:0]        maskExt_lo_144 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_144 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_144 = {maskExt_hi_144, maskExt_lo_144};
  wire [15:0]        maskExt_lo_145 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_145 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_145 = {maskExt_hi_145, maskExt_lo_145};
  wire [15:0]        maskExt_lo_146 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_146 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_146 = {maskExt_hi_146, maskExt_lo_146};
  wire [15:0]        maskExt_lo_147 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_147 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_147 = {maskExt_hi_147, maskExt_lo_147};
  wire [15:0]        maskExt_lo_148 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_148 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_148 = {maskExt_hi_148, maskExt_lo_148};
  wire [15:0]        maskExt_lo_149 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_149 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_149 = {maskExt_hi_149, maskExt_lo_149};
  wire [15:0]        maskExt_lo_150 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_150 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_150 = {maskExt_hi_150, maskExt_lo_150};
  wire [15:0]        maskExt_lo_151 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_151 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_151 = {maskExt_hi_151, maskExt_lo_151};
  wire [15:0]        maskExt_lo_152 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_152 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_152 = {maskExt_hi_152, maskExt_lo_152};
  wire [15:0]        maskExt_lo_153 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_153 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_153 = {maskExt_hi_153, maskExt_lo_153};
  wire [15:0]        maskExt_lo_154 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_154 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_154 = {maskExt_hi_154, maskExt_lo_154};
  wire [15:0]        maskExt_lo_155 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_155 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_155 = {maskExt_hi_155, maskExt_lo_155};
  wire [15:0]        maskExt_lo_156 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_156 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_156 = {maskExt_hi_156, maskExt_lo_156};
  wire [15:0]        maskExt_lo_157 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_157 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_157 = {maskExt_hi_157, maskExt_lo_157};
  wire [15:0]        maskExt_lo_158 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_158 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_158 = {maskExt_hi_158, maskExt_lo_158};
  wire [15:0]        maskExt_lo_159 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_159 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_159 = {maskExt_hi_159, maskExt_lo_159};
  wire [15:0]        maskExt_lo_160 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_160 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_160 = {maskExt_hi_160, maskExt_lo_160};
  wire [15:0]        maskExt_lo_161 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_161 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_161 = {maskExt_hi_161, maskExt_lo_161};
  wire [15:0]        maskExt_lo_162 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_162 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_162 = {maskExt_hi_162, maskExt_lo_162};
  wire [15:0]        maskExt_lo_163 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_163 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_163 = {maskExt_hi_163, maskExt_lo_163};
  wire [15:0]        maskExt_lo_164 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_164 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_164 = {maskExt_hi_164, maskExt_lo_164};
  wire [15:0]        maskExt_lo_165 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_165 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_165 = {maskExt_hi_165, maskExt_lo_165};
  wire [15:0]        maskExt_lo_166 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_166 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_166 = {maskExt_hi_166, maskExt_lo_166};
  wire [15:0]        maskExt_lo_167 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_167 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_167 = {maskExt_hi_167, maskExt_lo_167};
  wire [15:0]        maskExt_lo_168 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_168 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_168 = {maskExt_hi_168, maskExt_lo_168};
  wire [15:0]        maskExt_lo_169 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_169 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_169 = {maskExt_hi_169, maskExt_lo_169};
  wire [15:0]        maskExt_lo_170 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_170 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_170 = {maskExt_hi_170, maskExt_lo_170};
  wire [15:0]        maskExt_lo_171 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_171 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_171 = {maskExt_hi_171, maskExt_lo_171};
  wire [15:0]        maskExt_lo_172 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_172 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_172 = {maskExt_hi_172, maskExt_lo_172};
  wire [15:0]        maskExt_lo_173 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_173 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_173 = {maskExt_hi_173, maskExt_lo_173};
  wire [15:0]        maskExt_lo_174 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_174 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_174 = {maskExt_hi_174, maskExt_lo_174};
  wire [15:0]        maskExt_lo_175 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_175 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_175 = {maskExt_hi_175, maskExt_lo_175};
  wire [15:0]        maskExt_lo_176 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_176 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_176 = {maskExt_hi_176, maskExt_lo_176};
  wire [15:0]        maskExt_lo_177 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_177 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_177 = {maskExt_hi_177, maskExt_lo_177};
  wire [15:0]        maskExt_lo_178 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_178 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_178 = {maskExt_hi_178, maskExt_lo_178};
  wire [15:0]        maskExt_lo_179 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_179 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_179 = {maskExt_hi_179, maskExt_lo_179};
  wire [15:0]        maskExt_lo_180 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_180 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_180 = {maskExt_hi_180, maskExt_lo_180};
  wire [15:0]        maskExt_lo_181 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_181 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_181 = {maskExt_hi_181, maskExt_lo_181};
  wire [15:0]        maskExt_lo_182 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_182 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_182 = {maskExt_hi_182, maskExt_lo_182};
  wire [15:0]        maskExt_lo_183 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_183 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_183 = {maskExt_hi_183, maskExt_lo_183};
  wire [15:0]        maskExt_lo_184 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_184 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_184 = {maskExt_hi_184, maskExt_lo_184};
  wire [15:0]        maskExt_lo_185 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_185 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_185 = {maskExt_hi_185, maskExt_lo_185};
  wire [15:0]        maskExt_lo_186 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_186 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_186 = {maskExt_hi_186, maskExt_lo_186};
  wire [15:0]        maskExt_lo_187 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_187 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_187 = {maskExt_hi_187, maskExt_lo_187};
  wire [15:0]        maskExt_lo_188 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_188 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_188 = {maskExt_hi_188, maskExt_lo_188};
  wire [15:0]        maskExt_lo_189 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_189 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_189 = {maskExt_hi_189, maskExt_lo_189};
  wire [15:0]        maskExt_lo_190 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_190 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_190 = {maskExt_hi_190, maskExt_lo_190};
  wire [15:0]        maskExt_lo_191 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_191 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_191 = {maskExt_hi_191, maskExt_lo_191};
  wire [15:0]        maskExt_lo_192 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_192 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_192 = {maskExt_hi_192, maskExt_lo_192};
  wire [15:0]        maskExt_lo_193 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_193 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_193 = {maskExt_hi_193, maskExt_lo_193};
  wire [15:0]        maskExt_lo_194 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_194 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_194 = {maskExt_hi_194, maskExt_lo_194};
  wire [15:0]        maskExt_lo_195 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_195 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_195 = {maskExt_hi_195, maskExt_lo_195};
  wire [15:0]        maskExt_lo_196 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_196 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_196 = {maskExt_hi_196, maskExt_lo_196};
  wire [15:0]        maskExt_lo_197 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_197 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_197 = {maskExt_hi_197, maskExt_lo_197};
  wire [15:0]        maskExt_lo_198 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_198 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_198 = {maskExt_hi_198, maskExt_lo_198};
  wire [15:0]        maskExt_lo_199 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_199 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_199 = {maskExt_hi_199, maskExt_lo_199};
  wire [15:0]        maskExt_lo_200 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_200 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_200 = {maskExt_hi_200, maskExt_lo_200};
  wire [15:0]        maskExt_lo_201 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_201 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_201 = {maskExt_hi_201, maskExt_lo_201};
  wire [15:0]        maskExt_lo_202 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_202 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_202 = {maskExt_hi_202, maskExt_lo_202};
  wire [15:0]        maskExt_lo_203 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_203 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_203 = {maskExt_hi_203, maskExt_lo_203};
  wire [15:0]        maskExt_lo_204 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_204 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_204 = {maskExt_hi_204, maskExt_lo_204};
  wire [15:0]        maskExt_lo_205 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_205 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_205 = {maskExt_hi_205, maskExt_lo_205};
  wire [15:0]        maskExt_lo_206 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_206 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_206 = {maskExt_hi_206, maskExt_lo_206};
  wire [15:0]        maskExt_lo_207 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_207 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_207 = {maskExt_hi_207, maskExt_lo_207};
  wire [15:0]        maskExt_lo_208 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_208 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_208 = {maskExt_hi_208, maskExt_lo_208};
  wire [15:0]        maskExt_lo_209 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_209 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_209 = {maskExt_hi_209, maskExt_lo_209};
  wire [15:0]        maskExt_lo_210 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_210 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_210 = {maskExt_hi_210, maskExt_lo_210};
  wire [15:0]        maskExt_lo_211 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_211 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_211 = {maskExt_hi_211, maskExt_lo_211};
  wire [15:0]        maskExt_lo_212 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_212 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_212 = {maskExt_hi_212, maskExt_lo_212};
  wire [15:0]        maskExt_lo_213 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_213 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_213 = {maskExt_hi_213, maskExt_lo_213};
  wire [15:0]        maskExt_lo_214 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_214 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_214 = {maskExt_hi_214, maskExt_lo_214};
  wire [15:0]        maskExt_lo_215 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_215 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_215 = {maskExt_hi_215, maskExt_lo_215};
  wire [15:0]        maskExt_lo_216 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_216 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_216 = {maskExt_hi_216, maskExt_lo_216};
  wire [15:0]        maskExt_lo_217 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_217 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_217 = {maskExt_hi_217, maskExt_lo_217};
  wire [15:0]        maskExt_lo_218 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_218 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_218 = {maskExt_hi_218, maskExt_lo_218};
  wire [15:0]        maskExt_lo_219 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_219 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_219 = {maskExt_hi_219, maskExt_lo_219};
  wire [15:0]        maskExt_lo_220 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_220 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_220 = {maskExt_hi_220, maskExt_lo_220};
  wire [15:0]        maskExt_lo_221 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_221 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_221 = {maskExt_hi_221, maskExt_lo_221};
  wire [15:0]        maskExt_lo_222 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_222 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_222 = {maskExt_hi_222, maskExt_lo_222};
  wire [15:0]        maskExt_lo_223 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_223 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_223 = {maskExt_hi_223, maskExt_lo_223};
  wire [15:0]        maskExt_lo_224 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_224 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_224 = {maskExt_hi_224, maskExt_lo_224};
  wire [15:0]        maskExt_lo_225 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_225 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_225 = {maskExt_hi_225, maskExt_lo_225};
  wire [15:0]        maskExt_lo_226 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_226 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_226 = {maskExt_hi_226, maskExt_lo_226};
  wire [15:0]        maskExt_lo_227 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_227 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_227 = {maskExt_hi_227, maskExt_lo_227};
  wire [15:0]        maskExt_lo_228 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_228 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_228 = {maskExt_hi_228, maskExt_lo_228};
  wire [15:0]        maskExt_lo_229 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_229 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_229 = {maskExt_hi_229, maskExt_lo_229};
  wire [15:0]        maskExt_lo_230 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_230 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_230 = {maskExt_hi_230, maskExt_lo_230};
  wire [15:0]        maskExt_lo_231 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_231 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_231 = {maskExt_hi_231, maskExt_lo_231};
  wire [15:0]        maskExt_lo_232 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_232 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_232 = {maskExt_hi_232, maskExt_lo_232};
  wire [15:0]        maskExt_lo_233 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_233 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_233 = {maskExt_hi_233, maskExt_lo_233};
  wire [15:0]        maskExt_lo_234 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_234 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_234 = {maskExt_hi_234, maskExt_lo_234};
  wire [15:0]        maskExt_lo_235 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_235 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_235 = {maskExt_hi_235, maskExt_lo_235};
  wire [15:0]        maskExt_lo_236 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_236 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_236 = {maskExt_hi_236, maskExt_lo_236};
  wire [15:0]        maskExt_lo_237 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_237 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_237 = {maskExt_hi_237, maskExt_lo_237};
  wire [15:0]        maskExt_lo_238 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_238 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_238 = {maskExt_hi_238, maskExt_lo_238};
  wire [15:0]        maskExt_lo_239 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_239 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_239 = {maskExt_hi_239, maskExt_lo_239};
  wire [15:0]        maskExt_lo_240 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_240 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_240 = {maskExt_hi_240, maskExt_lo_240};
  wire [15:0]        maskExt_lo_241 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_241 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_241 = {maskExt_hi_241, maskExt_lo_241};
  wire [15:0]        maskExt_lo_242 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_242 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_242 = {maskExt_hi_242, maskExt_lo_242};
  wire [15:0]        maskExt_lo_243 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_243 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_243 = {maskExt_hi_243, maskExt_lo_243};
  wire [15:0]        maskExt_lo_244 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_244 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_244 = {maskExt_hi_244, maskExt_lo_244};
  wire [15:0]        maskExt_lo_245 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_245 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_245 = {maskExt_hi_245, maskExt_lo_245};
  wire [15:0]        maskExt_lo_246 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_246 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_246 = {maskExt_hi_246, maskExt_lo_246};
  wire [15:0]        maskExt_lo_247 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_247 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_247 = {maskExt_hi_247, maskExt_lo_247};
  wire [15:0]        maskExt_lo_248 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_248 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_248 = {maskExt_hi_248, maskExt_lo_248};
  wire [15:0]        maskExt_lo_249 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_249 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_249 = {maskExt_hi_249, maskExt_lo_249};
  wire [15:0]        maskExt_lo_250 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_250 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_250 = {maskExt_hi_250, maskExt_lo_250};
  wire [15:0]        maskExt_lo_251 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_251 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_251 = {maskExt_hi_251, maskExt_lo_251};
  wire [15:0]        maskExt_lo_252 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_252 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_252 = {maskExt_hi_252, maskExt_lo_252};
  wire [15:0]        maskExt_lo_253 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_253 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_253 = {maskExt_hi_253, maskExt_lo_253};
  wire [15:0]        maskExt_lo_254 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_254 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_254 = {maskExt_hi_254, maskExt_lo_254};
  wire [15:0]        maskExt_lo_255 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_255 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_255 = {maskExt_hi_255, maskExt_lo_255};
  wire [63:0]        _GEN = {v0_1, v0_0};
  wire [63:0]        regroupV0_lo_lo_lo_lo_lo_lo_lo;
  assign regroupV0_lo_lo_lo_lo_lo_lo_lo = _GEN;
  wire [63:0]        regroupV0_lo_lo_lo_lo_lo_lo_lo_5;
  assign regroupV0_lo_lo_lo_lo_lo_lo_lo_5 = _GEN;
  wire [63:0]        regroupV0_lo_lo_lo_lo_lo_lo_lo_10;
  assign regroupV0_lo_lo_lo_lo_lo_lo_lo_10 = _GEN;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_lo_lo_lo_lo_lo;
  assign slideAddressGen_slideMaskInput_lo_lo_lo_lo_lo_lo_lo = _GEN;
  wire [63:0]        selectReadStageMask_lo_lo_lo_lo_lo_lo_lo;
  assign selectReadStageMask_lo_lo_lo_lo_lo_lo_lo = _GEN;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_lo_lo_lo;
  assign maskSplit_maskSelect_lo_lo_lo_lo_lo_lo_lo = _GEN;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_lo_lo_lo_1;
  assign maskSplit_maskSelect_lo_lo_lo_lo_lo_lo_lo_1 = _GEN;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_lo_lo_lo_2;
  assign maskSplit_maskSelect_lo_lo_lo_lo_lo_lo_lo_2 = _GEN;
  wire [63:0]        maskForDestination_lo_lo_lo_lo_lo_lo_lo;
  assign maskForDestination_lo_lo_lo_lo_lo_lo_lo = _GEN;
  wire [63:0]        _GEN_0 = {v0_3, v0_2};
  wire [63:0]        regroupV0_lo_lo_lo_lo_lo_lo_hi;
  assign regroupV0_lo_lo_lo_lo_lo_lo_hi = _GEN_0;
  wire [63:0]        regroupV0_lo_lo_lo_lo_lo_lo_hi_5;
  assign regroupV0_lo_lo_lo_lo_lo_lo_hi_5 = _GEN_0;
  wire [63:0]        regroupV0_lo_lo_lo_lo_lo_lo_hi_10;
  assign regroupV0_lo_lo_lo_lo_lo_lo_hi_10 = _GEN_0;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_lo_lo_lo_lo_hi;
  assign slideAddressGen_slideMaskInput_lo_lo_lo_lo_lo_lo_hi = _GEN_0;
  wire [63:0]        selectReadStageMask_lo_lo_lo_lo_lo_lo_hi;
  assign selectReadStageMask_lo_lo_lo_lo_lo_lo_hi = _GEN_0;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_lo_lo_hi;
  assign maskSplit_maskSelect_lo_lo_lo_lo_lo_lo_hi = _GEN_0;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_lo_lo_hi_1;
  assign maskSplit_maskSelect_lo_lo_lo_lo_lo_lo_hi_1 = _GEN_0;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_lo_lo_hi_2;
  assign maskSplit_maskSelect_lo_lo_lo_lo_lo_lo_hi_2 = _GEN_0;
  wire [63:0]        maskForDestination_lo_lo_lo_lo_lo_lo_hi;
  assign maskForDestination_lo_lo_lo_lo_lo_lo_hi = _GEN_0;
  wire [127:0]       regroupV0_lo_lo_lo_lo_lo_lo = {regroupV0_lo_lo_lo_lo_lo_lo_hi, regroupV0_lo_lo_lo_lo_lo_lo_lo};
  wire [63:0]        _GEN_1 = {v0_5, v0_4};
  wire [63:0]        regroupV0_lo_lo_lo_lo_lo_hi_lo;
  assign regroupV0_lo_lo_lo_lo_lo_hi_lo = _GEN_1;
  wire [63:0]        regroupV0_lo_lo_lo_lo_lo_hi_lo_5;
  assign regroupV0_lo_lo_lo_lo_lo_hi_lo_5 = _GEN_1;
  wire [63:0]        regroupV0_lo_lo_lo_lo_lo_hi_lo_10;
  assign regroupV0_lo_lo_lo_lo_lo_hi_lo_10 = _GEN_1;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_lo_lo_lo_hi_lo;
  assign slideAddressGen_slideMaskInput_lo_lo_lo_lo_lo_hi_lo = _GEN_1;
  wire [63:0]        selectReadStageMask_lo_lo_lo_lo_lo_hi_lo;
  assign selectReadStageMask_lo_lo_lo_lo_lo_hi_lo = _GEN_1;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_lo_hi_lo;
  assign maskSplit_maskSelect_lo_lo_lo_lo_lo_hi_lo = _GEN_1;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_lo_hi_lo_1;
  assign maskSplit_maskSelect_lo_lo_lo_lo_lo_hi_lo_1 = _GEN_1;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_lo_hi_lo_2;
  assign maskSplit_maskSelect_lo_lo_lo_lo_lo_hi_lo_2 = _GEN_1;
  wire [63:0]        maskForDestination_lo_lo_lo_lo_lo_hi_lo;
  assign maskForDestination_lo_lo_lo_lo_lo_hi_lo = _GEN_1;
  wire [63:0]        _GEN_2 = {v0_7, v0_6};
  wire [63:0]        regroupV0_lo_lo_lo_lo_lo_hi_hi;
  assign regroupV0_lo_lo_lo_lo_lo_hi_hi = _GEN_2;
  wire [63:0]        regroupV0_lo_lo_lo_lo_lo_hi_hi_5;
  assign regroupV0_lo_lo_lo_lo_lo_hi_hi_5 = _GEN_2;
  wire [63:0]        regroupV0_lo_lo_lo_lo_lo_hi_hi_10;
  assign regroupV0_lo_lo_lo_lo_lo_hi_hi_10 = _GEN_2;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_lo_lo_lo_hi_hi;
  assign slideAddressGen_slideMaskInput_lo_lo_lo_lo_lo_hi_hi = _GEN_2;
  wire [63:0]        selectReadStageMask_lo_lo_lo_lo_lo_hi_hi;
  assign selectReadStageMask_lo_lo_lo_lo_lo_hi_hi = _GEN_2;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_lo_hi_hi;
  assign maskSplit_maskSelect_lo_lo_lo_lo_lo_hi_hi = _GEN_2;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_lo_hi_hi_1;
  assign maskSplit_maskSelect_lo_lo_lo_lo_lo_hi_hi_1 = _GEN_2;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_lo_hi_hi_2;
  assign maskSplit_maskSelect_lo_lo_lo_lo_lo_hi_hi_2 = _GEN_2;
  wire [63:0]        maskForDestination_lo_lo_lo_lo_lo_hi_hi;
  assign maskForDestination_lo_lo_lo_lo_lo_hi_hi = _GEN_2;
  wire [127:0]       regroupV0_lo_lo_lo_lo_lo_hi = {regroupV0_lo_lo_lo_lo_lo_hi_hi, regroupV0_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]       regroupV0_lo_lo_lo_lo_lo = {regroupV0_lo_lo_lo_lo_lo_hi, regroupV0_lo_lo_lo_lo_lo_lo};
  wire [63:0]        _GEN_3 = {v0_9, v0_8};
  wire [63:0]        regroupV0_lo_lo_lo_lo_hi_lo_lo;
  assign regroupV0_lo_lo_lo_lo_hi_lo_lo = _GEN_3;
  wire [63:0]        regroupV0_lo_lo_lo_lo_hi_lo_lo_5;
  assign regroupV0_lo_lo_lo_lo_hi_lo_lo_5 = _GEN_3;
  wire [63:0]        regroupV0_lo_lo_lo_lo_hi_lo_lo_10;
  assign regroupV0_lo_lo_lo_lo_hi_lo_lo_10 = _GEN_3;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_lo_lo_hi_lo_lo;
  assign slideAddressGen_slideMaskInput_lo_lo_lo_lo_hi_lo_lo = _GEN_3;
  wire [63:0]        selectReadStageMask_lo_lo_lo_lo_hi_lo_lo;
  assign selectReadStageMask_lo_lo_lo_lo_hi_lo_lo = _GEN_3;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_hi_lo_lo;
  assign maskSplit_maskSelect_lo_lo_lo_lo_hi_lo_lo = _GEN_3;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_hi_lo_lo_1;
  assign maskSplit_maskSelect_lo_lo_lo_lo_hi_lo_lo_1 = _GEN_3;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_hi_lo_lo_2;
  assign maskSplit_maskSelect_lo_lo_lo_lo_hi_lo_lo_2 = _GEN_3;
  wire [63:0]        maskForDestination_lo_lo_lo_lo_hi_lo_lo;
  assign maskForDestination_lo_lo_lo_lo_hi_lo_lo = _GEN_3;
  wire [63:0]        _GEN_4 = {v0_11, v0_10};
  wire [63:0]        regroupV0_lo_lo_lo_lo_hi_lo_hi;
  assign regroupV0_lo_lo_lo_lo_hi_lo_hi = _GEN_4;
  wire [63:0]        regroupV0_lo_lo_lo_lo_hi_lo_hi_5;
  assign regroupV0_lo_lo_lo_lo_hi_lo_hi_5 = _GEN_4;
  wire [63:0]        regroupV0_lo_lo_lo_lo_hi_lo_hi_10;
  assign regroupV0_lo_lo_lo_lo_hi_lo_hi_10 = _GEN_4;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_lo_lo_hi_lo_hi;
  assign slideAddressGen_slideMaskInput_lo_lo_lo_lo_hi_lo_hi = _GEN_4;
  wire [63:0]        selectReadStageMask_lo_lo_lo_lo_hi_lo_hi;
  assign selectReadStageMask_lo_lo_lo_lo_hi_lo_hi = _GEN_4;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_hi_lo_hi;
  assign maskSplit_maskSelect_lo_lo_lo_lo_hi_lo_hi = _GEN_4;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_hi_lo_hi_1;
  assign maskSplit_maskSelect_lo_lo_lo_lo_hi_lo_hi_1 = _GEN_4;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_hi_lo_hi_2;
  assign maskSplit_maskSelect_lo_lo_lo_lo_hi_lo_hi_2 = _GEN_4;
  wire [63:0]        maskForDestination_lo_lo_lo_lo_hi_lo_hi;
  assign maskForDestination_lo_lo_lo_lo_hi_lo_hi = _GEN_4;
  wire [127:0]       regroupV0_lo_lo_lo_lo_hi_lo = {regroupV0_lo_lo_lo_lo_hi_lo_hi, regroupV0_lo_lo_lo_lo_hi_lo_lo};
  wire [63:0]        _GEN_5 = {v0_13, v0_12};
  wire [63:0]        regroupV0_lo_lo_lo_lo_hi_hi_lo;
  assign regroupV0_lo_lo_lo_lo_hi_hi_lo = _GEN_5;
  wire [63:0]        regroupV0_lo_lo_lo_lo_hi_hi_lo_5;
  assign regroupV0_lo_lo_lo_lo_hi_hi_lo_5 = _GEN_5;
  wire [63:0]        regroupV0_lo_lo_lo_lo_hi_hi_lo_10;
  assign regroupV0_lo_lo_lo_lo_hi_hi_lo_10 = _GEN_5;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_lo_lo_hi_hi_lo;
  assign slideAddressGen_slideMaskInput_lo_lo_lo_lo_hi_hi_lo = _GEN_5;
  wire [63:0]        selectReadStageMask_lo_lo_lo_lo_hi_hi_lo;
  assign selectReadStageMask_lo_lo_lo_lo_hi_hi_lo = _GEN_5;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_hi_hi_lo;
  assign maskSplit_maskSelect_lo_lo_lo_lo_hi_hi_lo = _GEN_5;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_hi_hi_lo_1;
  assign maskSplit_maskSelect_lo_lo_lo_lo_hi_hi_lo_1 = _GEN_5;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_hi_hi_lo_2;
  assign maskSplit_maskSelect_lo_lo_lo_lo_hi_hi_lo_2 = _GEN_5;
  wire [63:0]        maskForDestination_lo_lo_lo_lo_hi_hi_lo;
  assign maskForDestination_lo_lo_lo_lo_hi_hi_lo = _GEN_5;
  wire [63:0]        _GEN_6 = {v0_15, v0_14};
  wire [63:0]        regroupV0_lo_lo_lo_lo_hi_hi_hi;
  assign regroupV0_lo_lo_lo_lo_hi_hi_hi = _GEN_6;
  wire [63:0]        regroupV0_lo_lo_lo_lo_hi_hi_hi_5;
  assign regroupV0_lo_lo_lo_lo_hi_hi_hi_5 = _GEN_6;
  wire [63:0]        regroupV0_lo_lo_lo_lo_hi_hi_hi_10;
  assign regroupV0_lo_lo_lo_lo_hi_hi_hi_10 = _GEN_6;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_lo_lo_hi_hi_hi;
  assign slideAddressGen_slideMaskInput_lo_lo_lo_lo_hi_hi_hi = _GEN_6;
  wire [63:0]        selectReadStageMask_lo_lo_lo_lo_hi_hi_hi;
  assign selectReadStageMask_lo_lo_lo_lo_hi_hi_hi = _GEN_6;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_hi_hi_hi;
  assign maskSplit_maskSelect_lo_lo_lo_lo_hi_hi_hi = _GEN_6;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_hi_hi_hi_1;
  assign maskSplit_maskSelect_lo_lo_lo_lo_hi_hi_hi_1 = _GEN_6;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_hi_hi_hi_2;
  assign maskSplit_maskSelect_lo_lo_lo_lo_hi_hi_hi_2 = _GEN_6;
  wire [63:0]        maskForDestination_lo_lo_lo_lo_hi_hi_hi;
  assign maskForDestination_lo_lo_lo_lo_hi_hi_hi = _GEN_6;
  wire [127:0]       regroupV0_lo_lo_lo_lo_hi_hi = {regroupV0_lo_lo_lo_lo_hi_hi_hi, regroupV0_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]       regroupV0_lo_lo_lo_lo_hi = {regroupV0_lo_lo_lo_lo_hi_hi, regroupV0_lo_lo_lo_lo_hi_lo};
  wire [511:0]       regroupV0_lo_lo_lo_lo = {regroupV0_lo_lo_lo_lo_hi, regroupV0_lo_lo_lo_lo_lo};
  wire [63:0]        _GEN_7 = {v0_17, v0_16};
  wire [63:0]        regroupV0_lo_lo_lo_hi_lo_lo_lo;
  assign regroupV0_lo_lo_lo_hi_lo_lo_lo = _GEN_7;
  wire [63:0]        regroupV0_lo_lo_lo_hi_lo_lo_lo_5;
  assign regroupV0_lo_lo_lo_hi_lo_lo_lo_5 = _GEN_7;
  wire [63:0]        regroupV0_lo_lo_lo_hi_lo_lo_lo_10;
  assign regroupV0_lo_lo_lo_hi_lo_lo_lo_10 = _GEN_7;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_lo_hi_lo_lo_lo;
  assign slideAddressGen_slideMaskInput_lo_lo_lo_hi_lo_lo_lo = _GEN_7;
  wire [63:0]        selectReadStageMask_lo_lo_lo_hi_lo_lo_lo;
  assign selectReadStageMask_lo_lo_lo_hi_lo_lo_lo = _GEN_7;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_lo_lo_lo;
  assign maskSplit_maskSelect_lo_lo_lo_hi_lo_lo_lo = _GEN_7;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_lo_lo_lo_1;
  assign maskSplit_maskSelect_lo_lo_lo_hi_lo_lo_lo_1 = _GEN_7;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_lo_lo_lo_2;
  assign maskSplit_maskSelect_lo_lo_lo_hi_lo_lo_lo_2 = _GEN_7;
  wire [63:0]        maskForDestination_lo_lo_lo_hi_lo_lo_lo;
  assign maskForDestination_lo_lo_lo_hi_lo_lo_lo = _GEN_7;
  wire [63:0]        _GEN_8 = {v0_19, v0_18};
  wire [63:0]        regroupV0_lo_lo_lo_hi_lo_lo_hi;
  assign regroupV0_lo_lo_lo_hi_lo_lo_hi = _GEN_8;
  wire [63:0]        regroupV0_lo_lo_lo_hi_lo_lo_hi_5;
  assign regroupV0_lo_lo_lo_hi_lo_lo_hi_5 = _GEN_8;
  wire [63:0]        regroupV0_lo_lo_lo_hi_lo_lo_hi_10;
  assign regroupV0_lo_lo_lo_hi_lo_lo_hi_10 = _GEN_8;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_lo_hi_lo_lo_hi;
  assign slideAddressGen_slideMaskInput_lo_lo_lo_hi_lo_lo_hi = _GEN_8;
  wire [63:0]        selectReadStageMask_lo_lo_lo_hi_lo_lo_hi;
  assign selectReadStageMask_lo_lo_lo_hi_lo_lo_hi = _GEN_8;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_lo_lo_hi;
  assign maskSplit_maskSelect_lo_lo_lo_hi_lo_lo_hi = _GEN_8;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_lo_lo_hi_1;
  assign maskSplit_maskSelect_lo_lo_lo_hi_lo_lo_hi_1 = _GEN_8;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_lo_lo_hi_2;
  assign maskSplit_maskSelect_lo_lo_lo_hi_lo_lo_hi_2 = _GEN_8;
  wire [63:0]        maskForDestination_lo_lo_lo_hi_lo_lo_hi;
  assign maskForDestination_lo_lo_lo_hi_lo_lo_hi = _GEN_8;
  wire [127:0]       regroupV0_lo_lo_lo_hi_lo_lo = {regroupV0_lo_lo_lo_hi_lo_lo_hi, regroupV0_lo_lo_lo_hi_lo_lo_lo};
  wire [63:0]        _GEN_9 = {v0_21, v0_20};
  wire [63:0]        regroupV0_lo_lo_lo_hi_lo_hi_lo;
  assign regroupV0_lo_lo_lo_hi_lo_hi_lo = _GEN_9;
  wire [63:0]        regroupV0_lo_lo_lo_hi_lo_hi_lo_5;
  assign regroupV0_lo_lo_lo_hi_lo_hi_lo_5 = _GEN_9;
  wire [63:0]        regroupV0_lo_lo_lo_hi_lo_hi_lo_10;
  assign regroupV0_lo_lo_lo_hi_lo_hi_lo_10 = _GEN_9;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_lo_hi_lo_hi_lo;
  assign slideAddressGen_slideMaskInput_lo_lo_lo_hi_lo_hi_lo = _GEN_9;
  wire [63:0]        selectReadStageMask_lo_lo_lo_hi_lo_hi_lo;
  assign selectReadStageMask_lo_lo_lo_hi_lo_hi_lo = _GEN_9;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_lo_hi_lo;
  assign maskSplit_maskSelect_lo_lo_lo_hi_lo_hi_lo = _GEN_9;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_lo_hi_lo_1;
  assign maskSplit_maskSelect_lo_lo_lo_hi_lo_hi_lo_1 = _GEN_9;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_lo_hi_lo_2;
  assign maskSplit_maskSelect_lo_lo_lo_hi_lo_hi_lo_2 = _GEN_9;
  wire [63:0]        maskForDestination_lo_lo_lo_hi_lo_hi_lo;
  assign maskForDestination_lo_lo_lo_hi_lo_hi_lo = _GEN_9;
  wire [63:0]        _GEN_10 = {v0_23, v0_22};
  wire [63:0]        regroupV0_lo_lo_lo_hi_lo_hi_hi;
  assign regroupV0_lo_lo_lo_hi_lo_hi_hi = _GEN_10;
  wire [63:0]        regroupV0_lo_lo_lo_hi_lo_hi_hi_5;
  assign regroupV0_lo_lo_lo_hi_lo_hi_hi_5 = _GEN_10;
  wire [63:0]        regroupV0_lo_lo_lo_hi_lo_hi_hi_10;
  assign regroupV0_lo_lo_lo_hi_lo_hi_hi_10 = _GEN_10;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_lo_hi_lo_hi_hi;
  assign slideAddressGen_slideMaskInput_lo_lo_lo_hi_lo_hi_hi = _GEN_10;
  wire [63:0]        selectReadStageMask_lo_lo_lo_hi_lo_hi_hi;
  assign selectReadStageMask_lo_lo_lo_hi_lo_hi_hi = _GEN_10;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_lo_hi_hi;
  assign maskSplit_maskSelect_lo_lo_lo_hi_lo_hi_hi = _GEN_10;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_lo_hi_hi_1;
  assign maskSplit_maskSelect_lo_lo_lo_hi_lo_hi_hi_1 = _GEN_10;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_lo_hi_hi_2;
  assign maskSplit_maskSelect_lo_lo_lo_hi_lo_hi_hi_2 = _GEN_10;
  wire [63:0]        maskForDestination_lo_lo_lo_hi_lo_hi_hi;
  assign maskForDestination_lo_lo_lo_hi_lo_hi_hi = _GEN_10;
  wire [127:0]       regroupV0_lo_lo_lo_hi_lo_hi = {regroupV0_lo_lo_lo_hi_lo_hi_hi, regroupV0_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]       regroupV0_lo_lo_lo_hi_lo = {regroupV0_lo_lo_lo_hi_lo_hi, regroupV0_lo_lo_lo_hi_lo_lo};
  wire [63:0]        _GEN_11 = {v0_25, v0_24};
  wire [63:0]        regroupV0_lo_lo_lo_hi_hi_lo_lo;
  assign regroupV0_lo_lo_lo_hi_hi_lo_lo = _GEN_11;
  wire [63:0]        regroupV0_lo_lo_lo_hi_hi_lo_lo_5;
  assign regroupV0_lo_lo_lo_hi_hi_lo_lo_5 = _GEN_11;
  wire [63:0]        regroupV0_lo_lo_lo_hi_hi_lo_lo_10;
  assign regroupV0_lo_lo_lo_hi_hi_lo_lo_10 = _GEN_11;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_lo_hi_hi_lo_lo;
  assign slideAddressGen_slideMaskInput_lo_lo_lo_hi_hi_lo_lo = _GEN_11;
  wire [63:0]        selectReadStageMask_lo_lo_lo_hi_hi_lo_lo;
  assign selectReadStageMask_lo_lo_lo_hi_hi_lo_lo = _GEN_11;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_hi_lo_lo;
  assign maskSplit_maskSelect_lo_lo_lo_hi_hi_lo_lo = _GEN_11;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_hi_lo_lo_1;
  assign maskSplit_maskSelect_lo_lo_lo_hi_hi_lo_lo_1 = _GEN_11;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_hi_lo_lo_2;
  assign maskSplit_maskSelect_lo_lo_lo_hi_hi_lo_lo_2 = _GEN_11;
  wire [63:0]        maskForDestination_lo_lo_lo_hi_hi_lo_lo;
  assign maskForDestination_lo_lo_lo_hi_hi_lo_lo = _GEN_11;
  wire [63:0]        _GEN_12 = {v0_27, v0_26};
  wire [63:0]        regroupV0_lo_lo_lo_hi_hi_lo_hi;
  assign regroupV0_lo_lo_lo_hi_hi_lo_hi = _GEN_12;
  wire [63:0]        regroupV0_lo_lo_lo_hi_hi_lo_hi_5;
  assign regroupV0_lo_lo_lo_hi_hi_lo_hi_5 = _GEN_12;
  wire [63:0]        regroupV0_lo_lo_lo_hi_hi_lo_hi_10;
  assign regroupV0_lo_lo_lo_hi_hi_lo_hi_10 = _GEN_12;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_lo_hi_hi_lo_hi;
  assign slideAddressGen_slideMaskInput_lo_lo_lo_hi_hi_lo_hi = _GEN_12;
  wire [63:0]        selectReadStageMask_lo_lo_lo_hi_hi_lo_hi;
  assign selectReadStageMask_lo_lo_lo_hi_hi_lo_hi = _GEN_12;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_hi_lo_hi;
  assign maskSplit_maskSelect_lo_lo_lo_hi_hi_lo_hi = _GEN_12;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_hi_lo_hi_1;
  assign maskSplit_maskSelect_lo_lo_lo_hi_hi_lo_hi_1 = _GEN_12;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_hi_lo_hi_2;
  assign maskSplit_maskSelect_lo_lo_lo_hi_hi_lo_hi_2 = _GEN_12;
  wire [63:0]        maskForDestination_lo_lo_lo_hi_hi_lo_hi;
  assign maskForDestination_lo_lo_lo_hi_hi_lo_hi = _GEN_12;
  wire [127:0]       regroupV0_lo_lo_lo_hi_hi_lo = {regroupV0_lo_lo_lo_hi_hi_lo_hi, regroupV0_lo_lo_lo_hi_hi_lo_lo};
  wire [63:0]        _GEN_13 = {v0_29, v0_28};
  wire [63:0]        regroupV0_lo_lo_lo_hi_hi_hi_lo;
  assign regroupV0_lo_lo_lo_hi_hi_hi_lo = _GEN_13;
  wire [63:0]        regroupV0_lo_lo_lo_hi_hi_hi_lo_5;
  assign regroupV0_lo_lo_lo_hi_hi_hi_lo_5 = _GEN_13;
  wire [63:0]        regroupV0_lo_lo_lo_hi_hi_hi_lo_10;
  assign regroupV0_lo_lo_lo_hi_hi_hi_lo_10 = _GEN_13;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_lo_hi_hi_hi_lo;
  assign slideAddressGen_slideMaskInput_lo_lo_lo_hi_hi_hi_lo = _GEN_13;
  wire [63:0]        selectReadStageMask_lo_lo_lo_hi_hi_hi_lo;
  assign selectReadStageMask_lo_lo_lo_hi_hi_hi_lo = _GEN_13;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_hi_hi_lo;
  assign maskSplit_maskSelect_lo_lo_lo_hi_hi_hi_lo = _GEN_13;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_hi_hi_lo_1;
  assign maskSplit_maskSelect_lo_lo_lo_hi_hi_hi_lo_1 = _GEN_13;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_hi_hi_lo_2;
  assign maskSplit_maskSelect_lo_lo_lo_hi_hi_hi_lo_2 = _GEN_13;
  wire [63:0]        maskForDestination_lo_lo_lo_hi_hi_hi_lo;
  assign maskForDestination_lo_lo_lo_hi_hi_hi_lo = _GEN_13;
  wire [63:0]        _GEN_14 = {v0_31, v0_30};
  wire [63:0]        regroupV0_lo_lo_lo_hi_hi_hi_hi;
  assign regroupV0_lo_lo_lo_hi_hi_hi_hi = _GEN_14;
  wire [63:0]        regroupV0_lo_lo_lo_hi_hi_hi_hi_5;
  assign regroupV0_lo_lo_lo_hi_hi_hi_hi_5 = _GEN_14;
  wire [63:0]        regroupV0_lo_lo_lo_hi_hi_hi_hi_10;
  assign regroupV0_lo_lo_lo_hi_hi_hi_hi_10 = _GEN_14;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_lo_hi_hi_hi_hi;
  assign slideAddressGen_slideMaskInput_lo_lo_lo_hi_hi_hi_hi = _GEN_14;
  wire [63:0]        selectReadStageMask_lo_lo_lo_hi_hi_hi_hi;
  assign selectReadStageMask_lo_lo_lo_hi_hi_hi_hi = _GEN_14;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_hi_hi_hi;
  assign maskSplit_maskSelect_lo_lo_lo_hi_hi_hi_hi = _GEN_14;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_hi_hi_hi_1;
  assign maskSplit_maskSelect_lo_lo_lo_hi_hi_hi_hi_1 = _GEN_14;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_hi_hi_hi_2;
  assign maskSplit_maskSelect_lo_lo_lo_hi_hi_hi_hi_2 = _GEN_14;
  wire [63:0]        maskForDestination_lo_lo_lo_hi_hi_hi_hi;
  assign maskForDestination_lo_lo_lo_hi_hi_hi_hi = _GEN_14;
  wire [127:0]       regroupV0_lo_lo_lo_hi_hi_hi = {regroupV0_lo_lo_lo_hi_hi_hi_hi, regroupV0_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]       regroupV0_lo_lo_lo_hi_hi = {regroupV0_lo_lo_lo_hi_hi_hi, regroupV0_lo_lo_lo_hi_hi_lo};
  wire [511:0]       regroupV0_lo_lo_lo_hi = {regroupV0_lo_lo_lo_hi_hi, regroupV0_lo_lo_lo_hi_lo};
  wire [1023:0]      regroupV0_lo_lo_lo = {regroupV0_lo_lo_lo_hi, regroupV0_lo_lo_lo_lo};
  wire [63:0]        _GEN_15 = {v0_33, v0_32};
  wire [63:0]        regroupV0_lo_lo_hi_lo_lo_lo_lo;
  assign regroupV0_lo_lo_hi_lo_lo_lo_lo = _GEN_15;
  wire [63:0]        regroupV0_lo_lo_hi_lo_lo_lo_lo_5;
  assign regroupV0_lo_lo_hi_lo_lo_lo_lo_5 = _GEN_15;
  wire [63:0]        regroupV0_lo_lo_hi_lo_lo_lo_lo_10;
  assign regroupV0_lo_lo_hi_lo_lo_lo_lo_10 = _GEN_15;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_hi_lo_lo_lo_lo;
  assign slideAddressGen_slideMaskInput_lo_lo_hi_lo_lo_lo_lo = _GEN_15;
  wire [63:0]        selectReadStageMask_lo_lo_hi_lo_lo_lo_lo;
  assign selectReadStageMask_lo_lo_hi_lo_lo_lo_lo = _GEN_15;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_lo_lo_lo;
  assign maskSplit_maskSelect_lo_lo_hi_lo_lo_lo_lo = _GEN_15;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_lo_lo_lo_1;
  assign maskSplit_maskSelect_lo_lo_hi_lo_lo_lo_lo_1 = _GEN_15;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_lo_lo_lo_2;
  assign maskSplit_maskSelect_lo_lo_hi_lo_lo_lo_lo_2 = _GEN_15;
  wire [63:0]        maskForDestination_lo_lo_hi_lo_lo_lo_lo;
  assign maskForDestination_lo_lo_hi_lo_lo_lo_lo = _GEN_15;
  wire [63:0]        _GEN_16 = {v0_35, v0_34};
  wire [63:0]        regroupV0_lo_lo_hi_lo_lo_lo_hi;
  assign regroupV0_lo_lo_hi_lo_lo_lo_hi = _GEN_16;
  wire [63:0]        regroupV0_lo_lo_hi_lo_lo_lo_hi_5;
  assign regroupV0_lo_lo_hi_lo_lo_lo_hi_5 = _GEN_16;
  wire [63:0]        regroupV0_lo_lo_hi_lo_lo_lo_hi_10;
  assign regroupV0_lo_lo_hi_lo_lo_lo_hi_10 = _GEN_16;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_hi_lo_lo_lo_hi;
  assign slideAddressGen_slideMaskInput_lo_lo_hi_lo_lo_lo_hi = _GEN_16;
  wire [63:0]        selectReadStageMask_lo_lo_hi_lo_lo_lo_hi;
  assign selectReadStageMask_lo_lo_hi_lo_lo_lo_hi = _GEN_16;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_lo_lo_hi;
  assign maskSplit_maskSelect_lo_lo_hi_lo_lo_lo_hi = _GEN_16;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_lo_lo_hi_1;
  assign maskSplit_maskSelect_lo_lo_hi_lo_lo_lo_hi_1 = _GEN_16;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_lo_lo_hi_2;
  assign maskSplit_maskSelect_lo_lo_hi_lo_lo_lo_hi_2 = _GEN_16;
  wire [63:0]        maskForDestination_lo_lo_hi_lo_lo_lo_hi;
  assign maskForDestination_lo_lo_hi_lo_lo_lo_hi = _GEN_16;
  wire [127:0]       regroupV0_lo_lo_hi_lo_lo_lo = {regroupV0_lo_lo_hi_lo_lo_lo_hi, regroupV0_lo_lo_hi_lo_lo_lo_lo};
  wire [63:0]        _GEN_17 = {v0_37, v0_36};
  wire [63:0]        regroupV0_lo_lo_hi_lo_lo_hi_lo;
  assign regroupV0_lo_lo_hi_lo_lo_hi_lo = _GEN_17;
  wire [63:0]        regroupV0_lo_lo_hi_lo_lo_hi_lo_5;
  assign regroupV0_lo_lo_hi_lo_lo_hi_lo_5 = _GEN_17;
  wire [63:0]        regroupV0_lo_lo_hi_lo_lo_hi_lo_10;
  assign regroupV0_lo_lo_hi_lo_lo_hi_lo_10 = _GEN_17;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_hi_lo_lo_hi_lo;
  assign slideAddressGen_slideMaskInput_lo_lo_hi_lo_lo_hi_lo = _GEN_17;
  wire [63:0]        selectReadStageMask_lo_lo_hi_lo_lo_hi_lo;
  assign selectReadStageMask_lo_lo_hi_lo_lo_hi_lo = _GEN_17;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_lo_hi_lo;
  assign maskSplit_maskSelect_lo_lo_hi_lo_lo_hi_lo = _GEN_17;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_lo_hi_lo_1;
  assign maskSplit_maskSelect_lo_lo_hi_lo_lo_hi_lo_1 = _GEN_17;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_lo_hi_lo_2;
  assign maskSplit_maskSelect_lo_lo_hi_lo_lo_hi_lo_2 = _GEN_17;
  wire [63:0]        maskForDestination_lo_lo_hi_lo_lo_hi_lo;
  assign maskForDestination_lo_lo_hi_lo_lo_hi_lo = _GEN_17;
  wire [63:0]        _GEN_18 = {v0_39, v0_38};
  wire [63:0]        regroupV0_lo_lo_hi_lo_lo_hi_hi;
  assign regroupV0_lo_lo_hi_lo_lo_hi_hi = _GEN_18;
  wire [63:0]        regroupV0_lo_lo_hi_lo_lo_hi_hi_5;
  assign regroupV0_lo_lo_hi_lo_lo_hi_hi_5 = _GEN_18;
  wire [63:0]        regroupV0_lo_lo_hi_lo_lo_hi_hi_10;
  assign regroupV0_lo_lo_hi_lo_lo_hi_hi_10 = _GEN_18;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_hi_lo_lo_hi_hi;
  assign slideAddressGen_slideMaskInput_lo_lo_hi_lo_lo_hi_hi = _GEN_18;
  wire [63:0]        selectReadStageMask_lo_lo_hi_lo_lo_hi_hi;
  assign selectReadStageMask_lo_lo_hi_lo_lo_hi_hi = _GEN_18;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_lo_hi_hi;
  assign maskSplit_maskSelect_lo_lo_hi_lo_lo_hi_hi = _GEN_18;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_lo_hi_hi_1;
  assign maskSplit_maskSelect_lo_lo_hi_lo_lo_hi_hi_1 = _GEN_18;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_lo_hi_hi_2;
  assign maskSplit_maskSelect_lo_lo_hi_lo_lo_hi_hi_2 = _GEN_18;
  wire [63:0]        maskForDestination_lo_lo_hi_lo_lo_hi_hi;
  assign maskForDestination_lo_lo_hi_lo_lo_hi_hi = _GEN_18;
  wire [127:0]       regroupV0_lo_lo_hi_lo_lo_hi = {regroupV0_lo_lo_hi_lo_lo_hi_hi, regroupV0_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]       regroupV0_lo_lo_hi_lo_lo = {regroupV0_lo_lo_hi_lo_lo_hi, regroupV0_lo_lo_hi_lo_lo_lo};
  wire [63:0]        _GEN_19 = {v0_41, v0_40};
  wire [63:0]        regroupV0_lo_lo_hi_lo_hi_lo_lo;
  assign regroupV0_lo_lo_hi_lo_hi_lo_lo = _GEN_19;
  wire [63:0]        regroupV0_lo_lo_hi_lo_hi_lo_lo_5;
  assign regroupV0_lo_lo_hi_lo_hi_lo_lo_5 = _GEN_19;
  wire [63:0]        regroupV0_lo_lo_hi_lo_hi_lo_lo_10;
  assign regroupV0_lo_lo_hi_lo_hi_lo_lo_10 = _GEN_19;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_hi_lo_hi_lo_lo;
  assign slideAddressGen_slideMaskInput_lo_lo_hi_lo_hi_lo_lo = _GEN_19;
  wire [63:0]        selectReadStageMask_lo_lo_hi_lo_hi_lo_lo;
  assign selectReadStageMask_lo_lo_hi_lo_hi_lo_lo = _GEN_19;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_hi_lo_lo;
  assign maskSplit_maskSelect_lo_lo_hi_lo_hi_lo_lo = _GEN_19;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_hi_lo_lo_1;
  assign maskSplit_maskSelect_lo_lo_hi_lo_hi_lo_lo_1 = _GEN_19;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_hi_lo_lo_2;
  assign maskSplit_maskSelect_lo_lo_hi_lo_hi_lo_lo_2 = _GEN_19;
  wire [63:0]        maskForDestination_lo_lo_hi_lo_hi_lo_lo;
  assign maskForDestination_lo_lo_hi_lo_hi_lo_lo = _GEN_19;
  wire [63:0]        _GEN_20 = {v0_43, v0_42};
  wire [63:0]        regroupV0_lo_lo_hi_lo_hi_lo_hi;
  assign regroupV0_lo_lo_hi_lo_hi_lo_hi = _GEN_20;
  wire [63:0]        regroupV0_lo_lo_hi_lo_hi_lo_hi_5;
  assign regroupV0_lo_lo_hi_lo_hi_lo_hi_5 = _GEN_20;
  wire [63:0]        regroupV0_lo_lo_hi_lo_hi_lo_hi_10;
  assign regroupV0_lo_lo_hi_lo_hi_lo_hi_10 = _GEN_20;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_hi_lo_hi_lo_hi;
  assign slideAddressGen_slideMaskInput_lo_lo_hi_lo_hi_lo_hi = _GEN_20;
  wire [63:0]        selectReadStageMask_lo_lo_hi_lo_hi_lo_hi;
  assign selectReadStageMask_lo_lo_hi_lo_hi_lo_hi = _GEN_20;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_hi_lo_hi;
  assign maskSplit_maskSelect_lo_lo_hi_lo_hi_lo_hi = _GEN_20;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_hi_lo_hi_1;
  assign maskSplit_maskSelect_lo_lo_hi_lo_hi_lo_hi_1 = _GEN_20;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_hi_lo_hi_2;
  assign maskSplit_maskSelect_lo_lo_hi_lo_hi_lo_hi_2 = _GEN_20;
  wire [63:0]        maskForDestination_lo_lo_hi_lo_hi_lo_hi;
  assign maskForDestination_lo_lo_hi_lo_hi_lo_hi = _GEN_20;
  wire [127:0]       regroupV0_lo_lo_hi_lo_hi_lo = {regroupV0_lo_lo_hi_lo_hi_lo_hi, regroupV0_lo_lo_hi_lo_hi_lo_lo};
  wire [63:0]        _GEN_21 = {v0_45, v0_44};
  wire [63:0]        regroupV0_lo_lo_hi_lo_hi_hi_lo;
  assign regroupV0_lo_lo_hi_lo_hi_hi_lo = _GEN_21;
  wire [63:0]        regroupV0_lo_lo_hi_lo_hi_hi_lo_5;
  assign regroupV0_lo_lo_hi_lo_hi_hi_lo_5 = _GEN_21;
  wire [63:0]        regroupV0_lo_lo_hi_lo_hi_hi_lo_10;
  assign regroupV0_lo_lo_hi_lo_hi_hi_lo_10 = _GEN_21;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_hi_lo_hi_hi_lo;
  assign slideAddressGen_slideMaskInput_lo_lo_hi_lo_hi_hi_lo = _GEN_21;
  wire [63:0]        selectReadStageMask_lo_lo_hi_lo_hi_hi_lo;
  assign selectReadStageMask_lo_lo_hi_lo_hi_hi_lo = _GEN_21;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_hi_hi_lo;
  assign maskSplit_maskSelect_lo_lo_hi_lo_hi_hi_lo = _GEN_21;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_hi_hi_lo_1;
  assign maskSplit_maskSelect_lo_lo_hi_lo_hi_hi_lo_1 = _GEN_21;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_hi_hi_lo_2;
  assign maskSplit_maskSelect_lo_lo_hi_lo_hi_hi_lo_2 = _GEN_21;
  wire [63:0]        maskForDestination_lo_lo_hi_lo_hi_hi_lo;
  assign maskForDestination_lo_lo_hi_lo_hi_hi_lo = _GEN_21;
  wire [63:0]        _GEN_22 = {v0_47, v0_46};
  wire [63:0]        regroupV0_lo_lo_hi_lo_hi_hi_hi;
  assign regroupV0_lo_lo_hi_lo_hi_hi_hi = _GEN_22;
  wire [63:0]        regroupV0_lo_lo_hi_lo_hi_hi_hi_5;
  assign regroupV0_lo_lo_hi_lo_hi_hi_hi_5 = _GEN_22;
  wire [63:0]        regroupV0_lo_lo_hi_lo_hi_hi_hi_10;
  assign regroupV0_lo_lo_hi_lo_hi_hi_hi_10 = _GEN_22;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_hi_lo_hi_hi_hi;
  assign slideAddressGen_slideMaskInput_lo_lo_hi_lo_hi_hi_hi = _GEN_22;
  wire [63:0]        selectReadStageMask_lo_lo_hi_lo_hi_hi_hi;
  assign selectReadStageMask_lo_lo_hi_lo_hi_hi_hi = _GEN_22;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_hi_hi_hi;
  assign maskSplit_maskSelect_lo_lo_hi_lo_hi_hi_hi = _GEN_22;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_hi_hi_hi_1;
  assign maskSplit_maskSelect_lo_lo_hi_lo_hi_hi_hi_1 = _GEN_22;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_hi_hi_hi_2;
  assign maskSplit_maskSelect_lo_lo_hi_lo_hi_hi_hi_2 = _GEN_22;
  wire [63:0]        maskForDestination_lo_lo_hi_lo_hi_hi_hi;
  assign maskForDestination_lo_lo_hi_lo_hi_hi_hi = _GEN_22;
  wire [127:0]       regroupV0_lo_lo_hi_lo_hi_hi = {regroupV0_lo_lo_hi_lo_hi_hi_hi, regroupV0_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]       regroupV0_lo_lo_hi_lo_hi = {regroupV0_lo_lo_hi_lo_hi_hi, regroupV0_lo_lo_hi_lo_hi_lo};
  wire [511:0]       regroupV0_lo_lo_hi_lo = {regroupV0_lo_lo_hi_lo_hi, regroupV0_lo_lo_hi_lo_lo};
  wire [63:0]        _GEN_23 = {v0_49, v0_48};
  wire [63:0]        regroupV0_lo_lo_hi_hi_lo_lo_lo;
  assign regroupV0_lo_lo_hi_hi_lo_lo_lo = _GEN_23;
  wire [63:0]        regroupV0_lo_lo_hi_hi_lo_lo_lo_5;
  assign regroupV0_lo_lo_hi_hi_lo_lo_lo_5 = _GEN_23;
  wire [63:0]        regroupV0_lo_lo_hi_hi_lo_lo_lo_10;
  assign regroupV0_lo_lo_hi_hi_lo_lo_lo_10 = _GEN_23;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_hi_hi_lo_lo_lo;
  assign slideAddressGen_slideMaskInput_lo_lo_hi_hi_lo_lo_lo = _GEN_23;
  wire [63:0]        selectReadStageMask_lo_lo_hi_hi_lo_lo_lo;
  assign selectReadStageMask_lo_lo_hi_hi_lo_lo_lo = _GEN_23;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_lo_lo_lo;
  assign maskSplit_maskSelect_lo_lo_hi_hi_lo_lo_lo = _GEN_23;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_lo_lo_lo_1;
  assign maskSplit_maskSelect_lo_lo_hi_hi_lo_lo_lo_1 = _GEN_23;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_lo_lo_lo_2;
  assign maskSplit_maskSelect_lo_lo_hi_hi_lo_lo_lo_2 = _GEN_23;
  wire [63:0]        maskForDestination_lo_lo_hi_hi_lo_lo_lo;
  assign maskForDestination_lo_lo_hi_hi_lo_lo_lo = _GEN_23;
  wire [63:0]        _GEN_24 = {v0_51, v0_50};
  wire [63:0]        regroupV0_lo_lo_hi_hi_lo_lo_hi;
  assign regroupV0_lo_lo_hi_hi_lo_lo_hi = _GEN_24;
  wire [63:0]        regroupV0_lo_lo_hi_hi_lo_lo_hi_5;
  assign regroupV0_lo_lo_hi_hi_lo_lo_hi_5 = _GEN_24;
  wire [63:0]        regroupV0_lo_lo_hi_hi_lo_lo_hi_10;
  assign regroupV0_lo_lo_hi_hi_lo_lo_hi_10 = _GEN_24;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_hi_hi_lo_lo_hi;
  assign slideAddressGen_slideMaskInput_lo_lo_hi_hi_lo_lo_hi = _GEN_24;
  wire [63:0]        selectReadStageMask_lo_lo_hi_hi_lo_lo_hi;
  assign selectReadStageMask_lo_lo_hi_hi_lo_lo_hi = _GEN_24;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_lo_lo_hi;
  assign maskSplit_maskSelect_lo_lo_hi_hi_lo_lo_hi = _GEN_24;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_lo_lo_hi_1;
  assign maskSplit_maskSelect_lo_lo_hi_hi_lo_lo_hi_1 = _GEN_24;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_lo_lo_hi_2;
  assign maskSplit_maskSelect_lo_lo_hi_hi_lo_lo_hi_2 = _GEN_24;
  wire [63:0]        maskForDestination_lo_lo_hi_hi_lo_lo_hi;
  assign maskForDestination_lo_lo_hi_hi_lo_lo_hi = _GEN_24;
  wire [127:0]       regroupV0_lo_lo_hi_hi_lo_lo = {regroupV0_lo_lo_hi_hi_lo_lo_hi, regroupV0_lo_lo_hi_hi_lo_lo_lo};
  wire [63:0]        _GEN_25 = {v0_53, v0_52};
  wire [63:0]        regroupV0_lo_lo_hi_hi_lo_hi_lo;
  assign regroupV0_lo_lo_hi_hi_lo_hi_lo = _GEN_25;
  wire [63:0]        regroupV0_lo_lo_hi_hi_lo_hi_lo_5;
  assign regroupV0_lo_lo_hi_hi_lo_hi_lo_5 = _GEN_25;
  wire [63:0]        regroupV0_lo_lo_hi_hi_lo_hi_lo_10;
  assign regroupV0_lo_lo_hi_hi_lo_hi_lo_10 = _GEN_25;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_hi_hi_lo_hi_lo;
  assign slideAddressGen_slideMaskInput_lo_lo_hi_hi_lo_hi_lo = _GEN_25;
  wire [63:0]        selectReadStageMask_lo_lo_hi_hi_lo_hi_lo;
  assign selectReadStageMask_lo_lo_hi_hi_lo_hi_lo = _GEN_25;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_lo_hi_lo;
  assign maskSplit_maskSelect_lo_lo_hi_hi_lo_hi_lo = _GEN_25;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_lo_hi_lo_1;
  assign maskSplit_maskSelect_lo_lo_hi_hi_lo_hi_lo_1 = _GEN_25;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_lo_hi_lo_2;
  assign maskSplit_maskSelect_lo_lo_hi_hi_lo_hi_lo_2 = _GEN_25;
  wire [63:0]        maskForDestination_lo_lo_hi_hi_lo_hi_lo;
  assign maskForDestination_lo_lo_hi_hi_lo_hi_lo = _GEN_25;
  wire [63:0]        _GEN_26 = {v0_55, v0_54};
  wire [63:0]        regroupV0_lo_lo_hi_hi_lo_hi_hi;
  assign regroupV0_lo_lo_hi_hi_lo_hi_hi = _GEN_26;
  wire [63:0]        regroupV0_lo_lo_hi_hi_lo_hi_hi_5;
  assign regroupV0_lo_lo_hi_hi_lo_hi_hi_5 = _GEN_26;
  wire [63:0]        regroupV0_lo_lo_hi_hi_lo_hi_hi_10;
  assign regroupV0_lo_lo_hi_hi_lo_hi_hi_10 = _GEN_26;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_hi_hi_lo_hi_hi;
  assign slideAddressGen_slideMaskInput_lo_lo_hi_hi_lo_hi_hi = _GEN_26;
  wire [63:0]        selectReadStageMask_lo_lo_hi_hi_lo_hi_hi;
  assign selectReadStageMask_lo_lo_hi_hi_lo_hi_hi = _GEN_26;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_lo_hi_hi;
  assign maskSplit_maskSelect_lo_lo_hi_hi_lo_hi_hi = _GEN_26;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_lo_hi_hi_1;
  assign maskSplit_maskSelect_lo_lo_hi_hi_lo_hi_hi_1 = _GEN_26;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_lo_hi_hi_2;
  assign maskSplit_maskSelect_lo_lo_hi_hi_lo_hi_hi_2 = _GEN_26;
  wire [63:0]        maskForDestination_lo_lo_hi_hi_lo_hi_hi;
  assign maskForDestination_lo_lo_hi_hi_lo_hi_hi = _GEN_26;
  wire [127:0]       regroupV0_lo_lo_hi_hi_lo_hi = {regroupV0_lo_lo_hi_hi_lo_hi_hi, regroupV0_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]       regroupV0_lo_lo_hi_hi_lo = {regroupV0_lo_lo_hi_hi_lo_hi, regroupV0_lo_lo_hi_hi_lo_lo};
  wire [63:0]        _GEN_27 = {v0_57, v0_56};
  wire [63:0]        regroupV0_lo_lo_hi_hi_hi_lo_lo;
  assign regroupV0_lo_lo_hi_hi_hi_lo_lo = _GEN_27;
  wire [63:0]        regroupV0_lo_lo_hi_hi_hi_lo_lo_5;
  assign regroupV0_lo_lo_hi_hi_hi_lo_lo_5 = _GEN_27;
  wire [63:0]        regroupV0_lo_lo_hi_hi_hi_lo_lo_10;
  assign regroupV0_lo_lo_hi_hi_hi_lo_lo_10 = _GEN_27;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_hi_hi_hi_lo_lo;
  assign slideAddressGen_slideMaskInput_lo_lo_hi_hi_hi_lo_lo = _GEN_27;
  wire [63:0]        selectReadStageMask_lo_lo_hi_hi_hi_lo_lo;
  assign selectReadStageMask_lo_lo_hi_hi_hi_lo_lo = _GEN_27;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_hi_lo_lo;
  assign maskSplit_maskSelect_lo_lo_hi_hi_hi_lo_lo = _GEN_27;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_hi_lo_lo_1;
  assign maskSplit_maskSelect_lo_lo_hi_hi_hi_lo_lo_1 = _GEN_27;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_hi_lo_lo_2;
  assign maskSplit_maskSelect_lo_lo_hi_hi_hi_lo_lo_2 = _GEN_27;
  wire [63:0]        maskForDestination_lo_lo_hi_hi_hi_lo_lo;
  assign maskForDestination_lo_lo_hi_hi_hi_lo_lo = _GEN_27;
  wire [63:0]        _GEN_28 = {v0_59, v0_58};
  wire [63:0]        regroupV0_lo_lo_hi_hi_hi_lo_hi;
  assign regroupV0_lo_lo_hi_hi_hi_lo_hi = _GEN_28;
  wire [63:0]        regroupV0_lo_lo_hi_hi_hi_lo_hi_5;
  assign regroupV0_lo_lo_hi_hi_hi_lo_hi_5 = _GEN_28;
  wire [63:0]        regroupV0_lo_lo_hi_hi_hi_lo_hi_10;
  assign regroupV0_lo_lo_hi_hi_hi_lo_hi_10 = _GEN_28;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_hi_hi_hi_lo_hi;
  assign slideAddressGen_slideMaskInput_lo_lo_hi_hi_hi_lo_hi = _GEN_28;
  wire [63:0]        selectReadStageMask_lo_lo_hi_hi_hi_lo_hi;
  assign selectReadStageMask_lo_lo_hi_hi_hi_lo_hi = _GEN_28;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_hi_lo_hi;
  assign maskSplit_maskSelect_lo_lo_hi_hi_hi_lo_hi = _GEN_28;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_hi_lo_hi_1;
  assign maskSplit_maskSelect_lo_lo_hi_hi_hi_lo_hi_1 = _GEN_28;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_hi_lo_hi_2;
  assign maskSplit_maskSelect_lo_lo_hi_hi_hi_lo_hi_2 = _GEN_28;
  wire [63:0]        maskForDestination_lo_lo_hi_hi_hi_lo_hi;
  assign maskForDestination_lo_lo_hi_hi_hi_lo_hi = _GEN_28;
  wire [127:0]       regroupV0_lo_lo_hi_hi_hi_lo = {regroupV0_lo_lo_hi_hi_hi_lo_hi, regroupV0_lo_lo_hi_hi_hi_lo_lo};
  wire [63:0]        _GEN_29 = {v0_61, v0_60};
  wire [63:0]        regroupV0_lo_lo_hi_hi_hi_hi_lo;
  assign regroupV0_lo_lo_hi_hi_hi_hi_lo = _GEN_29;
  wire [63:0]        regroupV0_lo_lo_hi_hi_hi_hi_lo_5;
  assign regroupV0_lo_lo_hi_hi_hi_hi_lo_5 = _GEN_29;
  wire [63:0]        regroupV0_lo_lo_hi_hi_hi_hi_lo_10;
  assign regroupV0_lo_lo_hi_hi_hi_hi_lo_10 = _GEN_29;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_hi_hi_hi_hi_lo;
  assign slideAddressGen_slideMaskInput_lo_lo_hi_hi_hi_hi_lo = _GEN_29;
  wire [63:0]        selectReadStageMask_lo_lo_hi_hi_hi_hi_lo;
  assign selectReadStageMask_lo_lo_hi_hi_hi_hi_lo = _GEN_29;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_hi_hi_lo;
  assign maskSplit_maskSelect_lo_lo_hi_hi_hi_hi_lo = _GEN_29;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_hi_hi_lo_1;
  assign maskSplit_maskSelect_lo_lo_hi_hi_hi_hi_lo_1 = _GEN_29;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_hi_hi_lo_2;
  assign maskSplit_maskSelect_lo_lo_hi_hi_hi_hi_lo_2 = _GEN_29;
  wire [63:0]        maskForDestination_lo_lo_hi_hi_hi_hi_lo;
  assign maskForDestination_lo_lo_hi_hi_hi_hi_lo = _GEN_29;
  wire [63:0]        _GEN_30 = {v0_63, v0_62};
  wire [63:0]        regroupV0_lo_lo_hi_hi_hi_hi_hi;
  assign regroupV0_lo_lo_hi_hi_hi_hi_hi = _GEN_30;
  wire [63:0]        regroupV0_lo_lo_hi_hi_hi_hi_hi_5;
  assign regroupV0_lo_lo_hi_hi_hi_hi_hi_5 = _GEN_30;
  wire [63:0]        regroupV0_lo_lo_hi_hi_hi_hi_hi_10;
  assign regroupV0_lo_lo_hi_hi_hi_hi_hi_10 = _GEN_30;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_hi_hi_hi_hi_hi;
  assign slideAddressGen_slideMaskInput_lo_lo_hi_hi_hi_hi_hi = _GEN_30;
  wire [63:0]        selectReadStageMask_lo_lo_hi_hi_hi_hi_hi;
  assign selectReadStageMask_lo_lo_hi_hi_hi_hi_hi = _GEN_30;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_hi_hi_hi;
  assign maskSplit_maskSelect_lo_lo_hi_hi_hi_hi_hi = _GEN_30;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_hi_hi_hi_1;
  assign maskSplit_maskSelect_lo_lo_hi_hi_hi_hi_hi_1 = _GEN_30;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_hi_hi_hi_2;
  assign maskSplit_maskSelect_lo_lo_hi_hi_hi_hi_hi_2 = _GEN_30;
  wire [63:0]        maskForDestination_lo_lo_hi_hi_hi_hi_hi;
  assign maskForDestination_lo_lo_hi_hi_hi_hi_hi = _GEN_30;
  wire [127:0]       regroupV0_lo_lo_hi_hi_hi_hi = {regroupV0_lo_lo_hi_hi_hi_hi_hi, regroupV0_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]       regroupV0_lo_lo_hi_hi_hi = {regroupV0_lo_lo_hi_hi_hi_hi, regroupV0_lo_lo_hi_hi_hi_lo};
  wire [511:0]       regroupV0_lo_lo_hi_hi = {regroupV0_lo_lo_hi_hi_hi, regroupV0_lo_lo_hi_hi_lo};
  wire [1023:0]      regroupV0_lo_lo_hi = {regroupV0_lo_lo_hi_hi, regroupV0_lo_lo_hi_lo};
  wire [2047:0]      regroupV0_lo_lo = {regroupV0_lo_lo_hi, regroupV0_lo_lo_lo};
  wire [63:0]        _GEN_31 = {v0_65, v0_64};
  wire [63:0]        regroupV0_lo_hi_lo_lo_lo_lo_lo;
  assign regroupV0_lo_hi_lo_lo_lo_lo_lo = _GEN_31;
  wire [63:0]        regroupV0_lo_hi_lo_lo_lo_lo_lo_5;
  assign regroupV0_lo_hi_lo_lo_lo_lo_lo_5 = _GEN_31;
  wire [63:0]        regroupV0_lo_hi_lo_lo_lo_lo_lo_10;
  assign regroupV0_lo_hi_lo_lo_lo_lo_lo_10 = _GEN_31;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_lo_lo_lo_lo_lo;
  assign slideAddressGen_slideMaskInput_lo_hi_lo_lo_lo_lo_lo = _GEN_31;
  wire [63:0]        selectReadStageMask_lo_hi_lo_lo_lo_lo_lo;
  assign selectReadStageMask_lo_hi_lo_lo_lo_lo_lo = _GEN_31;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_lo_lo_lo;
  assign maskSplit_maskSelect_lo_hi_lo_lo_lo_lo_lo = _GEN_31;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_lo_lo_lo_1;
  assign maskSplit_maskSelect_lo_hi_lo_lo_lo_lo_lo_1 = _GEN_31;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_lo_lo_lo_2;
  assign maskSplit_maskSelect_lo_hi_lo_lo_lo_lo_lo_2 = _GEN_31;
  wire [63:0]        maskForDestination_lo_hi_lo_lo_lo_lo_lo;
  assign maskForDestination_lo_hi_lo_lo_lo_lo_lo = _GEN_31;
  wire [63:0]        _GEN_32 = {v0_67, v0_66};
  wire [63:0]        regroupV0_lo_hi_lo_lo_lo_lo_hi;
  assign regroupV0_lo_hi_lo_lo_lo_lo_hi = _GEN_32;
  wire [63:0]        regroupV0_lo_hi_lo_lo_lo_lo_hi_5;
  assign regroupV0_lo_hi_lo_lo_lo_lo_hi_5 = _GEN_32;
  wire [63:0]        regroupV0_lo_hi_lo_lo_lo_lo_hi_10;
  assign regroupV0_lo_hi_lo_lo_lo_lo_hi_10 = _GEN_32;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_lo_lo_lo_lo_hi;
  assign slideAddressGen_slideMaskInput_lo_hi_lo_lo_lo_lo_hi = _GEN_32;
  wire [63:0]        selectReadStageMask_lo_hi_lo_lo_lo_lo_hi;
  assign selectReadStageMask_lo_hi_lo_lo_lo_lo_hi = _GEN_32;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_lo_lo_hi;
  assign maskSplit_maskSelect_lo_hi_lo_lo_lo_lo_hi = _GEN_32;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_lo_lo_hi_1;
  assign maskSplit_maskSelect_lo_hi_lo_lo_lo_lo_hi_1 = _GEN_32;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_lo_lo_hi_2;
  assign maskSplit_maskSelect_lo_hi_lo_lo_lo_lo_hi_2 = _GEN_32;
  wire [63:0]        maskForDestination_lo_hi_lo_lo_lo_lo_hi;
  assign maskForDestination_lo_hi_lo_lo_lo_lo_hi = _GEN_32;
  wire [127:0]       regroupV0_lo_hi_lo_lo_lo_lo = {regroupV0_lo_hi_lo_lo_lo_lo_hi, regroupV0_lo_hi_lo_lo_lo_lo_lo};
  wire [63:0]        _GEN_33 = {v0_69, v0_68};
  wire [63:0]        regroupV0_lo_hi_lo_lo_lo_hi_lo;
  assign regroupV0_lo_hi_lo_lo_lo_hi_lo = _GEN_33;
  wire [63:0]        regroupV0_lo_hi_lo_lo_lo_hi_lo_5;
  assign regroupV0_lo_hi_lo_lo_lo_hi_lo_5 = _GEN_33;
  wire [63:0]        regroupV0_lo_hi_lo_lo_lo_hi_lo_10;
  assign regroupV0_lo_hi_lo_lo_lo_hi_lo_10 = _GEN_33;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_lo_lo_lo_hi_lo;
  assign slideAddressGen_slideMaskInput_lo_hi_lo_lo_lo_hi_lo = _GEN_33;
  wire [63:0]        selectReadStageMask_lo_hi_lo_lo_lo_hi_lo;
  assign selectReadStageMask_lo_hi_lo_lo_lo_hi_lo = _GEN_33;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_lo_hi_lo;
  assign maskSplit_maskSelect_lo_hi_lo_lo_lo_hi_lo = _GEN_33;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_lo_hi_lo_1;
  assign maskSplit_maskSelect_lo_hi_lo_lo_lo_hi_lo_1 = _GEN_33;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_lo_hi_lo_2;
  assign maskSplit_maskSelect_lo_hi_lo_lo_lo_hi_lo_2 = _GEN_33;
  wire [63:0]        maskForDestination_lo_hi_lo_lo_lo_hi_lo;
  assign maskForDestination_lo_hi_lo_lo_lo_hi_lo = _GEN_33;
  wire [63:0]        _GEN_34 = {v0_71, v0_70};
  wire [63:0]        regroupV0_lo_hi_lo_lo_lo_hi_hi;
  assign regroupV0_lo_hi_lo_lo_lo_hi_hi = _GEN_34;
  wire [63:0]        regroupV0_lo_hi_lo_lo_lo_hi_hi_5;
  assign regroupV0_lo_hi_lo_lo_lo_hi_hi_5 = _GEN_34;
  wire [63:0]        regroupV0_lo_hi_lo_lo_lo_hi_hi_10;
  assign regroupV0_lo_hi_lo_lo_lo_hi_hi_10 = _GEN_34;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_lo_lo_lo_hi_hi;
  assign slideAddressGen_slideMaskInput_lo_hi_lo_lo_lo_hi_hi = _GEN_34;
  wire [63:0]        selectReadStageMask_lo_hi_lo_lo_lo_hi_hi;
  assign selectReadStageMask_lo_hi_lo_lo_lo_hi_hi = _GEN_34;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_lo_hi_hi;
  assign maskSplit_maskSelect_lo_hi_lo_lo_lo_hi_hi = _GEN_34;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_lo_hi_hi_1;
  assign maskSplit_maskSelect_lo_hi_lo_lo_lo_hi_hi_1 = _GEN_34;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_lo_hi_hi_2;
  assign maskSplit_maskSelect_lo_hi_lo_lo_lo_hi_hi_2 = _GEN_34;
  wire [63:0]        maskForDestination_lo_hi_lo_lo_lo_hi_hi;
  assign maskForDestination_lo_hi_lo_lo_lo_hi_hi = _GEN_34;
  wire [127:0]       regroupV0_lo_hi_lo_lo_lo_hi = {regroupV0_lo_hi_lo_lo_lo_hi_hi, regroupV0_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]       regroupV0_lo_hi_lo_lo_lo = {regroupV0_lo_hi_lo_lo_lo_hi, regroupV0_lo_hi_lo_lo_lo_lo};
  wire [63:0]        _GEN_35 = {v0_73, v0_72};
  wire [63:0]        regroupV0_lo_hi_lo_lo_hi_lo_lo;
  assign regroupV0_lo_hi_lo_lo_hi_lo_lo = _GEN_35;
  wire [63:0]        regroupV0_lo_hi_lo_lo_hi_lo_lo_5;
  assign regroupV0_lo_hi_lo_lo_hi_lo_lo_5 = _GEN_35;
  wire [63:0]        regroupV0_lo_hi_lo_lo_hi_lo_lo_10;
  assign regroupV0_lo_hi_lo_lo_hi_lo_lo_10 = _GEN_35;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_lo_lo_hi_lo_lo;
  assign slideAddressGen_slideMaskInput_lo_hi_lo_lo_hi_lo_lo = _GEN_35;
  wire [63:0]        selectReadStageMask_lo_hi_lo_lo_hi_lo_lo;
  assign selectReadStageMask_lo_hi_lo_lo_hi_lo_lo = _GEN_35;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_hi_lo_lo;
  assign maskSplit_maskSelect_lo_hi_lo_lo_hi_lo_lo = _GEN_35;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_hi_lo_lo_1;
  assign maskSplit_maskSelect_lo_hi_lo_lo_hi_lo_lo_1 = _GEN_35;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_hi_lo_lo_2;
  assign maskSplit_maskSelect_lo_hi_lo_lo_hi_lo_lo_2 = _GEN_35;
  wire [63:0]        maskForDestination_lo_hi_lo_lo_hi_lo_lo;
  assign maskForDestination_lo_hi_lo_lo_hi_lo_lo = _GEN_35;
  wire [63:0]        _GEN_36 = {v0_75, v0_74};
  wire [63:0]        regroupV0_lo_hi_lo_lo_hi_lo_hi;
  assign regroupV0_lo_hi_lo_lo_hi_lo_hi = _GEN_36;
  wire [63:0]        regroupV0_lo_hi_lo_lo_hi_lo_hi_5;
  assign regroupV0_lo_hi_lo_lo_hi_lo_hi_5 = _GEN_36;
  wire [63:0]        regroupV0_lo_hi_lo_lo_hi_lo_hi_10;
  assign regroupV0_lo_hi_lo_lo_hi_lo_hi_10 = _GEN_36;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_lo_lo_hi_lo_hi;
  assign slideAddressGen_slideMaskInput_lo_hi_lo_lo_hi_lo_hi = _GEN_36;
  wire [63:0]        selectReadStageMask_lo_hi_lo_lo_hi_lo_hi;
  assign selectReadStageMask_lo_hi_lo_lo_hi_lo_hi = _GEN_36;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_hi_lo_hi;
  assign maskSplit_maskSelect_lo_hi_lo_lo_hi_lo_hi = _GEN_36;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_hi_lo_hi_1;
  assign maskSplit_maskSelect_lo_hi_lo_lo_hi_lo_hi_1 = _GEN_36;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_hi_lo_hi_2;
  assign maskSplit_maskSelect_lo_hi_lo_lo_hi_lo_hi_2 = _GEN_36;
  wire [63:0]        maskForDestination_lo_hi_lo_lo_hi_lo_hi;
  assign maskForDestination_lo_hi_lo_lo_hi_lo_hi = _GEN_36;
  wire [127:0]       regroupV0_lo_hi_lo_lo_hi_lo = {regroupV0_lo_hi_lo_lo_hi_lo_hi, regroupV0_lo_hi_lo_lo_hi_lo_lo};
  wire [63:0]        _GEN_37 = {v0_77, v0_76};
  wire [63:0]        regroupV0_lo_hi_lo_lo_hi_hi_lo;
  assign regroupV0_lo_hi_lo_lo_hi_hi_lo = _GEN_37;
  wire [63:0]        regroupV0_lo_hi_lo_lo_hi_hi_lo_5;
  assign regroupV0_lo_hi_lo_lo_hi_hi_lo_5 = _GEN_37;
  wire [63:0]        regroupV0_lo_hi_lo_lo_hi_hi_lo_10;
  assign regroupV0_lo_hi_lo_lo_hi_hi_lo_10 = _GEN_37;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_lo_lo_hi_hi_lo;
  assign slideAddressGen_slideMaskInput_lo_hi_lo_lo_hi_hi_lo = _GEN_37;
  wire [63:0]        selectReadStageMask_lo_hi_lo_lo_hi_hi_lo;
  assign selectReadStageMask_lo_hi_lo_lo_hi_hi_lo = _GEN_37;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_hi_hi_lo;
  assign maskSplit_maskSelect_lo_hi_lo_lo_hi_hi_lo = _GEN_37;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_hi_hi_lo_1;
  assign maskSplit_maskSelect_lo_hi_lo_lo_hi_hi_lo_1 = _GEN_37;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_hi_hi_lo_2;
  assign maskSplit_maskSelect_lo_hi_lo_lo_hi_hi_lo_2 = _GEN_37;
  wire [63:0]        maskForDestination_lo_hi_lo_lo_hi_hi_lo;
  assign maskForDestination_lo_hi_lo_lo_hi_hi_lo = _GEN_37;
  wire [63:0]        _GEN_38 = {v0_79, v0_78};
  wire [63:0]        regroupV0_lo_hi_lo_lo_hi_hi_hi;
  assign regroupV0_lo_hi_lo_lo_hi_hi_hi = _GEN_38;
  wire [63:0]        regroupV0_lo_hi_lo_lo_hi_hi_hi_5;
  assign regroupV0_lo_hi_lo_lo_hi_hi_hi_5 = _GEN_38;
  wire [63:0]        regroupV0_lo_hi_lo_lo_hi_hi_hi_10;
  assign regroupV0_lo_hi_lo_lo_hi_hi_hi_10 = _GEN_38;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_lo_lo_hi_hi_hi;
  assign slideAddressGen_slideMaskInput_lo_hi_lo_lo_hi_hi_hi = _GEN_38;
  wire [63:0]        selectReadStageMask_lo_hi_lo_lo_hi_hi_hi;
  assign selectReadStageMask_lo_hi_lo_lo_hi_hi_hi = _GEN_38;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_hi_hi_hi;
  assign maskSplit_maskSelect_lo_hi_lo_lo_hi_hi_hi = _GEN_38;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_hi_hi_hi_1;
  assign maskSplit_maskSelect_lo_hi_lo_lo_hi_hi_hi_1 = _GEN_38;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_hi_hi_hi_2;
  assign maskSplit_maskSelect_lo_hi_lo_lo_hi_hi_hi_2 = _GEN_38;
  wire [63:0]        maskForDestination_lo_hi_lo_lo_hi_hi_hi;
  assign maskForDestination_lo_hi_lo_lo_hi_hi_hi = _GEN_38;
  wire [127:0]       regroupV0_lo_hi_lo_lo_hi_hi = {regroupV0_lo_hi_lo_lo_hi_hi_hi, regroupV0_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]       regroupV0_lo_hi_lo_lo_hi = {regroupV0_lo_hi_lo_lo_hi_hi, regroupV0_lo_hi_lo_lo_hi_lo};
  wire [511:0]       regroupV0_lo_hi_lo_lo = {regroupV0_lo_hi_lo_lo_hi, regroupV0_lo_hi_lo_lo_lo};
  wire [63:0]        _GEN_39 = {v0_81, v0_80};
  wire [63:0]        regroupV0_lo_hi_lo_hi_lo_lo_lo;
  assign regroupV0_lo_hi_lo_hi_lo_lo_lo = _GEN_39;
  wire [63:0]        regroupV0_lo_hi_lo_hi_lo_lo_lo_5;
  assign regroupV0_lo_hi_lo_hi_lo_lo_lo_5 = _GEN_39;
  wire [63:0]        regroupV0_lo_hi_lo_hi_lo_lo_lo_10;
  assign regroupV0_lo_hi_lo_hi_lo_lo_lo_10 = _GEN_39;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_lo_hi_lo_lo_lo;
  assign slideAddressGen_slideMaskInput_lo_hi_lo_hi_lo_lo_lo = _GEN_39;
  wire [63:0]        selectReadStageMask_lo_hi_lo_hi_lo_lo_lo;
  assign selectReadStageMask_lo_hi_lo_hi_lo_lo_lo = _GEN_39;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_lo_lo_lo;
  assign maskSplit_maskSelect_lo_hi_lo_hi_lo_lo_lo = _GEN_39;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_lo_lo_lo_1;
  assign maskSplit_maskSelect_lo_hi_lo_hi_lo_lo_lo_1 = _GEN_39;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_lo_lo_lo_2;
  assign maskSplit_maskSelect_lo_hi_lo_hi_lo_lo_lo_2 = _GEN_39;
  wire [63:0]        maskForDestination_lo_hi_lo_hi_lo_lo_lo;
  assign maskForDestination_lo_hi_lo_hi_lo_lo_lo = _GEN_39;
  wire [63:0]        _GEN_40 = {v0_83, v0_82};
  wire [63:0]        regroupV0_lo_hi_lo_hi_lo_lo_hi;
  assign regroupV0_lo_hi_lo_hi_lo_lo_hi = _GEN_40;
  wire [63:0]        regroupV0_lo_hi_lo_hi_lo_lo_hi_5;
  assign regroupV0_lo_hi_lo_hi_lo_lo_hi_5 = _GEN_40;
  wire [63:0]        regroupV0_lo_hi_lo_hi_lo_lo_hi_10;
  assign regroupV0_lo_hi_lo_hi_lo_lo_hi_10 = _GEN_40;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_lo_hi_lo_lo_hi;
  assign slideAddressGen_slideMaskInput_lo_hi_lo_hi_lo_lo_hi = _GEN_40;
  wire [63:0]        selectReadStageMask_lo_hi_lo_hi_lo_lo_hi;
  assign selectReadStageMask_lo_hi_lo_hi_lo_lo_hi = _GEN_40;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_lo_lo_hi;
  assign maskSplit_maskSelect_lo_hi_lo_hi_lo_lo_hi = _GEN_40;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_lo_lo_hi_1;
  assign maskSplit_maskSelect_lo_hi_lo_hi_lo_lo_hi_1 = _GEN_40;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_lo_lo_hi_2;
  assign maskSplit_maskSelect_lo_hi_lo_hi_lo_lo_hi_2 = _GEN_40;
  wire [63:0]        maskForDestination_lo_hi_lo_hi_lo_lo_hi;
  assign maskForDestination_lo_hi_lo_hi_lo_lo_hi = _GEN_40;
  wire [127:0]       regroupV0_lo_hi_lo_hi_lo_lo = {regroupV0_lo_hi_lo_hi_lo_lo_hi, regroupV0_lo_hi_lo_hi_lo_lo_lo};
  wire [63:0]        _GEN_41 = {v0_85, v0_84};
  wire [63:0]        regroupV0_lo_hi_lo_hi_lo_hi_lo;
  assign regroupV0_lo_hi_lo_hi_lo_hi_lo = _GEN_41;
  wire [63:0]        regroupV0_lo_hi_lo_hi_lo_hi_lo_5;
  assign regroupV0_lo_hi_lo_hi_lo_hi_lo_5 = _GEN_41;
  wire [63:0]        regroupV0_lo_hi_lo_hi_lo_hi_lo_10;
  assign regroupV0_lo_hi_lo_hi_lo_hi_lo_10 = _GEN_41;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_lo_hi_lo_hi_lo;
  assign slideAddressGen_slideMaskInput_lo_hi_lo_hi_lo_hi_lo = _GEN_41;
  wire [63:0]        selectReadStageMask_lo_hi_lo_hi_lo_hi_lo;
  assign selectReadStageMask_lo_hi_lo_hi_lo_hi_lo = _GEN_41;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_lo_hi_lo;
  assign maskSplit_maskSelect_lo_hi_lo_hi_lo_hi_lo = _GEN_41;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_lo_hi_lo_1;
  assign maskSplit_maskSelect_lo_hi_lo_hi_lo_hi_lo_1 = _GEN_41;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_lo_hi_lo_2;
  assign maskSplit_maskSelect_lo_hi_lo_hi_lo_hi_lo_2 = _GEN_41;
  wire [63:0]        maskForDestination_lo_hi_lo_hi_lo_hi_lo;
  assign maskForDestination_lo_hi_lo_hi_lo_hi_lo = _GEN_41;
  wire [63:0]        _GEN_42 = {v0_87, v0_86};
  wire [63:0]        regroupV0_lo_hi_lo_hi_lo_hi_hi;
  assign regroupV0_lo_hi_lo_hi_lo_hi_hi = _GEN_42;
  wire [63:0]        regroupV0_lo_hi_lo_hi_lo_hi_hi_5;
  assign regroupV0_lo_hi_lo_hi_lo_hi_hi_5 = _GEN_42;
  wire [63:0]        regroupV0_lo_hi_lo_hi_lo_hi_hi_10;
  assign regroupV0_lo_hi_lo_hi_lo_hi_hi_10 = _GEN_42;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_lo_hi_lo_hi_hi;
  assign slideAddressGen_slideMaskInput_lo_hi_lo_hi_lo_hi_hi = _GEN_42;
  wire [63:0]        selectReadStageMask_lo_hi_lo_hi_lo_hi_hi;
  assign selectReadStageMask_lo_hi_lo_hi_lo_hi_hi = _GEN_42;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_lo_hi_hi;
  assign maskSplit_maskSelect_lo_hi_lo_hi_lo_hi_hi = _GEN_42;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_lo_hi_hi_1;
  assign maskSplit_maskSelect_lo_hi_lo_hi_lo_hi_hi_1 = _GEN_42;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_lo_hi_hi_2;
  assign maskSplit_maskSelect_lo_hi_lo_hi_lo_hi_hi_2 = _GEN_42;
  wire [63:0]        maskForDestination_lo_hi_lo_hi_lo_hi_hi;
  assign maskForDestination_lo_hi_lo_hi_lo_hi_hi = _GEN_42;
  wire [127:0]       regroupV0_lo_hi_lo_hi_lo_hi = {regroupV0_lo_hi_lo_hi_lo_hi_hi, regroupV0_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]       regroupV0_lo_hi_lo_hi_lo = {regroupV0_lo_hi_lo_hi_lo_hi, regroupV0_lo_hi_lo_hi_lo_lo};
  wire [63:0]        _GEN_43 = {v0_89, v0_88};
  wire [63:0]        regroupV0_lo_hi_lo_hi_hi_lo_lo;
  assign regroupV0_lo_hi_lo_hi_hi_lo_lo = _GEN_43;
  wire [63:0]        regroupV0_lo_hi_lo_hi_hi_lo_lo_5;
  assign regroupV0_lo_hi_lo_hi_hi_lo_lo_5 = _GEN_43;
  wire [63:0]        regroupV0_lo_hi_lo_hi_hi_lo_lo_10;
  assign regroupV0_lo_hi_lo_hi_hi_lo_lo_10 = _GEN_43;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_lo_hi_hi_lo_lo;
  assign slideAddressGen_slideMaskInput_lo_hi_lo_hi_hi_lo_lo = _GEN_43;
  wire [63:0]        selectReadStageMask_lo_hi_lo_hi_hi_lo_lo;
  assign selectReadStageMask_lo_hi_lo_hi_hi_lo_lo = _GEN_43;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_hi_lo_lo;
  assign maskSplit_maskSelect_lo_hi_lo_hi_hi_lo_lo = _GEN_43;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_hi_lo_lo_1;
  assign maskSplit_maskSelect_lo_hi_lo_hi_hi_lo_lo_1 = _GEN_43;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_hi_lo_lo_2;
  assign maskSplit_maskSelect_lo_hi_lo_hi_hi_lo_lo_2 = _GEN_43;
  wire [63:0]        maskForDestination_lo_hi_lo_hi_hi_lo_lo;
  assign maskForDestination_lo_hi_lo_hi_hi_lo_lo = _GEN_43;
  wire [63:0]        _GEN_44 = {v0_91, v0_90};
  wire [63:0]        regroupV0_lo_hi_lo_hi_hi_lo_hi;
  assign regroupV0_lo_hi_lo_hi_hi_lo_hi = _GEN_44;
  wire [63:0]        regroupV0_lo_hi_lo_hi_hi_lo_hi_5;
  assign regroupV0_lo_hi_lo_hi_hi_lo_hi_5 = _GEN_44;
  wire [63:0]        regroupV0_lo_hi_lo_hi_hi_lo_hi_10;
  assign regroupV0_lo_hi_lo_hi_hi_lo_hi_10 = _GEN_44;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_lo_hi_hi_lo_hi;
  assign slideAddressGen_slideMaskInput_lo_hi_lo_hi_hi_lo_hi = _GEN_44;
  wire [63:0]        selectReadStageMask_lo_hi_lo_hi_hi_lo_hi;
  assign selectReadStageMask_lo_hi_lo_hi_hi_lo_hi = _GEN_44;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_hi_lo_hi;
  assign maskSplit_maskSelect_lo_hi_lo_hi_hi_lo_hi = _GEN_44;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_hi_lo_hi_1;
  assign maskSplit_maskSelect_lo_hi_lo_hi_hi_lo_hi_1 = _GEN_44;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_hi_lo_hi_2;
  assign maskSplit_maskSelect_lo_hi_lo_hi_hi_lo_hi_2 = _GEN_44;
  wire [63:0]        maskForDestination_lo_hi_lo_hi_hi_lo_hi;
  assign maskForDestination_lo_hi_lo_hi_hi_lo_hi = _GEN_44;
  wire [127:0]       regroupV0_lo_hi_lo_hi_hi_lo = {regroupV0_lo_hi_lo_hi_hi_lo_hi, regroupV0_lo_hi_lo_hi_hi_lo_lo};
  wire [63:0]        _GEN_45 = {v0_93, v0_92};
  wire [63:0]        regroupV0_lo_hi_lo_hi_hi_hi_lo;
  assign regroupV0_lo_hi_lo_hi_hi_hi_lo = _GEN_45;
  wire [63:0]        regroupV0_lo_hi_lo_hi_hi_hi_lo_5;
  assign regroupV0_lo_hi_lo_hi_hi_hi_lo_5 = _GEN_45;
  wire [63:0]        regroupV0_lo_hi_lo_hi_hi_hi_lo_10;
  assign regroupV0_lo_hi_lo_hi_hi_hi_lo_10 = _GEN_45;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_lo_hi_hi_hi_lo;
  assign slideAddressGen_slideMaskInput_lo_hi_lo_hi_hi_hi_lo = _GEN_45;
  wire [63:0]        selectReadStageMask_lo_hi_lo_hi_hi_hi_lo;
  assign selectReadStageMask_lo_hi_lo_hi_hi_hi_lo = _GEN_45;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_hi_hi_lo;
  assign maskSplit_maskSelect_lo_hi_lo_hi_hi_hi_lo = _GEN_45;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_hi_hi_lo_1;
  assign maskSplit_maskSelect_lo_hi_lo_hi_hi_hi_lo_1 = _GEN_45;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_hi_hi_lo_2;
  assign maskSplit_maskSelect_lo_hi_lo_hi_hi_hi_lo_2 = _GEN_45;
  wire [63:0]        maskForDestination_lo_hi_lo_hi_hi_hi_lo;
  assign maskForDestination_lo_hi_lo_hi_hi_hi_lo = _GEN_45;
  wire [63:0]        _GEN_46 = {v0_95, v0_94};
  wire [63:0]        regroupV0_lo_hi_lo_hi_hi_hi_hi;
  assign regroupV0_lo_hi_lo_hi_hi_hi_hi = _GEN_46;
  wire [63:0]        regroupV0_lo_hi_lo_hi_hi_hi_hi_5;
  assign regroupV0_lo_hi_lo_hi_hi_hi_hi_5 = _GEN_46;
  wire [63:0]        regroupV0_lo_hi_lo_hi_hi_hi_hi_10;
  assign regroupV0_lo_hi_lo_hi_hi_hi_hi_10 = _GEN_46;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_lo_hi_hi_hi_hi;
  assign slideAddressGen_slideMaskInput_lo_hi_lo_hi_hi_hi_hi = _GEN_46;
  wire [63:0]        selectReadStageMask_lo_hi_lo_hi_hi_hi_hi;
  assign selectReadStageMask_lo_hi_lo_hi_hi_hi_hi = _GEN_46;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_hi_hi_hi;
  assign maskSplit_maskSelect_lo_hi_lo_hi_hi_hi_hi = _GEN_46;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_hi_hi_hi_1;
  assign maskSplit_maskSelect_lo_hi_lo_hi_hi_hi_hi_1 = _GEN_46;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_hi_hi_hi_2;
  assign maskSplit_maskSelect_lo_hi_lo_hi_hi_hi_hi_2 = _GEN_46;
  wire [63:0]        maskForDestination_lo_hi_lo_hi_hi_hi_hi;
  assign maskForDestination_lo_hi_lo_hi_hi_hi_hi = _GEN_46;
  wire [127:0]       regroupV0_lo_hi_lo_hi_hi_hi = {regroupV0_lo_hi_lo_hi_hi_hi_hi, regroupV0_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]       regroupV0_lo_hi_lo_hi_hi = {regroupV0_lo_hi_lo_hi_hi_hi, regroupV0_lo_hi_lo_hi_hi_lo};
  wire [511:0]       regroupV0_lo_hi_lo_hi = {regroupV0_lo_hi_lo_hi_hi, regroupV0_lo_hi_lo_hi_lo};
  wire [1023:0]      regroupV0_lo_hi_lo = {regroupV0_lo_hi_lo_hi, regroupV0_lo_hi_lo_lo};
  wire [63:0]        _GEN_47 = {v0_97, v0_96};
  wire [63:0]        regroupV0_lo_hi_hi_lo_lo_lo_lo;
  assign regroupV0_lo_hi_hi_lo_lo_lo_lo = _GEN_47;
  wire [63:0]        regroupV0_lo_hi_hi_lo_lo_lo_lo_5;
  assign regroupV0_lo_hi_hi_lo_lo_lo_lo_5 = _GEN_47;
  wire [63:0]        regroupV0_lo_hi_hi_lo_lo_lo_lo_10;
  assign regroupV0_lo_hi_hi_lo_lo_lo_lo_10 = _GEN_47;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_hi_lo_lo_lo_lo;
  assign slideAddressGen_slideMaskInput_lo_hi_hi_lo_lo_lo_lo = _GEN_47;
  wire [63:0]        selectReadStageMask_lo_hi_hi_lo_lo_lo_lo;
  assign selectReadStageMask_lo_hi_hi_lo_lo_lo_lo = _GEN_47;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_lo_lo_lo;
  assign maskSplit_maskSelect_lo_hi_hi_lo_lo_lo_lo = _GEN_47;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_lo_lo_lo_1;
  assign maskSplit_maskSelect_lo_hi_hi_lo_lo_lo_lo_1 = _GEN_47;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_lo_lo_lo_2;
  assign maskSplit_maskSelect_lo_hi_hi_lo_lo_lo_lo_2 = _GEN_47;
  wire [63:0]        maskForDestination_lo_hi_hi_lo_lo_lo_lo;
  assign maskForDestination_lo_hi_hi_lo_lo_lo_lo = _GEN_47;
  wire [63:0]        _GEN_48 = {v0_99, v0_98};
  wire [63:0]        regroupV0_lo_hi_hi_lo_lo_lo_hi;
  assign regroupV0_lo_hi_hi_lo_lo_lo_hi = _GEN_48;
  wire [63:0]        regroupV0_lo_hi_hi_lo_lo_lo_hi_5;
  assign regroupV0_lo_hi_hi_lo_lo_lo_hi_5 = _GEN_48;
  wire [63:0]        regroupV0_lo_hi_hi_lo_lo_lo_hi_10;
  assign regroupV0_lo_hi_hi_lo_lo_lo_hi_10 = _GEN_48;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_hi_lo_lo_lo_hi;
  assign slideAddressGen_slideMaskInput_lo_hi_hi_lo_lo_lo_hi = _GEN_48;
  wire [63:0]        selectReadStageMask_lo_hi_hi_lo_lo_lo_hi;
  assign selectReadStageMask_lo_hi_hi_lo_lo_lo_hi = _GEN_48;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_lo_lo_hi;
  assign maskSplit_maskSelect_lo_hi_hi_lo_lo_lo_hi = _GEN_48;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_lo_lo_hi_1;
  assign maskSplit_maskSelect_lo_hi_hi_lo_lo_lo_hi_1 = _GEN_48;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_lo_lo_hi_2;
  assign maskSplit_maskSelect_lo_hi_hi_lo_lo_lo_hi_2 = _GEN_48;
  wire [63:0]        maskForDestination_lo_hi_hi_lo_lo_lo_hi;
  assign maskForDestination_lo_hi_hi_lo_lo_lo_hi = _GEN_48;
  wire [127:0]       regroupV0_lo_hi_hi_lo_lo_lo = {regroupV0_lo_hi_hi_lo_lo_lo_hi, regroupV0_lo_hi_hi_lo_lo_lo_lo};
  wire [63:0]        _GEN_49 = {v0_101, v0_100};
  wire [63:0]        regroupV0_lo_hi_hi_lo_lo_hi_lo;
  assign regroupV0_lo_hi_hi_lo_lo_hi_lo = _GEN_49;
  wire [63:0]        regroupV0_lo_hi_hi_lo_lo_hi_lo_5;
  assign regroupV0_lo_hi_hi_lo_lo_hi_lo_5 = _GEN_49;
  wire [63:0]        regroupV0_lo_hi_hi_lo_lo_hi_lo_10;
  assign regroupV0_lo_hi_hi_lo_lo_hi_lo_10 = _GEN_49;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_hi_lo_lo_hi_lo;
  assign slideAddressGen_slideMaskInput_lo_hi_hi_lo_lo_hi_lo = _GEN_49;
  wire [63:0]        selectReadStageMask_lo_hi_hi_lo_lo_hi_lo;
  assign selectReadStageMask_lo_hi_hi_lo_lo_hi_lo = _GEN_49;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_lo_hi_lo;
  assign maskSplit_maskSelect_lo_hi_hi_lo_lo_hi_lo = _GEN_49;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_lo_hi_lo_1;
  assign maskSplit_maskSelect_lo_hi_hi_lo_lo_hi_lo_1 = _GEN_49;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_lo_hi_lo_2;
  assign maskSplit_maskSelect_lo_hi_hi_lo_lo_hi_lo_2 = _GEN_49;
  wire [63:0]        maskForDestination_lo_hi_hi_lo_lo_hi_lo;
  assign maskForDestination_lo_hi_hi_lo_lo_hi_lo = _GEN_49;
  wire [63:0]        _GEN_50 = {v0_103, v0_102};
  wire [63:0]        regroupV0_lo_hi_hi_lo_lo_hi_hi;
  assign regroupV0_lo_hi_hi_lo_lo_hi_hi = _GEN_50;
  wire [63:0]        regroupV0_lo_hi_hi_lo_lo_hi_hi_5;
  assign regroupV0_lo_hi_hi_lo_lo_hi_hi_5 = _GEN_50;
  wire [63:0]        regroupV0_lo_hi_hi_lo_lo_hi_hi_10;
  assign regroupV0_lo_hi_hi_lo_lo_hi_hi_10 = _GEN_50;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_hi_lo_lo_hi_hi;
  assign slideAddressGen_slideMaskInput_lo_hi_hi_lo_lo_hi_hi = _GEN_50;
  wire [63:0]        selectReadStageMask_lo_hi_hi_lo_lo_hi_hi;
  assign selectReadStageMask_lo_hi_hi_lo_lo_hi_hi = _GEN_50;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_lo_hi_hi;
  assign maskSplit_maskSelect_lo_hi_hi_lo_lo_hi_hi = _GEN_50;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_lo_hi_hi_1;
  assign maskSplit_maskSelect_lo_hi_hi_lo_lo_hi_hi_1 = _GEN_50;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_lo_hi_hi_2;
  assign maskSplit_maskSelect_lo_hi_hi_lo_lo_hi_hi_2 = _GEN_50;
  wire [63:0]        maskForDestination_lo_hi_hi_lo_lo_hi_hi;
  assign maskForDestination_lo_hi_hi_lo_lo_hi_hi = _GEN_50;
  wire [127:0]       regroupV0_lo_hi_hi_lo_lo_hi = {regroupV0_lo_hi_hi_lo_lo_hi_hi, regroupV0_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]       regroupV0_lo_hi_hi_lo_lo = {regroupV0_lo_hi_hi_lo_lo_hi, regroupV0_lo_hi_hi_lo_lo_lo};
  wire [63:0]        _GEN_51 = {v0_105, v0_104};
  wire [63:0]        regroupV0_lo_hi_hi_lo_hi_lo_lo;
  assign regroupV0_lo_hi_hi_lo_hi_lo_lo = _GEN_51;
  wire [63:0]        regroupV0_lo_hi_hi_lo_hi_lo_lo_5;
  assign regroupV0_lo_hi_hi_lo_hi_lo_lo_5 = _GEN_51;
  wire [63:0]        regroupV0_lo_hi_hi_lo_hi_lo_lo_10;
  assign regroupV0_lo_hi_hi_lo_hi_lo_lo_10 = _GEN_51;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_hi_lo_hi_lo_lo;
  assign slideAddressGen_slideMaskInput_lo_hi_hi_lo_hi_lo_lo = _GEN_51;
  wire [63:0]        selectReadStageMask_lo_hi_hi_lo_hi_lo_lo;
  assign selectReadStageMask_lo_hi_hi_lo_hi_lo_lo = _GEN_51;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_hi_lo_lo;
  assign maskSplit_maskSelect_lo_hi_hi_lo_hi_lo_lo = _GEN_51;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_hi_lo_lo_1;
  assign maskSplit_maskSelect_lo_hi_hi_lo_hi_lo_lo_1 = _GEN_51;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_hi_lo_lo_2;
  assign maskSplit_maskSelect_lo_hi_hi_lo_hi_lo_lo_2 = _GEN_51;
  wire [63:0]        maskForDestination_lo_hi_hi_lo_hi_lo_lo;
  assign maskForDestination_lo_hi_hi_lo_hi_lo_lo = _GEN_51;
  wire [63:0]        _GEN_52 = {v0_107, v0_106};
  wire [63:0]        regroupV0_lo_hi_hi_lo_hi_lo_hi;
  assign regroupV0_lo_hi_hi_lo_hi_lo_hi = _GEN_52;
  wire [63:0]        regroupV0_lo_hi_hi_lo_hi_lo_hi_5;
  assign regroupV0_lo_hi_hi_lo_hi_lo_hi_5 = _GEN_52;
  wire [63:0]        regroupV0_lo_hi_hi_lo_hi_lo_hi_10;
  assign regroupV0_lo_hi_hi_lo_hi_lo_hi_10 = _GEN_52;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_hi_lo_hi_lo_hi;
  assign slideAddressGen_slideMaskInput_lo_hi_hi_lo_hi_lo_hi = _GEN_52;
  wire [63:0]        selectReadStageMask_lo_hi_hi_lo_hi_lo_hi;
  assign selectReadStageMask_lo_hi_hi_lo_hi_lo_hi = _GEN_52;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_hi_lo_hi;
  assign maskSplit_maskSelect_lo_hi_hi_lo_hi_lo_hi = _GEN_52;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_hi_lo_hi_1;
  assign maskSplit_maskSelect_lo_hi_hi_lo_hi_lo_hi_1 = _GEN_52;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_hi_lo_hi_2;
  assign maskSplit_maskSelect_lo_hi_hi_lo_hi_lo_hi_2 = _GEN_52;
  wire [63:0]        maskForDestination_lo_hi_hi_lo_hi_lo_hi;
  assign maskForDestination_lo_hi_hi_lo_hi_lo_hi = _GEN_52;
  wire [127:0]       regroupV0_lo_hi_hi_lo_hi_lo = {regroupV0_lo_hi_hi_lo_hi_lo_hi, regroupV0_lo_hi_hi_lo_hi_lo_lo};
  wire [63:0]        _GEN_53 = {v0_109, v0_108};
  wire [63:0]        regroupV0_lo_hi_hi_lo_hi_hi_lo;
  assign regroupV0_lo_hi_hi_lo_hi_hi_lo = _GEN_53;
  wire [63:0]        regroupV0_lo_hi_hi_lo_hi_hi_lo_5;
  assign regroupV0_lo_hi_hi_lo_hi_hi_lo_5 = _GEN_53;
  wire [63:0]        regroupV0_lo_hi_hi_lo_hi_hi_lo_10;
  assign regroupV0_lo_hi_hi_lo_hi_hi_lo_10 = _GEN_53;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_hi_lo_hi_hi_lo;
  assign slideAddressGen_slideMaskInput_lo_hi_hi_lo_hi_hi_lo = _GEN_53;
  wire [63:0]        selectReadStageMask_lo_hi_hi_lo_hi_hi_lo;
  assign selectReadStageMask_lo_hi_hi_lo_hi_hi_lo = _GEN_53;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_hi_hi_lo;
  assign maskSplit_maskSelect_lo_hi_hi_lo_hi_hi_lo = _GEN_53;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_hi_hi_lo_1;
  assign maskSplit_maskSelect_lo_hi_hi_lo_hi_hi_lo_1 = _GEN_53;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_hi_hi_lo_2;
  assign maskSplit_maskSelect_lo_hi_hi_lo_hi_hi_lo_2 = _GEN_53;
  wire [63:0]        maskForDestination_lo_hi_hi_lo_hi_hi_lo;
  assign maskForDestination_lo_hi_hi_lo_hi_hi_lo = _GEN_53;
  wire [63:0]        _GEN_54 = {v0_111, v0_110};
  wire [63:0]        regroupV0_lo_hi_hi_lo_hi_hi_hi;
  assign regroupV0_lo_hi_hi_lo_hi_hi_hi = _GEN_54;
  wire [63:0]        regroupV0_lo_hi_hi_lo_hi_hi_hi_5;
  assign regroupV0_lo_hi_hi_lo_hi_hi_hi_5 = _GEN_54;
  wire [63:0]        regroupV0_lo_hi_hi_lo_hi_hi_hi_10;
  assign regroupV0_lo_hi_hi_lo_hi_hi_hi_10 = _GEN_54;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_hi_lo_hi_hi_hi;
  assign slideAddressGen_slideMaskInput_lo_hi_hi_lo_hi_hi_hi = _GEN_54;
  wire [63:0]        selectReadStageMask_lo_hi_hi_lo_hi_hi_hi;
  assign selectReadStageMask_lo_hi_hi_lo_hi_hi_hi = _GEN_54;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_hi_hi_hi;
  assign maskSplit_maskSelect_lo_hi_hi_lo_hi_hi_hi = _GEN_54;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_hi_hi_hi_1;
  assign maskSplit_maskSelect_lo_hi_hi_lo_hi_hi_hi_1 = _GEN_54;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_hi_hi_hi_2;
  assign maskSplit_maskSelect_lo_hi_hi_lo_hi_hi_hi_2 = _GEN_54;
  wire [63:0]        maskForDestination_lo_hi_hi_lo_hi_hi_hi;
  assign maskForDestination_lo_hi_hi_lo_hi_hi_hi = _GEN_54;
  wire [127:0]       regroupV0_lo_hi_hi_lo_hi_hi = {regroupV0_lo_hi_hi_lo_hi_hi_hi, regroupV0_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]       regroupV0_lo_hi_hi_lo_hi = {regroupV0_lo_hi_hi_lo_hi_hi, regroupV0_lo_hi_hi_lo_hi_lo};
  wire [511:0]       regroupV0_lo_hi_hi_lo = {regroupV0_lo_hi_hi_lo_hi, regroupV0_lo_hi_hi_lo_lo};
  wire [63:0]        _GEN_55 = {v0_113, v0_112};
  wire [63:0]        regroupV0_lo_hi_hi_hi_lo_lo_lo;
  assign regroupV0_lo_hi_hi_hi_lo_lo_lo = _GEN_55;
  wire [63:0]        regroupV0_lo_hi_hi_hi_lo_lo_lo_5;
  assign regroupV0_lo_hi_hi_hi_lo_lo_lo_5 = _GEN_55;
  wire [63:0]        regroupV0_lo_hi_hi_hi_lo_lo_lo_10;
  assign regroupV0_lo_hi_hi_hi_lo_lo_lo_10 = _GEN_55;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_hi_hi_lo_lo_lo;
  assign slideAddressGen_slideMaskInput_lo_hi_hi_hi_lo_lo_lo = _GEN_55;
  wire [63:0]        selectReadStageMask_lo_hi_hi_hi_lo_lo_lo;
  assign selectReadStageMask_lo_hi_hi_hi_lo_lo_lo = _GEN_55;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_lo_lo_lo;
  assign maskSplit_maskSelect_lo_hi_hi_hi_lo_lo_lo = _GEN_55;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_lo_lo_lo_1;
  assign maskSplit_maskSelect_lo_hi_hi_hi_lo_lo_lo_1 = _GEN_55;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_lo_lo_lo_2;
  assign maskSplit_maskSelect_lo_hi_hi_hi_lo_lo_lo_2 = _GEN_55;
  wire [63:0]        maskForDestination_lo_hi_hi_hi_lo_lo_lo;
  assign maskForDestination_lo_hi_hi_hi_lo_lo_lo = _GEN_55;
  wire [63:0]        _GEN_56 = {v0_115, v0_114};
  wire [63:0]        regroupV0_lo_hi_hi_hi_lo_lo_hi;
  assign regroupV0_lo_hi_hi_hi_lo_lo_hi = _GEN_56;
  wire [63:0]        regroupV0_lo_hi_hi_hi_lo_lo_hi_5;
  assign regroupV0_lo_hi_hi_hi_lo_lo_hi_5 = _GEN_56;
  wire [63:0]        regroupV0_lo_hi_hi_hi_lo_lo_hi_10;
  assign regroupV0_lo_hi_hi_hi_lo_lo_hi_10 = _GEN_56;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_hi_hi_lo_lo_hi;
  assign slideAddressGen_slideMaskInput_lo_hi_hi_hi_lo_lo_hi = _GEN_56;
  wire [63:0]        selectReadStageMask_lo_hi_hi_hi_lo_lo_hi;
  assign selectReadStageMask_lo_hi_hi_hi_lo_lo_hi = _GEN_56;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_lo_lo_hi;
  assign maskSplit_maskSelect_lo_hi_hi_hi_lo_lo_hi = _GEN_56;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_lo_lo_hi_1;
  assign maskSplit_maskSelect_lo_hi_hi_hi_lo_lo_hi_1 = _GEN_56;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_lo_lo_hi_2;
  assign maskSplit_maskSelect_lo_hi_hi_hi_lo_lo_hi_2 = _GEN_56;
  wire [63:0]        maskForDestination_lo_hi_hi_hi_lo_lo_hi;
  assign maskForDestination_lo_hi_hi_hi_lo_lo_hi = _GEN_56;
  wire [127:0]       regroupV0_lo_hi_hi_hi_lo_lo = {regroupV0_lo_hi_hi_hi_lo_lo_hi, regroupV0_lo_hi_hi_hi_lo_lo_lo};
  wire [63:0]        _GEN_57 = {v0_117, v0_116};
  wire [63:0]        regroupV0_lo_hi_hi_hi_lo_hi_lo;
  assign regroupV0_lo_hi_hi_hi_lo_hi_lo = _GEN_57;
  wire [63:0]        regroupV0_lo_hi_hi_hi_lo_hi_lo_5;
  assign regroupV0_lo_hi_hi_hi_lo_hi_lo_5 = _GEN_57;
  wire [63:0]        regroupV0_lo_hi_hi_hi_lo_hi_lo_10;
  assign regroupV0_lo_hi_hi_hi_lo_hi_lo_10 = _GEN_57;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_hi_hi_lo_hi_lo;
  assign slideAddressGen_slideMaskInput_lo_hi_hi_hi_lo_hi_lo = _GEN_57;
  wire [63:0]        selectReadStageMask_lo_hi_hi_hi_lo_hi_lo;
  assign selectReadStageMask_lo_hi_hi_hi_lo_hi_lo = _GEN_57;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_lo_hi_lo;
  assign maskSplit_maskSelect_lo_hi_hi_hi_lo_hi_lo = _GEN_57;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_lo_hi_lo_1;
  assign maskSplit_maskSelect_lo_hi_hi_hi_lo_hi_lo_1 = _GEN_57;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_lo_hi_lo_2;
  assign maskSplit_maskSelect_lo_hi_hi_hi_lo_hi_lo_2 = _GEN_57;
  wire [63:0]        maskForDestination_lo_hi_hi_hi_lo_hi_lo;
  assign maskForDestination_lo_hi_hi_hi_lo_hi_lo = _GEN_57;
  wire [63:0]        _GEN_58 = {v0_119, v0_118};
  wire [63:0]        regroupV0_lo_hi_hi_hi_lo_hi_hi;
  assign regroupV0_lo_hi_hi_hi_lo_hi_hi = _GEN_58;
  wire [63:0]        regroupV0_lo_hi_hi_hi_lo_hi_hi_5;
  assign regroupV0_lo_hi_hi_hi_lo_hi_hi_5 = _GEN_58;
  wire [63:0]        regroupV0_lo_hi_hi_hi_lo_hi_hi_10;
  assign regroupV0_lo_hi_hi_hi_lo_hi_hi_10 = _GEN_58;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_hi_hi_lo_hi_hi;
  assign slideAddressGen_slideMaskInput_lo_hi_hi_hi_lo_hi_hi = _GEN_58;
  wire [63:0]        selectReadStageMask_lo_hi_hi_hi_lo_hi_hi;
  assign selectReadStageMask_lo_hi_hi_hi_lo_hi_hi = _GEN_58;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_lo_hi_hi;
  assign maskSplit_maskSelect_lo_hi_hi_hi_lo_hi_hi = _GEN_58;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_lo_hi_hi_1;
  assign maskSplit_maskSelect_lo_hi_hi_hi_lo_hi_hi_1 = _GEN_58;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_lo_hi_hi_2;
  assign maskSplit_maskSelect_lo_hi_hi_hi_lo_hi_hi_2 = _GEN_58;
  wire [63:0]        maskForDestination_lo_hi_hi_hi_lo_hi_hi;
  assign maskForDestination_lo_hi_hi_hi_lo_hi_hi = _GEN_58;
  wire [127:0]       regroupV0_lo_hi_hi_hi_lo_hi = {regroupV0_lo_hi_hi_hi_lo_hi_hi, regroupV0_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]       regroupV0_lo_hi_hi_hi_lo = {regroupV0_lo_hi_hi_hi_lo_hi, regroupV0_lo_hi_hi_hi_lo_lo};
  wire [63:0]        _GEN_59 = {v0_121, v0_120};
  wire [63:0]        regroupV0_lo_hi_hi_hi_hi_lo_lo;
  assign regroupV0_lo_hi_hi_hi_hi_lo_lo = _GEN_59;
  wire [63:0]        regroupV0_lo_hi_hi_hi_hi_lo_lo_5;
  assign regroupV0_lo_hi_hi_hi_hi_lo_lo_5 = _GEN_59;
  wire [63:0]        regroupV0_lo_hi_hi_hi_hi_lo_lo_10;
  assign regroupV0_lo_hi_hi_hi_hi_lo_lo_10 = _GEN_59;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_hi_hi_hi_lo_lo;
  assign slideAddressGen_slideMaskInput_lo_hi_hi_hi_hi_lo_lo = _GEN_59;
  wire [63:0]        selectReadStageMask_lo_hi_hi_hi_hi_lo_lo;
  assign selectReadStageMask_lo_hi_hi_hi_hi_lo_lo = _GEN_59;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_hi_lo_lo;
  assign maskSplit_maskSelect_lo_hi_hi_hi_hi_lo_lo = _GEN_59;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_hi_lo_lo_1;
  assign maskSplit_maskSelect_lo_hi_hi_hi_hi_lo_lo_1 = _GEN_59;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_hi_lo_lo_2;
  assign maskSplit_maskSelect_lo_hi_hi_hi_hi_lo_lo_2 = _GEN_59;
  wire [63:0]        maskForDestination_lo_hi_hi_hi_hi_lo_lo;
  assign maskForDestination_lo_hi_hi_hi_hi_lo_lo = _GEN_59;
  wire [63:0]        _GEN_60 = {v0_123, v0_122};
  wire [63:0]        regroupV0_lo_hi_hi_hi_hi_lo_hi;
  assign regroupV0_lo_hi_hi_hi_hi_lo_hi = _GEN_60;
  wire [63:0]        regroupV0_lo_hi_hi_hi_hi_lo_hi_5;
  assign regroupV0_lo_hi_hi_hi_hi_lo_hi_5 = _GEN_60;
  wire [63:0]        regroupV0_lo_hi_hi_hi_hi_lo_hi_10;
  assign regroupV0_lo_hi_hi_hi_hi_lo_hi_10 = _GEN_60;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_hi_hi_hi_lo_hi;
  assign slideAddressGen_slideMaskInput_lo_hi_hi_hi_hi_lo_hi = _GEN_60;
  wire [63:0]        selectReadStageMask_lo_hi_hi_hi_hi_lo_hi;
  assign selectReadStageMask_lo_hi_hi_hi_hi_lo_hi = _GEN_60;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_hi_lo_hi;
  assign maskSplit_maskSelect_lo_hi_hi_hi_hi_lo_hi = _GEN_60;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_hi_lo_hi_1;
  assign maskSplit_maskSelect_lo_hi_hi_hi_hi_lo_hi_1 = _GEN_60;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_hi_lo_hi_2;
  assign maskSplit_maskSelect_lo_hi_hi_hi_hi_lo_hi_2 = _GEN_60;
  wire [63:0]        maskForDestination_lo_hi_hi_hi_hi_lo_hi;
  assign maskForDestination_lo_hi_hi_hi_hi_lo_hi = _GEN_60;
  wire [127:0]       regroupV0_lo_hi_hi_hi_hi_lo = {regroupV0_lo_hi_hi_hi_hi_lo_hi, regroupV0_lo_hi_hi_hi_hi_lo_lo};
  wire [63:0]        _GEN_61 = {v0_125, v0_124};
  wire [63:0]        regroupV0_lo_hi_hi_hi_hi_hi_lo;
  assign regroupV0_lo_hi_hi_hi_hi_hi_lo = _GEN_61;
  wire [63:0]        regroupV0_lo_hi_hi_hi_hi_hi_lo_5;
  assign regroupV0_lo_hi_hi_hi_hi_hi_lo_5 = _GEN_61;
  wire [63:0]        regroupV0_lo_hi_hi_hi_hi_hi_lo_10;
  assign regroupV0_lo_hi_hi_hi_hi_hi_lo_10 = _GEN_61;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_hi_hi_hi_hi_lo;
  assign slideAddressGen_slideMaskInput_lo_hi_hi_hi_hi_hi_lo = _GEN_61;
  wire [63:0]        selectReadStageMask_lo_hi_hi_hi_hi_hi_lo;
  assign selectReadStageMask_lo_hi_hi_hi_hi_hi_lo = _GEN_61;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_hi_hi_lo;
  assign maskSplit_maskSelect_lo_hi_hi_hi_hi_hi_lo = _GEN_61;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_hi_hi_lo_1;
  assign maskSplit_maskSelect_lo_hi_hi_hi_hi_hi_lo_1 = _GEN_61;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_hi_hi_lo_2;
  assign maskSplit_maskSelect_lo_hi_hi_hi_hi_hi_lo_2 = _GEN_61;
  wire [63:0]        maskForDestination_lo_hi_hi_hi_hi_hi_lo;
  assign maskForDestination_lo_hi_hi_hi_hi_hi_lo = _GEN_61;
  wire [63:0]        _GEN_62 = {v0_127, v0_126};
  wire [63:0]        regroupV0_lo_hi_hi_hi_hi_hi_hi;
  assign regroupV0_lo_hi_hi_hi_hi_hi_hi = _GEN_62;
  wire [63:0]        regroupV0_lo_hi_hi_hi_hi_hi_hi_5;
  assign regroupV0_lo_hi_hi_hi_hi_hi_hi_5 = _GEN_62;
  wire [63:0]        regroupV0_lo_hi_hi_hi_hi_hi_hi_10;
  assign regroupV0_lo_hi_hi_hi_hi_hi_hi_10 = _GEN_62;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_hi_hi_hi_hi_hi;
  assign slideAddressGen_slideMaskInput_lo_hi_hi_hi_hi_hi_hi = _GEN_62;
  wire [63:0]        selectReadStageMask_lo_hi_hi_hi_hi_hi_hi;
  assign selectReadStageMask_lo_hi_hi_hi_hi_hi_hi = _GEN_62;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_hi_hi_hi;
  assign maskSplit_maskSelect_lo_hi_hi_hi_hi_hi_hi = _GEN_62;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_hi_hi_hi_1;
  assign maskSplit_maskSelect_lo_hi_hi_hi_hi_hi_hi_1 = _GEN_62;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_hi_hi_hi_2;
  assign maskSplit_maskSelect_lo_hi_hi_hi_hi_hi_hi_2 = _GEN_62;
  wire [63:0]        maskForDestination_lo_hi_hi_hi_hi_hi_hi;
  assign maskForDestination_lo_hi_hi_hi_hi_hi_hi = _GEN_62;
  wire [127:0]       regroupV0_lo_hi_hi_hi_hi_hi = {regroupV0_lo_hi_hi_hi_hi_hi_hi, regroupV0_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]       regroupV0_lo_hi_hi_hi_hi = {regroupV0_lo_hi_hi_hi_hi_hi, regroupV0_lo_hi_hi_hi_hi_lo};
  wire [511:0]       regroupV0_lo_hi_hi_hi = {regroupV0_lo_hi_hi_hi_hi, regroupV0_lo_hi_hi_hi_lo};
  wire [1023:0]      regroupV0_lo_hi_hi = {regroupV0_lo_hi_hi_hi, regroupV0_lo_hi_hi_lo};
  wire [2047:0]      regroupV0_lo_hi = {regroupV0_lo_hi_hi, regroupV0_lo_hi_lo};
  wire [4095:0]      regroupV0_lo = {regroupV0_lo_hi, regroupV0_lo_lo};
  wire [63:0]        _GEN_63 = {v0_129, v0_128};
  wire [63:0]        regroupV0_hi_lo_lo_lo_lo_lo_lo;
  assign regroupV0_hi_lo_lo_lo_lo_lo_lo = _GEN_63;
  wire [63:0]        regroupV0_hi_lo_lo_lo_lo_lo_lo_5;
  assign regroupV0_hi_lo_lo_lo_lo_lo_lo_5 = _GEN_63;
  wire [63:0]        regroupV0_hi_lo_lo_lo_lo_lo_lo_10;
  assign regroupV0_hi_lo_lo_lo_lo_lo_lo_10 = _GEN_63;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_lo_lo_lo_lo_lo;
  assign slideAddressGen_slideMaskInput_hi_lo_lo_lo_lo_lo_lo = _GEN_63;
  wire [63:0]        selectReadStageMask_hi_lo_lo_lo_lo_lo_lo;
  assign selectReadStageMask_hi_lo_lo_lo_lo_lo_lo = _GEN_63;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_lo_lo_lo;
  assign maskSplit_maskSelect_hi_lo_lo_lo_lo_lo_lo = _GEN_63;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_lo_lo_lo_1;
  assign maskSplit_maskSelect_hi_lo_lo_lo_lo_lo_lo_1 = _GEN_63;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_lo_lo_lo_2;
  assign maskSplit_maskSelect_hi_lo_lo_lo_lo_lo_lo_2 = _GEN_63;
  wire [63:0]        maskForDestination_hi_lo_lo_lo_lo_lo_lo;
  assign maskForDestination_hi_lo_lo_lo_lo_lo_lo = _GEN_63;
  wire [63:0]        _GEN_64 = {v0_131, v0_130};
  wire [63:0]        regroupV0_hi_lo_lo_lo_lo_lo_hi;
  assign regroupV0_hi_lo_lo_lo_lo_lo_hi = _GEN_64;
  wire [63:0]        regroupV0_hi_lo_lo_lo_lo_lo_hi_5;
  assign regroupV0_hi_lo_lo_lo_lo_lo_hi_5 = _GEN_64;
  wire [63:0]        regroupV0_hi_lo_lo_lo_lo_lo_hi_10;
  assign regroupV0_hi_lo_lo_lo_lo_lo_hi_10 = _GEN_64;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_lo_lo_lo_lo_hi;
  assign slideAddressGen_slideMaskInput_hi_lo_lo_lo_lo_lo_hi = _GEN_64;
  wire [63:0]        selectReadStageMask_hi_lo_lo_lo_lo_lo_hi;
  assign selectReadStageMask_hi_lo_lo_lo_lo_lo_hi = _GEN_64;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_lo_lo_hi;
  assign maskSplit_maskSelect_hi_lo_lo_lo_lo_lo_hi = _GEN_64;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_lo_lo_hi_1;
  assign maskSplit_maskSelect_hi_lo_lo_lo_lo_lo_hi_1 = _GEN_64;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_lo_lo_hi_2;
  assign maskSplit_maskSelect_hi_lo_lo_lo_lo_lo_hi_2 = _GEN_64;
  wire [63:0]        maskForDestination_hi_lo_lo_lo_lo_lo_hi;
  assign maskForDestination_hi_lo_lo_lo_lo_lo_hi = _GEN_64;
  wire [127:0]       regroupV0_hi_lo_lo_lo_lo_lo = {regroupV0_hi_lo_lo_lo_lo_lo_hi, regroupV0_hi_lo_lo_lo_lo_lo_lo};
  wire [63:0]        _GEN_65 = {v0_133, v0_132};
  wire [63:0]        regroupV0_hi_lo_lo_lo_lo_hi_lo;
  assign regroupV0_hi_lo_lo_lo_lo_hi_lo = _GEN_65;
  wire [63:0]        regroupV0_hi_lo_lo_lo_lo_hi_lo_5;
  assign regroupV0_hi_lo_lo_lo_lo_hi_lo_5 = _GEN_65;
  wire [63:0]        regroupV0_hi_lo_lo_lo_lo_hi_lo_10;
  assign regroupV0_hi_lo_lo_lo_lo_hi_lo_10 = _GEN_65;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_lo_lo_lo_hi_lo;
  assign slideAddressGen_slideMaskInput_hi_lo_lo_lo_lo_hi_lo = _GEN_65;
  wire [63:0]        selectReadStageMask_hi_lo_lo_lo_lo_hi_lo;
  assign selectReadStageMask_hi_lo_lo_lo_lo_hi_lo = _GEN_65;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_lo_hi_lo;
  assign maskSplit_maskSelect_hi_lo_lo_lo_lo_hi_lo = _GEN_65;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_lo_hi_lo_1;
  assign maskSplit_maskSelect_hi_lo_lo_lo_lo_hi_lo_1 = _GEN_65;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_lo_hi_lo_2;
  assign maskSplit_maskSelect_hi_lo_lo_lo_lo_hi_lo_2 = _GEN_65;
  wire [63:0]        maskForDestination_hi_lo_lo_lo_lo_hi_lo;
  assign maskForDestination_hi_lo_lo_lo_lo_hi_lo = _GEN_65;
  wire [63:0]        _GEN_66 = {v0_135, v0_134};
  wire [63:0]        regroupV0_hi_lo_lo_lo_lo_hi_hi;
  assign regroupV0_hi_lo_lo_lo_lo_hi_hi = _GEN_66;
  wire [63:0]        regroupV0_hi_lo_lo_lo_lo_hi_hi_5;
  assign regroupV0_hi_lo_lo_lo_lo_hi_hi_5 = _GEN_66;
  wire [63:0]        regroupV0_hi_lo_lo_lo_lo_hi_hi_10;
  assign regroupV0_hi_lo_lo_lo_lo_hi_hi_10 = _GEN_66;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_lo_lo_lo_hi_hi;
  assign slideAddressGen_slideMaskInput_hi_lo_lo_lo_lo_hi_hi = _GEN_66;
  wire [63:0]        selectReadStageMask_hi_lo_lo_lo_lo_hi_hi;
  assign selectReadStageMask_hi_lo_lo_lo_lo_hi_hi = _GEN_66;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_lo_hi_hi;
  assign maskSplit_maskSelect_hi_lo_lo_lo_lo_hi_hi = _GEN_66;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_lo_hi_hi_1;
  assign maskSplit_maskSelect_hi_lo_lo_lo_lo_hi_hi_1 = _GEN_66;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_lo_hi_hi_2;
  assign maskSplit_maskSelect_hi_lo_lo_lo_lo_hi_hi_2 = _GEN_66;
  wire [63:0]        maskForDestination_hi_lo_lo_lo_lo_hi_hi;
  assign maskForDestination_hi_lo_lo_lo_lo_hi_hi = _GEN_66;
  wire [127:0]       regroupV0_hi_lo_lo_lo_lo_hi = {regroupV0_hi_lo_lo_lo_lo_hi_hi, regroupV0_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]       regroupV0_hi_lo_lo_lo_lo = {regroupV0_hi_lo_lo_lo_lo_hi, regroupV0_hi_lo_lo_lo_lo_lo};
  wire [63:0]        _GEN_67 = {v0_137, v0_136};
  wire [63:0]        regroupV0_hi_lo_lo_lo_hi_lo_lo;
  assign regroupV0_hi_lo_lo_lo_hi_lo_lo = _GEN_67;
  wire [63:0]        regroupV0_hi_lo_lo_lo_hi_lo_lo_5;
  assign regroupV0_hi_lo_lo_lo_hi_lo_lo_5 = _GEN_67;
  wire [63:0]        regroupV0_hi_lo_lo_lo_hi_lo_lo_10;
  assign regroupV0_hi_lo_lo_lo_hi_lo_lo_10 = _GEN_67;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_lo_lo_hi_lo_lo;
  assign slideAddressGen_slideMaskInput_hi_lo_lo_lo_hi_lo_lo = _GEN_67;
  wire [63:0]        selectReadStageMask_hi_lo_lo_lo_hi_lo_lo;
  assign selectReadStageMask_hi_lo_lo_lo_hi_lo_lo = _GEN_67;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_hi_lo_lo;
  assign maskSplit_maskSelect_hi_lo_lo_lo_hi_lo_lo = _GEN_67;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_hi_lo_lo_1;
  assign maskSplit_maskSelect_hi_lo_lo_lo_hi_lo_lo_1 = _GEN_67;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_hi_lo_lo_2;
  assign maskSplit_maskSelect_hi_lo_lo_lo_hi_lo_lo_2 = _GEN_67;
  wire [63:0]        maskForDestination_hi_lo_lo_lo_hi_lo_lo;
  assign maskForDestination_hi_lo_lo_lo_hi_lo_lo = _GEN_67;
  wire [63:0]        _GEN_68 = {v0_139, v0_138};
  wire [63:0]        regroupV0_hi_lo_lo_lo_hi_lo_hi;
  assign regroupV0_hi_lo_lo_lo_hi_lo_hi = _GEN_68;
  wire [63:0]        regroupV0_hi_lo_lo_lo_hi_lo_hi_5;
  assign regroupV0_hi_lo_lo_lo_hi_lo_hi_5 = _GEN_68;
  wire [63:0]        regroupV0_hi_lo_lo_lo_hi_lo_hi_10;
  assign regroupV0_hi_lo_lo_lo_hi_lo_hi_10 = _GEN_68;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_lo_lo_hi_lo_hi;
  assign slideAddressGen_slideMaskInput_hi_lo_lo_lo_hi_lo_hi = _GEN_68;
  wire [63:0]        selectReadStageMask_hi_lo_lo_lo_hi_lo_hi;
  assign selectReadStageMask_hi_lo_lo_lo_hi_lo_hi = _GEN_68;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_hi_lo_hi;
  assign maskSplit_maskSelect_hi_lo_lo_lo_hi_lo_hi = _GEN_68;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_hi_lo_hi_1;
  assign maskSplit_maskSelect_hi_lo_lo_lo_hi_lo_hi_1 = _GEN_68;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_hi_lo_hi_2;
  assign maskSplit_maskSelect_hi_lo_lo_lo_hi_lo_hi_2 = _GEN_68;
  wire [63:0]        maskForDestination_hi_lo_lo_lo_hi_lo_hi;
  assign maskForDestination_hi_lo_lo_lo_hi_lo_hi = _GEN_68;
  wire [127:0]       regroupV0_hi_lo_lo_lo_hi_lo = {regroupV0_hi_lo_lo_lo_hi_lo_hi, regroupV0_hi_lo_lo_lo_hi_lo_lo};
  wire [63:0]        _GEN_69 = {v0_141, v0_140};
  wire [63:0]        regroupV0_hi_lo_lo_lo_hi_hi_lo;
  assign regroupV0_hi_lo_lo_lo_hi_hi_lo = _GEN_69;
  wire [63:0]        regroupV0_hi_lo_lo_lo_hi_hi_lo_5;
  assign regroupV0_hi_lo_lo_lo_hi_hi_lo_5 = _GEN_69;
  wire [63:0]        regroupV0_hi_lo_lo_lo_hi_hi_lo_10;
  assign regroupV0_hi_lo_lo_lo_hi_hi_lo_10 = _GEN_69;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_lo_lo_hi_hi_lo;
  assign slideAddressGen_slideMaskInput_hi_lo_lo_lo_hi_hi_lo = _GEN_69;
  wire [63:0]        selectReadStageMask_hi_lo_lo_lo_hi_hi_lo;
  assign selectReadStageMask_hi_lo_lo_lo_hi_hi_lo = _GEN_69;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_hi_hi_lo;
  assign maskSplit_maskSelect_hi_lo_lo_lo_hi_hi_lo = _GEN_69;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_hi_hi_lo_1;
  assign maskSplit_maskSelect_hi_lo_lo_lo_hi_hi_lo_1 = _GEN_69;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_hi_hi_lo_2;
  assign maskSplit_maskSelect_hi_lo_lo_lo_hi_hi_lo_2 = _GEN_69;
  wire [63:0]        maskForDestination_hi_lo_lo_lo_hi_hi_lo;
  assign maskForDestination_hi_lo_lo_lo_hi_hi_lo = _GEN_69;
  wire [63:0]        _GEN_70 = {v0_143, v0_142};
  wire [63:0]        regroupV0_hi_lo_lo_lo_hi_hi_hi;
  assign regroupV0_hi_lo_lo_lo_hi_hi_hi = _GEN_70;
  wire [63:0]        regroupV0_hi_lo_lo_lo_hi_hi_hi_5;
  assign regroupV0_hi_lo_lo_lo_hi_hi_hi_5 = _GEN_70;
  wire [63:0]        regroupV0_hi_lo_lo_lo_hi_hi_hi_10;
  assign regroupV0_hi_lo_lo_lo_hi_hi_hi_10 = _GEN_70;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_lo_lo_hi_hi_hi;
  assign slideAddressGen_slideMaskInput_hi_lo_lo_lo_hi_hi_hi = _GEN_70;
  wire [63:0]        selectReadStageMask_hi_lo_lo_lo_hi_hi_hi;
  assign selectReadStageMask_hi_lo_lo_lo_hi_hi_hi = _GEN_70;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_hi_hi_hi;
  assign maskSplit_maskSelect_hi_lo_lo_lo_hi_hi_hi = _GEN_70;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_hi_hi_hi_1;
  assign maskSplit_maskSelect_hi_lo_lo_lo_hi_hi_hi_1 = _GEN_70;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_hi_hi_hi_2;
  assign maskSplit_maskSelect_hi_lo_lo_lo_hi_hi_hi_2 = _GEN_70;
  wire [63:0]        maskForDestination_hi_lo_lo_lo_hi_hi_hi;
  assign maskForDestination_hi_lo_lo_lo_hi_hi_hi = _GEN_70;
  wire [127:0]       regroupV0_hi_lo_lo_lo_hi_hi = {regroupV0_hi_lo_lo_lo_hi_hi_hi, regroupV0_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]       regroupV0_hi_lo_lo_lo_hi = {regroupV0_hi_lo_lo_lo_hi_hi, regroupV0_hi_lo_lo_lo_hi_lo};
  wire [511:0]       regroupV0_hi_lo_lo_lo = {regroupV0_hi_lo_lo_lo_hi, regroupV0_hi_lo_lo_lo_lo};
  wire [63:0]        _GEN_71 = {v0_145, v0_144};
  wire [63:0]        regroupV0_hi_lo_lo_hi_lo_lo_lo;
  assign regroupV0_hi_lo_lo_hi_lo_lo_lo = _GEN_71;
  wire [63:0]        regroupV0_hi_lo_lo_hi_lo_lo_lo_5;
  assign regroupV0_hi_lo_lo_hi_lo_lo_lo_5 = _GEN_71;
  wire [63:0]        regroupV0_hi_lo_lo_hi_lo_lo_lo_10;
  assign regroupV0_hi_lo_lo_hi_lo_lo_lo_10 = _GEN_71;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_lo_hi_lo_lo_lo;
  assign slideAddressGen_slideMaskInput_hi_lo_lo_hi_lo_lo_lo = _GEN_71;
  wire [63:0]        selectReadStageMask_hi_lo_lo_hi_lo_lo_lo;
  assign selectReadStageMask_hi_lo_lo_hi_lo_lo_lo = _GEN_71;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_lo_lo_lo;
  assign maskSplit_maskSelect_hi_lo_lo_hi_lo_lo_lo = _GEN_71;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_lo_lo_lo_1;
  assign maskSplit_maskSelect_hi_lo_lo_hi_lo_lo_lo_1 = _GEN_71;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_lo_lo_lo_2;
  assign maskSplit_maskSelect_hi_lo_lo_hi_lo_lo_lo_2 = _GEN_71;
  wire [63:0]        maskForDestination_hi_lo_lo_hi_lo_lo_lo;
  assign maskForDestination_hi_lo_lo_hi_lo_lo_lo = _GEN_71;
  wire [63:0]        _GEN_72 = {v0_147, v0_146};
  wire [63:0]        regroupV0_hi_lo_lo_hi_lo_lo_hi;
  assign regroupV0_hi_lo_lo_hi_lo_lo_hi = _GEN_72;
  wire [63:0]        regroupV0_hi_lo_lo_hi_lo_lo_hi_5;
  assign regroupV0_hi_lo_lo_hi_lo_lo_hi_5 = _GEN_72;
  wire [63:0]        regroupV0_hi_lo_lo_hi_lo_lo_hi_10;
  assign regroupV0_hi_lo_lo_hi_lo_lo_hi_10 = _GEN_72;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_lo_hi_lo_lo_hi;
  assign slideAddressGen_slideMaskInput_hi_lo_lo_hi_lo_lo_hi = _GEN_72;
  wire [63:0]        selectReadStageMask_hi_lo_lo_hi_lo_lo_hi;
  assign selectReadStageMask_hi_lo_lo_hi_lo_lo_hi = _GEN_72;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_lo_lo_hi;
  assign maskSplit_maskSelect_hi_lo_lo_hi_lo_lo_hi = _GEN_72;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_lo_lo_hi_1;
  assign maskSplit_maskSelect_hi_lo_lo_hi_lo_lo_hi_1 = _GEN_72;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_lo_lo_hi_2;
  assign maskSplit_maskSelect_hi_lo_lo_hi_lo_lo_hi_2 = _GEN_72;
  wire [63:0]        maskForDestination_hi_lo_lo_hi_lo_lo_hi;
  assign maskForDestination_hi_lo_lo_hi_lo_lo_hi = _GEN_72;
  wire [127:0]       regroupV0_hi_lo_lo_hi_lo_lo = {regroupV0_hi_lo_lo_hi_lo_lo_hi, regroupV0_hi_lo_lo_hi_lo_lo_lo};
  wire [63:0]        _GEN_73 = {v0_149, v0_148};
  wire [63:0]        regroupV0_hi_lo_lo_hi_lo_hi_lo;
  assign regroupV0_hi_lo_lo_hi_lo_hi_lo = _GEN_73;
  wire [63:0]        regroupV0_hi_lo_lo_hi_lo_hi_lo_5;
  assign regroupV0_hi_lo_lo_hi_lo_hi_lo_5 = _GEN_73;
  wire [63:0]        regroupV0_hi_lo_lo_hi_lo_hi_lo_10;
  assign regroupV0_hi_lo_lo_hi_lo_hi_lo_10 = _GEN_73;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_lo_hi_lo_hi_lo;
  assign slideAddressGen_slideMaskInput_hi_lo_lo_hi_lo_hi_lo = _GEN_73;
  wire [63:0]        selectReadStageMask_hi_lo_lo_hi_lo_hi_lo;
  assign selectReadStageMask_hi_lo_lo_hi_lo_hi_lo = _GEN_73;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_lo_hi_lo;
  assign maskSplit_maskSelect_hi_lo_lo_hi_lo_hi_lo = _GEN_73;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_lo_hi_lo_1;
  assign maskSplit_maskSelect_hi_lo_lo_hi_lo_hi_lo_1 = _GEN_73;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_lo_hi_lo_2;
  assign maskSplit_maskSelect_hi_lo_lo_hi_lo_hi_lo_2 = _GEN_73;
  wire [63:0]        maskForDestination_hi_lo_lo_hi_lo_hi_lo;
  assign maskForDestination_hi_lo_lo_hi_lo_hi_lo = _GEN_73;
  wire [63:0]        _GEN_74 = {v0_151, v0_150};
  wire [63:0]        regroupV0_hi_lo_lo_hi_lo_hi_hi;
  assign regroupV0_hi_lo_lo_hi_lo_hi_hi = _GEN_74;
  wire [63:0]        regroupV0_hi_lo_lo_hi_lo_hi_hi_5;
  assign regroupV0_hi_lo_lo_hi_lo_hi_hi_5 = _GEN_74;
  wire [63:0]        regroupV0_hi_lo_lo_hi_lo_hi_hi_10;
  assign regroupV0_hi_lo_lo_hi_lo_hi_hi_10 = _GEN_74;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_lo_hi_lo_hi_hi;
  assign slideAddressGen_slideMaskInput_hi_lo_lo_hi_lo_hi_hi = _GEN_74;
  wire [63:0]        selectReadStageMask_hi_lo_lo_hi_lo_hi_hi;
  assign selectReadStageMask_hi_lo_lo_hi_lo_hi_hi = _GEN_74;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_lo_hi_hi;
  assign maskSplit_maskSelect_hi_lo_lo_hi_lo_hi_hi = _GEN_74;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_lo_hi_hi_1;
  assign maskSplit_maskSelect_hi_lo_lo_hi_lo_hi_hi_1 = _GEN_74;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_lo_hi_hi_2;
  assign maskSplit_maskSelect_hi_lo_lo_hi_lo_hi_hi_2 = _GEN_74;
  wire [63:0]        maskForDestination_hi_lo_lo_hi_lo_hi_hi;
  assign maskForDestination_hi_lo_lo_hi_lo_hi_hi = _GEN_74;
  wire [127:0]       regroupV0_hi_lo_lo_hi_lo_hi = {regroupV0_hi_lo_lo_hi_lo_hi_hi, regroupV0_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]       regroupV0_hi_lo_lo_hi_lo = {regroupV0_hi_lo_lo_hi_lo_hi, regroupV0_hi_lo_lo_hi_lo_lo};
  wire [63:0]        _GEN_75 = {v0_153, v0_152};
  wire [63:0]        regroupV0_hi_lo_lo_hi_hi_lo_lo;
  assign regroupV0_hi_lo_lo_hi_hi_lo_lo = _GEN_75;
  wire [63:0]        regroupV0_hi_lo_lo_hi_hi_lo_lo_5;
  assign regroupV0_hi_lo_lo_hi_hi_lo_lo_5 = _GEN_75;
  wire [63:0]        regroupV0_hi_lo_lo_hi_hi_lo_lo_10;
  assign regroupV0_hi_lo_lo_hi_hi_lo_lo_10 = _GEN_75;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_lo_hi_hi_lo_lo;
  assign slideAddressGen_slideMaskInput_hi_lo_lo_hi_hi_lo_lo = _GEN_75;
  wire [63:0]        selectReadStageMask_hi_lo_lo_hi_hi_lo_lo;
  assign selectReadStageMask_hi_lo_lo_hi_hi_lo_lo = _GEN_75;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_hi_lo_lo;
  assign maskSplit_maskSelect_hi_lo_lo_hi_hi_lo_lo = _GEN_75;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_hi_lo_lo_1;
  assign maskSplit_maskSelect_hi_lo_lo_hi_hi_lo_lo_1 = _GEN_75;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_hi_lo_lo_2;
  assign maskSplit_maskSelect_hi_lo_lo_hi_hi_lo_lo_2 = _GEN_75;
  wire [63:0]        maskForDestination_hi_lo_lo_hi_hi_lo_lo;
  assign maskForDestination_hi_lo_lo_hi_hi_lo_lo = _GEN_75;
  wire [63:0]        _GEN_76 = {v0_155, v0_154};
  wire [63:0]        regroupV0_hi_lo_lo_hi_hi_lo_hi;
  assign regroupV0_hi_lo_lo_hi_hi_lo_hi = _GEN_76;
  wire [63:0]        regroupV0_hi_lo_lo_hi_hi_lo_hi_5;
  assign regroupV0_hi_lo_lo_hi_hi_lo_hi_5 = _GEN_76;
  wire [63:0]        regroupV0_hi_lo_lo_hi_hi_lo_hi_10;
  assign regroupV0_hi_lo_lo_hi_hi_lo_hi_10 = _GEN_76;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_lo_hi_hi_lo_hi;
  assign slideAddressGen_slideMaskInput_hi_lo_lo_hi_hi_lo_hi = _GEN_76;
  wire [63:0]        selectReadStageMask_hi_lo_lo_hi_hi_lo_hi;
  assign selectReadStageMask_hi_lo_lo_hi_hi_lo_hi = _GEN_76;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_hi_lo_hi;
  assign maskSplit_maskSelect_hi_lo_lo_hi_hi_lo_hi = _GEN_76;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_hi_lo_hi_1;
  assign maskSplit_maskSelect_hi_lo_lo_hi_hi_lo_hi_1 = _GEN_76;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_hi_lo_hi_2;
  assign maskSplit_maskSelect_hi_lo_lo_hi_hi_lo_hi_2 = _GEN_76;
  wire [63:0]        maskForDestination_hi_lo_lo_hi_hi_lo_hi;
  assign maskForDestination_hi_lo_lo_hi_hi_lo_hi = _GEN_76;
  wire [127:0]       regroupV0_hi_lo_lo_hi_hi_lo = {regroupV0_hi_lo_lo_hi_hi_lo_hi, regroupV0_hi_lo_lo_hi_hi_lo_lo};
  wire [63:0]        _GEN_77 = {v0_157, v0_156};
  wire [63:0]        regroupV0_hi_lo_lo_hi_hi_hi_lo;
  assign regroupV0_hi_lo_lo_hi_hi_hi_lo = _GEN_77;
  wire [63:0]        regroupV0_hi_lo_lo_hi_hi_hi_lo_5;
  assign regroupV0_hi_lo_lo_hi_hi_hi_lo_5 = _GEN_77;
  wire [63:0]        regroupV0_hi_lo_lo_hi_hi_hi_lo_10;
  assign regroupV0_hi_lo_lo_hi_hi_hi_lo_10 = _GEN_77;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_lo_hi_hi_hi_lo;
  assign slideAddressGen_slideMaskInput_hi_lo_lo_hi_hi_hi_lo = _GEN_77;
  wire [63:0]        selectReadStageMask_hi_lo_lo_hi_hi_hi_lo;
  assign selectReadStageMask_hi_lo_lo_hi_hi_hi_lo = _GEN_77;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_hi_hi_lo;
  assign maskSplit_maskSelect_hi_lo_lo_hi_hi_hi_lo = _GEN_77;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_hi_hi_lo_1;
  assign maskSplit_maskSelect_hi_lo_lo_hi_hi_hi_lo_1 = _GEN_77;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_hi_hi_lo_2;
  assign maskSplit_maskSelect_hi_lo_lo_hi_hi_hi_lo_2 = _GEN_77;
  wire [63:0]        maskForDestination_hi_lo_lo_hi_hi_hi_lo;
  assign maskForDestination_hi_lo_lo_hi_hi_hi_lo = _GEN_77;
  wire [63:0]        _GEN_78 = {v0_159, v0_158};
  wire [63:0]        regroupV0_hi_lo_lo_hi_hi_hi_hi;
  assign regroupV0_hi_lo_lo_hi_hi_hi_hi = _GEN_78;
  wire [63:0]        regroupV0_hi_lo_lo_hi_hi_hi_hi_5;
  assign regroupV0_hi_lo_lo_hi_hi_hi_hi_5 = _GEN_78;
  wire [63:0]        regroupV0_hi_lo_lo_hi_hi_hi_hi_10;
  assign regroupV0_hi_lo_lo_hi_hi_hi_hi_10 = _GEN_78;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_lo_hi_hi_hi_hi;
  assign slideAddressGen_slideMaskInput_hi_lo_lo_hi_hi_hi_hi = _GEN_78;
  wire [63:0]        selectReadStageMask_hi_lo_lo_hi_hi_hi_hi;
  assign selectReadStageMask_hi_lo_lo_hi_hi_hi_hi = _GEN_78;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_hi_hi_hi;
  assign maskSplit_maskSelect_hi_lo_lo_hi_hi_hi_hi = _GEN_78;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_hi_hi_hi_1;
  assign maskSplit_maskSelect_hi_lo_lo_hi_hi_hi_hi_1 = _GEN_78;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_hi_hi_hi_2;
  assign maskSplit_maskSelect_hi_lo_lo_hi_hi_hi_hi_2 = _GEN_78;
  wire [63:0]        maskForDestination_hi_lo_lo_hi_hi_hi_hi;
  assign maskForDestination_hi_lo_lo_hi_hi_hi_hi = _GEN_78;
  wire [127:0]       regroupV0_hi_lo_lo_hi_hi_hi = {regroupV0_hi_lo_lo_hi_hi_hi_hi, regroupV0_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]       regroupV0_hi_lo_lo_hi_hi = {regroupV0_hi_lo_lo_hi_hi_hi, regroupV0_hi_lo_lo_hi_hi_lo};
  wire [511:0]       regroupV0_hi_lo_lo_hi = {regroupV0_hi_lo_lo_hi_hi, regroupV0_hi_lo_lo_hi_lo};
  wire [1023:0]      regroupV0_hi_lo_lo = {regroupV0_hi_lo_lo_hi, regroupV0_hi_lo_lo_lo};
  wire [63:0]        _GEN_79 = {v0_161, v0_160};
  wire [63:0]        regroupV0_hi_lo_hi_lo_lo_lo_lo;
  assign regroupV0_hi_lo_hi_lo_lo_lo_lo = _GEN_79;
  wire [63:0]        regroupV0_hi_lo_hi_lo_lo_lo_lo_5;
  assign regroupV0_hi_lo_hi_lo_lo_lo_lo_5 = _GEN_79;
  wire [63:0]        regroupV0_hi_lo_hi_lo_lo_lo_lo_10;
  assign regroupV0_hi_lo_hi_lo_lo_lo_lo_10 = _GEN_79;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_hi_lo_lo_lo_lo;
  assign slideAddressGen_slideMaskInput_hi_lo_hi_lo_lo_lo_lo = _GEN_79;
  wire [63:0]        selectReadStageMask_hi_lo_hi_lo_lo_lo_lo;
  assign selectReadStageMask_hi_lo_hi_lo_lo_lo_lo = _GEN_79;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_lo_lo_lo;
  assign maskSplit_maskSelect_hi_lo_hi_lo_lo_lo_lo = _GEN_79;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_lo_lo_lo_1;
  assign maskSplit_maskSelect_hi_lo_hi_lo_lo_lo_lo_1 = _GEN_79;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_lo_lo_lo_2;
  assign maskSplit_maskSelect_hi_lo_hi_lo_lo_lo_lo_2 = _GEN_79;
  wire [63:0]        maskForDestination_hi_lo_hi_lo_lo_lo_lo;
  assign maskForDestination_hi_lo_hi_lo_lo_lo_lo = _GEN_79;
  wire [63:0]        _GEN_80 = {v0_163, v0_162};
  wire [63:0]        regroupV0_hi_lo_hi_lo_lo_lo_hi;
  assign regroupV0_hi_lo_hi_lo_lo_lo_hi = _GEN_80;
  wire [63:0]        regroupV0_hi_lo_hi_lo_lo_lo_hi_5;
  assign regroupV0_hi_lo_hi_lo_lo_lo_hi_5 = _GEN_80;
  wire [63:0]        regroupV0_hi_lo_hi_lo_lo_lo_hi_10;
  assign regroupV0_hi_lo_hi_lo_lo_lo_hi_10 = _GEN_80;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_hi_lo_lo_lo_hi;
  assign slideAddressGen_slideMaskInput_hi_lo_hi_lo_lo_lo_hi = _GEN_80;
  wire [63:0]        selectReadStageMask_hi_lo_hi_lo_lo_lo_hi;
  assign selectReadStageMask_hi_lo_hi_lo_lo_lo_hi = _GEN_80;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_lo_lo_hi;
  assign maskSplit_maskSelect_hi_lo_hi_lo_lo_lo_hi = _GEN_80;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_lo_lo_hi_1;
  assign maskSplit_maskSelect_hi_lo_hi_lo_lo_lo_hi_1 = _GEN_80;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_lo_lo_hi_2;
  assign maskSplit_maskSelect_hi_lo_hi_lo_lo_lo_hi_2 = _GEN_80;
  wire [63:0]        maskForDestination_hi_lo_hi_lo_lo_lo_hi;
  assign maskForDestination_hi_lo_hi_lo_lo_lo_hi = _GEN_80;
  wire [127:0]       regroupV0_hi_lo_hi_lo_lo_lo = {regroupV0_hi_lo_hi_lo_lo_lo_hi, regroupV0_hi_lo_hi_lo_lo_lo_lo};
  wire [63:0]        _GEN_81 = {v0_165, v0_164};
  wire [63:0]        regroupV0_hi_lo_hi_lo_lo_hi_lo;
  assign regroupV0_hi_lo_hi_lo_lo_hi_lo = _GEN_81;
  wire [63:0]        regroupV0_hi_lo_hi_lo_lo_hi_lo_5;
  assign regroupV0_hi_lo_hi_lo_lo_hi_lo_5 = _GEN_81;
  wire [63:0]        regroupV0_hi_lo_hi_lo_lo_hi_lo_10;
  assign regroupV0_hi_lo_hi_lo_lo_hi_lo_10 = _GEN_81;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_hi_lo_lo_hi_lo;
  assign slideAddressGen_slideMaskInput_hi_lo_hi_lo_lo_hi_lo = _GEN_81;
  wire [63:0]        selectReadStageMask_hi_lo_hi_lo_lo_hi_lo;
  assign selectReadStageMask_hi_lo_hi_lo_lo_hi_lo = _GEN_81;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_lo_hi_lo;
  assign maskSplit_maskSelect_hi_lo_hi_lo_lo_hi_lo = _GEN_81;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_lo_hi_lo_1;
  assign maskSplit_maskSelect_hi_lo_hi_lo_lo_hi_lo_1 = _GEN_81;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_lo_hi_lo_2;
  assign maskSplit_maskSelect_hi_lo_hi_lo_lo_hi_lo_2 = _GEN_81;
  wire [63:0]        maskForDestination_hi_lo_hi_lo_lo_hi_lo;
  assign maskForDestination_hi_lo_hi_lo_lo_hi_lo = _GEN_81;
  wire [63:0]        _GEN_82 = {v0_167, v0_166};
  wire [63:0]        regroupV0_hi_lo_hi_lo_lo_hi_hi;
  assign regroupV0_hi_lo_hi_lo_lo_hi_hi = _GEN_82;
  wire [63:0]        regroupV0_hi_lo_hi_lo_lo_hi_hi_5;
  assign regroupV0_hi_lo_hi_lo_lo_hi_hi_5 = _GEN_82;
  wire [63:0]        regroupV0_hi_lo_hi_lo_lo_hi_hi_10;
  assign regroupV0_hi_lo_hi_lo_lo_hi_hi_10 = _GEN_82;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_hi_lo_lo_hi_hi;
  assign slideAddressGen_slideMaskInput_hi_lo_hi_lo_lo_hi_hi = _GEN_82;
  wire [63:0]        selectReadStageMask_hi_lo_hi_lo_lo_hi_hi;
  assign selectReadStageMask_hi_lo_hi_lo_lo_hi_hi = _GEN_82;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_lo_hi_hi;
  assign maskSplit_maskSelect_hi_lo_hi_lo_lo_hi_hi = _GEN_82;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_lo_hi_hi_1;
  assign maskSplit_maskSelect_hi_lo_hi_lo_lo_hi_hi_1 = _GEN_82;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_lo_hi_hi_2;
  assign maskSplit_maskSelect_hi_lo_hi_lo_lo_hi_hi_2 = _GEN_82;
  wire [63:0]        maskForDestination_hi_lo_hi_lo_lo_hi_hi;
  assign maskForDestination_hi_lo_hi_lo_lo_hi_hi = _GEN_82;
  wire [127:0]       regroupV0_hi_lo_hi_lo_lo_hi = {regroupV0_hi_lo_hi_lo_lo_hi_hi, regroupV0_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]       regroupV0_hi_lo_hi_lo_lo = {regroupV0_hi_lo_hi_lo_lo_hi, regroupV0_hi_lo_hi_lo_lo_lo};
  wire [63:0]        _GEN_83 = {v0_169, v0_168};
  wire [63:0]        regroupV0_hi_lo_hi_lo_hi_lo_lo;
  assign regroupV0_hi_lo_hi_lo_hi_lo_lo = _GEN_83;
  wire [63:0]        regroupV0_hi_lo_hi_lo_hi_lo_lo_5;
  assign regroupV0_hi_lo_hi_lo_hi_lo_lo_5 = _GEN_83;
  wire [63:0]        regroupV0_hi_lo_hi_lo_hi_lo_lo_10;
  assign regroupV0_hi_lo_hi_lo_hi_lo_lo_10 = _GEN_83;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_hi_lo_hi_lo_lo;
  assign slideAddressGen_slideMaskInput_hi_lo_hi_lo_hi_lo_lo = _GEN_83;
  wire [63:0]        selectReadStageMask_hi_lo_hi_lo_hi_lo_lo;
  assign selectReadStageMask_hi_lo_hi_lo_hi_lo_lo = _GEN_83;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_hi_lo_lo;
  assign maskSplit_maskSelect_hi_lo_hi_lo_hi_lo_lo = _GEN_83;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_hi_lo_lo_1;
  assign maskSplit_maskSelect_hi_lo_hi_lo_hi_lo_lo_1 = _GEN_83;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_hi_lo_lo_2;
  assign maskSplit_maskSelect_hi_lo_hi_lo_hi_lo_lo_2 = _GEN_83;
  wire [63:0]        maskForDestination_hi_lo_hi_lo_hi_lo_lo;
  assign maskForDestination_hi_lo_hi_lo_hi_lo_lo = _GEN_83;
  wire [63:0]        _GEN_84 = {v0_171, v0_170};
  wire [63:0]        regroupV0_hi_lo_hi_lo_hi_lo_hi;
  assign regroupV0_hi_lo_hi_lo_hi_lo_hi = _GEN_84;
  wire [63:0]        regroupV0_hi_lo_hi_lo_hi_lo_hi_5;
  assign regroupV0_hi_lo_hi_lo_hi_lo_hi_5 = _GEN_84;
  wire [63:0]        regroupV0_hi_lo_hi_lo_hi_lo_hi_10;
  assign regroupV0_hi_lo_hi_lo_hi_lo_hi_10 = _GEN_84;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_hi_lo_hi_lo_hi;
  assign slideAddressGen_slideMaskInput_hi_lo_hi_lo_hi_lo_hi = _GEN_84;
  wire [63:0]        selectReadStageMask_hi_lo_hi_lo_hi_lo_hi;
  assign selectReadStageMask_hi_lo_hi_lo_hi_lo_hi = _GEN_84;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_hi_lo_hi;
  assign maskSplit_maskSelect_hi_lo_hi_lo_hi_lo_hi = _GEN_84;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_hi_lo_hi_1;
  assign maskSplit_maskSelect_hi_lo_hi_lo_hi_lo_hi_1 = _GEN_84;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_hi_lo_hi_2;
  assign maskSplit_maskSelect_hi_lo_hi_lo_hi_lo_hi_2 = _GEN_84;
  wire [63:0]        maskForDestination_hi_lo_hi_lo_hi_lo_hi;
  assign maskForDestination_hi_lo_hi_lo_hi_lo_hi = _GEN_84;
  wire [127:0]       regroupV0_hi_lo_hi_lo_hi_lo = {regroupV0_hi_lo_hi_lo_hi_lo_hi, regroupV0_hi_lo_hi_lo_hi_lo_lo};
  wire [63:0]        _GEN_85 = {v0_173, v0_172};
  wire [63:0]        regroupV0_hi_lo_hi_lo_hi_hi_lo;
  assign regroupV0_hi_lo_hi_lo_hi_hi_lo = _GEN_85;
  wire [63:0]        regroupV0_hi_lo_hi_lo_hi_hi_lo_5;
  assign regroupV0_hi_lo_hi_lo_hi_hi_lo_5 = _GEN_85;
  wire [63:0]        regroupV0_hi_lo_hi_lo_hi_hi_lo_10;
  assign regroupV0_hi_lo_hi_lo_hi_hi_lo_10 = _GEN_85;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_hi_lo_hi_hi_lo;
  assign slideAddressGen_slideMaskInput_hi_lo_hi_lo_hi_hi_lo = _GEN_85;
  wire [63:0]        selectReadStageMask_hi_lo_hi_lo_hi_hi_lo;
  assign selectReadStageMask_hi_lo_hi_lo_hi_hi_lo = _GEN_85;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_hi_hi_lo;
  assign maskSplit_maskSelect_hi_lo_hi_lo_hi_hi_lo = _GEN_85;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_hi_hi_lo_1;
  assign maskSplit_maskSelect_hi_lo_hi_lo_hi_hi_lo_1 = _GEN_85;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_hi_hi_lo_2;
  assign maskSplit_maskSelect_hi_lo_hi_lo_hi_hi_lo_2 = _GEN_85;
  wire [63:0]        maskForDestination_hi_lo_hi_lo_hi_hi_lo;
  assign maskForDestination_hi_lo_hi_lo_hi_hi_lo = _GEN_85;
  wire [63:0]        _GEN_86 = {v0_175, v0_174};
  wire [63:0]        regroupV0_hi_lo_hi_lo_hi_hi_hi;
  assign regroupV0_hi_lo_hi_lo_hi_hi_hi = _GEN_86;
  wire [63:0]        regroupV0_hi_lo_hi_lo_hi_hi_hi_5;
  assign regroupV0_hi_lo_hi_lo_hi_hi_hi_5 = _GEN_86;
  wire [63:0]        regroupV0_hi_lo_hi_lo_hi_hi_hi_10;
  assign regroupV0_hi_lo_hi_lo_hi_hi_hi_10 = _GEN_86;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_hi_lo_hi_hi_hi;
  assign slideAddressGen_slideMaskInput_hi_lo_hi_lo_hi_hi_hi = _GEN_86;
  wire [63:0]        selectReadStageMask_hi_lo_hi_lo_hi_hi_hi;
  assign selectReadStageMask_hi_lo_hi_lo_hi_hi_hi = _GEN_86;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_hi_hi_hi;
  assign maskSplit_maskSelect_hi_lo_hi_lo_hi_hi_hi = _GEN_86;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_hi_hi_hi_1;
  assign maskSplit_maskSelect_hi_lo_hi_lo_hi_hi_hi_1 = _GEN_86;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_hi_hi_hi_2;
  assign maskSplit_maskSelect_hi_lo_hi_lo_hi_hi_hi_2 = _GEN_86;
  wire [63:0]        maskForDestination_hi_lo_hi_lo_hi_hi_hi;
  assign maskForDestination_hi_lo_hi_lo_hi_hi_hi = _GEN_86;
  wire [127:0]       regroupV0_hi_lo_hi_lo_hi_hi = {regroupV0_hi_lo_hi_lo_hi_hi_hi, regroupV0_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]       regroupV0_hi_lo_hi_lo_hi = {regroupV0_hi_lo_hi_lo_hi_hi, regroupV0_hi_lo_hi_lo_hi_lo};
  wire [511:0]       regroupV0_hi_lo_hi_lo = {regroupV0_hi_lo_hi_lo_hi, regroupV0_hi_lo_hi_lo_lo};
  wire [63:0]        _GEN_87 = {v0_177, v0_176};
  wire [63:0]        regroupV0_hi_lo_hi_hi_lo_lo_lo;
  assign regroupV0_hi_lo_hi_hi_lo_lo_lo = _GEN_87;
  wire [63:0]        regroupV0_hi_lo_hi_hi_lo_lo_lo_5;
  assign regroupV0_hi_lo_hi_hi_lo_lo_lo_5 = _GEN_87;
  wire [63:0]        regroupV0_hi_lo_hi_hi_lo_lo_lo_10;
  assign regroupV0_hi_lo_hi_hi_lo_lo_lo_10 = _GEN_87;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_hi_hi_lo_lo_lo;
  assign slideAddressGen_slideMaskInput_hi_lo_hi_hi_lo_lo_lo = _GEN_87;
  wire [63:0]        selectReadStageMask_hi_lo_hi_hi_lo_lo_lo;
  assign selectReadStageMask_hi_lo_hi_hi_lo_lo_lo = _GEN_87;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_lo_lo_lo;
  assign maskSplit_maskSelect_hi_lo_hi_hi_lo_lo_lo = _GEN_87;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_lo_lo_lo_1;
  assign maskSplit_maskSelect_hi_lo_hi_hi_lo_lo_lo_1 = _GEN_87;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_lo_lo_lo_2;
  assign maskSplit_maskSelect_hi_lo_hi_hi_lo_lo_lo_2 = _GEN_87;
  wire [63:0]        maskForDestination_hi_lo_hi_hi_lo_lo_lo;
  assign maskForDestination_hi_lo_hi_hi_lo_lo_lo = _GEN_87;
  wire [63:0]        _GEN_88 = {v0_179, v0_178};
  wire [63:0]        regroupV0_hi_lo_hi_hi_lo_lo_hi;
  assign regroupV0_hi_lo_hi_hi_lo_lo_hi = _GEN_88;
  wire [63:0]        regroupV0_hi_lo_hi_hi_lo_lo_hi_5;
  assign regroupV0_hi_lo_hi_hi_lo_lo_hi_5 = _GEN_88;
  wire [63:0]        regroupV0_hi_lo_hi_hi_lo_lo_hi_10;
  assign regroupV0_hi_lo_hi_hi_lo_lo_hi_10 = _GEN_88;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_hi_hi_lo_lo_hi;
  assign slideAddressGen_slideMaskInput_hi_lo_hi_hi_lo_lo_hi = _GEN_88;
  wire [63:0]        selectReadStageMask_hi_lo_hi_hi_lo_lo_hi;
  assign selectReadStageMask_hi_lo_hi_hi_lo_lo_hi = _GEN_88;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_lo_lo_hi;
  assign maskSplit_maskSelect_hi_lo_hi_hi_lo_lo_hi = _GEN_88;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_lo_lo_hi_1;
  assign maskSplit_maskSelect_hi_lo_hi_hi_lo_lo_hi_1 = _GEN_88;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_lo_lo_hi_2;
  assign maskSplit_maskSelect_hi_lo_hi_hi_lo_lo_hi_2 = _GEN_88;
  wire [63:0]        maskForDestination_hi_lo_hi_hi_lo_lo_hi;
  assign maskForDestination_hi_lo_hi_hi_lo_lo_hi = _GEN_88;
  wire [127:0]       regroupV0_hi_lo_hi_hi_lo_lo = {regroupV0_hi_lo_hi_hi_lo_lo_hi, regroupV0_hi_lo_hi_hi_lo_lo_lo};
  wire [63:0]        _GEN_89 = {v0_181, v0_180};
  wire [63:0]        regroupV0_hi_lo_hi_hi_lo_hi_lo;
  assign regroupV0_hi_lo_hi_hi_lo_hi_lo = _GEN_89;
  wire [63:0]        regroupV0_hi_lo_hi_hi_lo_hi_lo_5;
  assign regroupV0_hi_lo_hi_hi_lo_hi_lo_5 = _GEN_89;
  wire [63:0]        regroupV0_hi_lo_hi_hi_lo_hi_lo_10;
  assign regroupV0_hi_lo_hi_hi_lo_hi_lo_10 = _GEN_89;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_hi_hi_lo_hi_lo;
  assign slideAddressGen_slideMaskInput_hi_lo_hi_hi_lo_hi_lo = _GEN_89;
  wire [63:0]        selectReadStageMask_hi_lo_hi_hi_lo_hi_lo;
  assign selectReadStageMask_hi_lo_hi_hi_lo_hi_lo = _GEN_89;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_lo_hi_lo;
  assign maskSplit_maskSelect_hi_lo_hi_hi_lo_hi_lo = _GEN_89;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_lo_hi_lo_1;
  assign maskSplit_maskSelect_hi_lo_hi_hi_lo_hi_lo_1 = _GEN_89;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_lo_hi_lo_2;
  assign maskSplit_maskSelect_hi_lo_hi_hi_lo_hi_lo_2 = _GEN_89;
  wire [63:0]        maskForDestination_hi_lo_hi_hi_lo_hi_lo;
  assign maskForDestination_hi_lo_hi_hi_lo_hi_lo = _GEN_89;
  wire [63:0]        _GEN_90 = {v0_183, v0_182};
  wire [63:0]        regroupV0_hi_lo_hi_hi_lo_hi_hi;
  assign regroupV0_hi_lo_hi_hi_lo_hi_hi = _GEN_90;
  wire [63:0]        regroupV0_hi_lo_hi_hi_lo_hi_hi_5;
  assign regroupV0_hi_lo_hi_hi_lo_hi_hi_5 = _GEN_90;
  wire [63:0]        regroupV0_hi_lo_hi_hi_lo_hi_hi_10;
  assign regroupV0_hi_lo_hi_hi_lo_hi_hi_10 = _GEN_90;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_hi_hi_lo_hi_hi;
  assign slideAddressGen_slideMaskInput_hi_lo_hi_hi_lo_hi_hi = _GEN_90;
  wire [63:0]        selectReadStageMask_hi_lo_hi_hi_lo_hi_hi;
  assign selectReadStageMask_hi_lo_hi_hi_lo_hi_hi = _GEN_90;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_lo_hi_hi;
  assign maskSplit_maskSelect_hi_lo_hi_hi_lo_hi_hi = _GEN_90;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_lo_hi_hi_1;
  assign maskSplit_maskSelect_hi_lo_hi_hi_lo_hi_hi_1 = _GEN_90;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_lo_hi_hi_2;
  assign maskSplit_maskSelect_hi_lo_hi_hi_lo_hi_hi_2 = _GEN_90;
  wire [63:0]        maskForDestination_hi_lo_hi_hi_lo_hi_hi;
  assign maskForDestination_hi_lo_hi_hi_lo_hi_hi = _GEN_90;
  wire [127:0]       regroupV0_hi_lo_hi_hi_lo_hi = {regroupV0_hi_lo_hi_hi_lo_hi_hi, regroupV0_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]       regroupV0_hi_lo_hi_hi_lo = {regroupV0_hi_lo_hi_hi_lo_hi, regroupV0_hi_lo_hi_hi_lo_lo};
  wire [63:0]        _GEN_91 = {v0_185, v0_184};
  wire [63:0]        regroupV0_hi_lo_hi_hi_hi_lo_lo;
  assign regroupV0_hi_lo_hi_hi_hi_lo_lo = _GEN_91;
  wire [63:0]        regroupV0_hi_lo_hi_hi_hi_lo_lo_5;
  assign regroupV0_hi_lo_hi_hi_hi_lo_lo_5 = _GEN_91;
  wire [63:0]        regroupV0_hi_lo_hi_hi_hi_lo_lo_10;
  assign regroupV0_hi_lo_hi_hi_hi_lo_lo_10 = _GEN_91;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_hi_hi_hi_lo_lo;
  assign slideAddressGen_slideMaskInput_hi_lo_hi_hi_hi_lo_lo = _GEN_91;
  wire [63:0]        selectReadStageMask_hi_lo_hi_hi_hi_lo_lo;
  assign selectReadStageMask_hi_lo_hi_hi_hi_lo_lo = _GEN_91;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_hi_lo_lo;
  assign maskSplit_maskSelect_hi_lo_hi_hi_hi_lo_lo = _GEN_91;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_hi_lo_lo_1;
  assign maskSplit_maskSelect_hi_lo_hi_hi_hi_lo_lo_1 = _GEN_91;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_hi_lo_lo_2;
  assign maskSplit_maskSelect_hi_lo_hi_hi_hi_lo_lo_2 = _GEN_91;
  wire [63:0]        maskForDestination_hi_lo_hi_hi_hi_lo_lo;
  assign maskForDestination_hi_lo_hi_hi_hi_lo_lo = _GEN_91;
  wire [63:0]        _GEN_92 = {v0_187, v0_186};
  wire [63:0]        regroupV0_hi_lo_hi_hi_hi_lo_hi;
  assign regroupV0_hi_lo_hi_hi_hi_lo_hi = _GEN_92;
  wire [63:0]        regroupV0_hi_lo_hi_hi_hi_lo_hi_5;
  assign regroupV0_hi_lo_hi_hi_hi_lo_hi_5 = _GEN_92;
  wire [63:0]        regroupV0_hi_lo_hi_hi_hi_lo_hi_10;
  assign regroupV0_hi_lo_hi_hi_hi_lo_hi_10 = _GEN_92;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_hi_hi_hi_lo_hi;
  assign slideAddressGen_slideMaskInput_hi_lo_hi_hi_hi_lo_hi = _GEN_92;
  wire [63:0]        selectReadStageMask_hi_lo_hi_hi_hi_lo_hi;
  assign selectReadStageMask_hi_lo_hi_hi_hi_lo_hi = _GEN_92;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_hi_lo_hi;
  assign maskSplit_maskSelect_hi_lo_hi_hi_hi_lo_hi = _GEN_92;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_hi_lo_hi_1;
  assign maskSplit_maskSelect_hi_lo_hi_hi_hi_lo_hi_1 = _GEN_92;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_hi_lo_hi_2;
  assign maskSplit_maskSelect_hi_lo_hi_hi_hi_lo_hi_2 = _GEN_92;
  wire [63:0]        maskForDestination_hi_lo_hi_hi_hi_lo_hi;
  assign maskForDestination_hi_lo_hi_hi_hi_lo_hi = _GEN_92;
  wire [127:0]       regroupV0_hi_lo_hi_hi_hi_lo = {regroupV0_hi_lo_hi_hi_hi_lo_hi, regroupV0_hi_lo_hi_hi_hi_lo_lo};
  wire [63:0]        _GEN_93 = {v0_189, v0_188};
  wire [63:0]        regroupV0_hi_lo_hi_hi_hi_hi_lo;
  assign regroupV0_hi_lo_hi_hi_hi_hi_lo = _GEN_93;
  wire [63:0]        regroupV0_hi_lo_hi_hi_hi_hi_lo_5;
  assign regroupV0_hi_lo_hi_hi_hi_hi_lo_5 = _GEN_93;
  wire [63:0]        regroupV0_hi_lo_hi_hi_hi_hi_lo_10;
  assign regroupV0_hi_lo_hi_hi_hi_hi_lo_10 = _GEN_93;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_hi_hi_hi_hi_lo;
  assign slideAddressGen_slideMaskInput_hi_lo_hi_hi_hi_hi_lo = _GEN_93;
  wire [63:0]        selectReadStageMask_hi_lo_hi_hi_hi_hi_lo;
  assign selectReadStageMask_hi_lo_hi_hi_hi_hi_lo = _GEN_93;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_hi_hi_lo;
  assign maskSplit_maskSelect_hi_lo_hi_hi_hi_hi_lo = _GEN_93;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_hi_hi_lo_1;
  assign maskSplit_maskSelect_hi_lo_hi_hi_hi_hi_lo_1 = _GEN_93;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_hi_hi_lo_2;
  assign maskSplit_maskSelect_hi_lo_hi_hi_hi_hi_lo_2 = _GEN_93;
  wire [63:0]        maskForDestination_hi_lo_hi_hi_hi_hi_lo;
  assign maskForDestination_hi_lo_hi_hi_hi_hi_lo = _GEN_93;
  wire [63:0]        _GEN_94 = {v0_191, v0_190};
  wire [63:0]        regroupV0_hi_lo_hi_hi_hi_hi_hi;
  assign regroupV0_hi_lo_hi_hi_hi_hi_hi = _GEN_94;
  wire [63:0]        regroupV0_hi_lo_hi_hi_hi_hi_hi_5;
  assign regroupV0_hi_lo_hi_hi_hi_hi_hi_5 = _GEN_94;
  wire [63:0]        regroupV0_hi_lo_hi_hi_hi_hi_hi_10;
  assign regroupV0_hi_lo_hi_hi_hi_hi_hi_10 = _GEN_94;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_hi_hi_hi_hi_hi;
  assign slideAddressGen_slideMaskInput_hi_lo_hi_hi_hi_hi_hi = _GEN_94;
  wire [63:0]        selectReadStageMask_hi_lo_hi_hi_hi_hi_hi;
  assign selectReadStageMask_hi_lo_hi_hi_hi_hi_hi = _GEN_94;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_hi_hi_hi;
  assign maskSplit_maskSelect_hi_lo_hi_hi_hi_hi_hi = _GEN_94;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_hi_hi_hi_1;
  assign maskSplit_maskSelect_hi_lo_hi_hi_hi_hi_hi_1 = _GEN_94;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_hi_hi_hi_2;
  assign maskSplit_maskSelect_hi_lo_hi_hi_hi_hi_hi_2 = _GEN_94;
  wire [63:0]        maskForDestination_hi_lo_hi_hi_hi_hi_hi;
  assign maskForDestination_hi_lo_hi_hi_hi_hi_hi = _GEN_94;
  wire [127:0]       regroupV0_hi_lo_hi_hi_hi_hi = {regroupV0_hi_lo_hi_hi_hi_hi_hi, regroupV0_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]       regroupV0_hi_lo_hi_hi_hi = {regroupV0_hi_lo_hi_hi_hi_hi, regroupV0_hi_lo_hi_hi_hi_lo};
  wire [511:0]       regroupV0_hi_lo_hi_hi = {regroupV0_hi_lo_hi_hi_hi, regroupV0_hi_lo_hi_hi_lo};
  wire [1023:0]      regroupV0_hi_lo_hi = {regroupV0_hi_lo_hi_hi, regroupV0_hi_lo_hi_lo};
  wire [2047:0]      regroupV0_hi_lo = {regroupV0_hi_lo_hi, regroupV0_hi_lo_lo};
  wire [63:0]        _GEN_95 = {v0_193, v0_192};
  wire [63:0]        regroupV0_hi_hi_lo_lo_lo_lo_lo;
  assign regroupV0_hi_hi_lo_lo_lo_lo_lo = _GEN_95;
  wire [63:0]        regroupV0_hi_hi_lo_lo_lo_lo_lo_5;
  assign regroupV0_hi_hi_lo_lo_lo_lo_lo_5 = _GEN_95;
  wire [63:0]        regroupV0_hi_hi_lo_lo_lo_lo_lo_10;
  assign regroupV0_hi_hi_lo_lo_lo_lo_lo_10 = _GEN_95;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_lo_lo_lo_lo_lo;
  assign slideAddressGen_slideMaskInput_hi_hi_lo_lo_lo_lo_lo = _GEN_95;
  wire [63:0]        selectReadStageMask_hi_hi_lo_lo_lo_lo_lo;
  assign selectReadStageMask_hi_hi_lo_lo_lo_lo_lo = _GEN_95;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_lo_lo_lo;
  assign maskSplit_maskSelect_hi_hi_lo_lo_lo_lo_lo = _GEN_95;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_lo_lo_lo_1;
  assign maskSplit_maskSelect_hi_hi_lo_lo_lo_lo_lo_1 = _GEN_95;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_lo_lo_lo_2;
  assign maskSplit_maskSelect_hi_hi_lo_lo_lo_lo_lo_2 = _GEN_95;
  wire [63:0]        maskForDestination_hi_hi_lo_lo_lo_lo_lo;
  assign maskForDestination_hi_hi_lo_lo_lo_lo_lo = _GEN_95;
  wire [63:0]        _GEN_96 = {v0_195, v0_194};
  wire [63:0]        regroupV0_hi_hi_lo_lo_lo_lo_hi;
  assign regroupV0_hi_hi_lo_lo_lo_lo_hi = _GEN_96;
  wire [63:0]        regroupV0_hi_hi_lo_lo_lo_lo_hi_5;
  assign regroupV0_hi_hi_lo_lo_lo_lo_hi_5 = _GEN_96;
  wire [63:0]        regroupV0_hi_hi_lo_lo_lo_lo_hi_10;
  assign regroupV0_hi_hi_lo_lo_lo_lo_hi_10 = _GEN_96;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_lo_lo_lo_lo_hi;
  assign slideAddressGen_slideMaskInput_hi_hi_lo_lo_lo_lo_hi = _GEN_96;
  wire [63:0]        selectReadStageMask_hi_hi_lo_lo_lo_lo_hi;
  assign selectReadStageMask_hi_hi_lo_lo_lo_lo_hi = _GEN_96;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_lo_lo_hi;
  assign maskSplit_maskSelect_hi_hi_lo_lo_lo_lo_hi = _GEN_96;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_lo_lo_hi_1;
  assign maskSplit_maskSelect_hi_hi_lo_lo_lo_lo_hi_1 = _GEN_96;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_lo_lo_hi_2;
  assign maskSplit_maskSelect_hi_hi_lo_lo_lo_lo_hi_2 = _GEN_96;
  wire [63:0]        maskForDestination_hi_hi_lo_lo_lo_lo_hi;
  assign maskForDestination_hi_hi_lo_lo_lo_lo_hi = _GEN_96;
  wire [127:0]       regroupV0_hi_hi_lo_lo_lo_lo = {regroupV0_hi_hi_lo_lo_lo_lo_hi, regroupV0_hi_hi_lo_lo_lo_lo_lo};
  wire [63:0]        _GEN_97 = {v0_197, v0_196};
  wire [63:0]        regroupV0_hi_hi_lo_lo_lo_hi_lo;
  assign regroupV0_hi_hi_lo_lo_lo_hi_lo = _GEN_97;
  wire [63:0]        regroupV0_hi_hi_lo_lo_lo_hi_lo_5;
  assign regroupV0_hi_hi_lo_lo_lo_hi_lo_5 = _GEN_97;
  wire [63:0]        regroupV0_hi_hi_lo_lo_lo_hi_lo_10;
  assign regroupV0_hi_hi_lo_lo_lo_hi_lo_10 = _GEN_97;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_lo_lo_lo_hi_lo;
  assign slideAddressGen_slideMaskInput_hi_hi_lo_lo_lo_hi_lo = _GEN_97;
  wire [63:0]        selectReadStageMask_hi_hi_lo_lo_lo_hi_lo;
  assign selectReadStageMask_hi_hi_lo_lo_lo_hi_lo = _GEN_97;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_lo_hi_lo;
  assign maskSplit_maskSelect_hi_hi_lo_lo_lo_hi_lo = _GEN_97;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_lo_hi_lo_1;
  assign maskSplit_maskSelect_hi_hi_lo_lo_lo_hi_lo_1 = _GEN_97;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_lo_hi_lo_2;
  assign maskSplit_maskSelect_hi_hi_lo_lo_lo_hi_lo_2 = _GEN_97;
  wire [63:0]        maskForDestination_hi_hi_lo_lo_lo_hi_lo;
  assign maskForDestination_hi_hi_lo_lo_lo_hi_lo = _GEN_97;
  wire [63:0]        _GEN_98 = {v0_199, v0_198};
  wire [63:0]        regroupV0_hi_hi_lo_lo_lo_hi_hi;
  assign regroupV0_hi_hi_lo_lo_lo_hi_hi = _GEN_98;
  wire [63:0]        regroupV0_hi_hi_lo_lo_lo_hi_hi_5;
  assign regroupV0_hi_hi_lo_lo_lo_hi_hi_5 = _GEN_98;
  wire [63:0]        regroupV0_hi_hi_lo_lo_lo_hi_hi_10;
  assign regroupV0_hi_hi_lo_lo_lo_hi_hi_10 = _GEN_98;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_lo_lo_lo_hi_hi;
  assign slideAddressGen_slideMaskInput_hi_hi_lo_lo_lo_hi_hi = _GEN_98;
  wire [63:0]        selectReadStageMask_hi_hi_lo_lo_lo_hi_hi;
  assign selectReadStageMask_hi_hi_lo_lo_lo_hi_hi = _GEN_98;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_lo_hi_hi;
  assign maskSplit_maskSelect_hi_hi_lo_lo_lo_hi_hi = _GEN_98;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_lo_hi_hi_1;
  assign maskSplit_maskSelect_hi_hi_lo_lo_lo_hi_hi_1 = _GEN_98;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_lo_hi_hi_2;
  assign maskSplit_maskSelect_hi_hi_lo_lo_lo_hi_hi_2 = _GEN_98;
  wire [63:0]        maskForDestination_hi_hi_lo_lo_lo_hi_hi;
  assign maskForDestination_hi_hi_lo_lo_lo_hi_hi = _GEN_98;
  wire [127:0]       regroupV0_hi_hi_lo_lo_lo_hi = {regroupV0_hi_hi_lo_lo_lo_hi_hi, regroupV0_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]       regroupV0_hi_hi_lo_lo_lo = {regroupV0_hi_hi_lo_lo_lo_hi, regroupV0_hi_hi_lo_lo_lo_lo};
  wire [63:0]        _GEN_99 = {v0_201, v0_200};
  wire [63:0]        regroupV0_hi_hi_lo_lo_hi_lo_lo;
  assign regroupV0_hi_hi_lo_lo_hi_lo_lo = _GEN_99;
  wire [63:0]        regroupV0_hi_hi_lo_lo_hi_lo_lo_5;
  assign regroupV0_hi_hi_lo_lo_hi_lo_lo_5 = _GEN_99;
  wire [63:0]        regroupV0_hi_hi_lo_lo_hi_lo_lo_10;
  assign regroupV0_hi_hi_lo_lo_hi_lo_lo_10 = _GEN_99;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_lo_lo_hi_lo_lo;
  assign slideAddressGen_slideMaskInput_hi_hi_lo_lo_hi_lo_lo = _GEN_99;
  wire [63:0]        selectReadStageMask_hi_hi_lo_lo_hi_lo_lo;
  assign selectReadStageMask_hi_hi_lo_lo_hi_lo_lo = _GEN_99;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_hi_lo_lo;
  assign maskSplit_maskSelect_hi_hi_lo_lo_hi_lo_lo = _GEN_99;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_hi_lo_lo_1;
  assign maskSplit_maskSelect_hi_hi_lo_lo_hi_lo_lo_1 = _GEN_99;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_hi_lo_lo_2;
  assign maskSplit_maskSelect_hi_hi_lo_lo_hi_lo_lo_2 = _GEN_99;
  wire [63:0]        maskForDestination_hi_hi_lo_lo_hi_lo_lo;
  assign maskForDestination_hi_hi_lo_lo_hi_lo_lo = _GEN_99;
  wire [63:0]        _GEN_100 = {v0_203, v0_202};
  wire [63:0]        regroupV0_hi_hi_lo_lo_hi_lo_hi;
  assign regroupV0_hi_hi_lo_lo_hi_lo_hi = _GEN_100;
  wire [63:0]        regroupV0_hi_hi_lo_lo_hi_lo_hi_5;
  assign regroupV0_hi_hi_lo_lo_hi_lo_hi_5 = _GEN_100;
  wire [63:0]        regroupV0_hi_hi_lo_lo_hi_lo_hi_10;
  assign regroupV0_hi_hi_lo_lo_hi_lo_hi_10 = _GEN_100;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_lo_lo_hi_lo_hi;
  assign slideAddressGen_slideMaskInput_hi_hi_lo_lo_hi_lo_hi = _GEN_100;
  wire [63:0]        selectReadStageMask_hi_hi_lo_lo_hi_lo_hi;
  assign selectReadStageMask_hi_hi_lo_lo_hi_lo_hi = _GEN_100;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_hi_lo_hi;
  assign maskSplit_maskSelect_hi_hi_lo_lo_hi_lo_hi = _GEN_100;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_hi_lo_hi_1;
  assign maskSplit_maskSelect_hi_hi_lo_lo_hi_lo_hi_1 = _GEN_100;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_hi_lo_hi_2;
  assign maskSplit_maskSelect_hi_hi_lo_lo_hi_lo_hi_2 = _GEN_100;
  wire [63:0]        maskForDestination_hi_hi_lo_lo_hi_lo_hi;
  assign maskForDestination_hi_hi_lo_lo_hi_lo_hi = _GEN_100;
  wire [127:0]       regroupV0_hi_hi_lo_lo_hi_lo = {regroupV0_hi_hi_lo_lo_hi_lo_hi, regroupV0_hi_hi_lo_lo_hi_lo_lo};
  wire [63:0]        _GEN_101 = {v0_205, v0_204};
  wire [63:0]        regroupV0_hi_hi_lo_lo_hi_hi_lo;
  assign regroupV0_hi_hi_lo_lo_hi_hi_lo = _GEN_101;
  wire [63:0]        regroupV0_hi_hi_lo_lo_hi_hi_lo_5;
  assign regroupV0_hi_hi_lo_lo_hi_hi_lo_5 = _GEN_101;
  wire [63:0]        regroupV0_hi_hi_lo_lo_hi_hi_lo_10;
  assign regroupV0_hi_hi_lo_lo_hi_hi_lo_10 = _GEN_101;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_lo_lo_hi_hi_lo;
  assign slideAddressGen_slideMaskInput_hi_hi_lo_lo_hi_hi_lo = _GEN_101;
  wire [63:0]        selectReadStageMask_hi_hi_lo_lo_hi_hi_lo;
  assign selectReadStageMask_hi_hi_lo_lo_hi_hi_lo = _GEN_101;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_hi_hi_lo;
  assign maskSplit_maskSelect_hi_hi_lo_lo_hi_hi_lo = _GEN_101;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_hi_hi_lo_1;
  assign maskSplit_maskSelect_hi_hi_lo_lo_hi_hi_lo_1 = _GEN_101;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_hi_hi_lo_2;
  assign maskSplit_maskSelect_hi_hi_lo_lo_hi_hi_lo_2 = _GEN_101;
  wire [63:0]        maskForDestination_hi_hi_lo_lo_hi_hi_lo;
  assign maskForDestination_hi_hi_lo_lo_hi_hi_lo = _GEN_101;
  wire [63:0]        _GEN_102 = {v0_207, v0_206};
  wire [63:0]        regroupV0_hi_hi_lo_lo_hi_hi_hi;
  assign regroupV0_hi_hi_lo_lo_hi_hi_hi = _GEN_102;
  wire [63:0]        regroupV0_hi_hi_lo_lo_hi_hi_hi_5;
  assign regroupV0_hi_hi_lo_lo_hi_hi_hi_5 = _GEN_102;
  wire [63:0]        regroupV0_hi_hi_lo_lo_hi_hi_hi_10;
  assign regroupV0_hi_hi_lo_lo_hi_hi_hi_10 = _GEN_102;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_lo_lo_hi_hi_hi;
  assign slideAddressGen_slideMaskInput_hi_hi_lo_lo_hi_hi_hi = _GEN_102;
  wire [63:0]        selectReadStageMask_hi_hi_lo_lo_hi_hi_hi;
  assign selectReadStageMask_hi_hi_lo_lo_hi_hi_hi = _GEN_102;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_hi_hi_hi;
  assign maskSplit_maskSelect_hi_hi_lo_lo_hi_hi_hi = _GEN_102;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_hi_hi_hi_1;
  assign maskSplit_maskSelect_hi_hi_lo_lo_hi_hi_hi_1 = _GEN_102;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_hi_hi_hi_2;
  assign maskSplit_maskSelect_hi_hi_lo_lo_hi_hi_hi_2 = _GEN_102;
  wire [63:0]        maskForDestination_hi_hi_lo_lo_hi_hi_hi;
  assign maskForDestination_hi_hi_lo_lo_hi_hi_hi = _GEN_102;
  wire [127:0]       regroupV0_hi_hi_lo_lo_hi_hi = {regroupV0_hi_hi_lo_lo_hi_hi_hi, regroupV0_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]       regroupV0_hi_hi_lo_lo_hi = {regroupV0_hi_hi_lo_lo_hi_hi, regroupV0_hi_hi_lo_lo_hi_lo};
  wire [511:0]       regroupV0_hi_hi_lo_lo = {regroupV0_hi_hi_lo_lo_hi, regroupV0_hi_hi_lo_lo_lo};
  wire [63:0]        _GEN_103 = {v0_209, v0_208};
  wire [63:0]        regroupV0_hi_hi_lo_hi_lo_lo_lo;
  assign regroupV0_hi_hi_lo_hi_lo_lo_lo = _GEN_103;
  wire [63:0]        regroupV0_hi_hi_lo_hi_lo_lo_lo_5;
  assign regroupV0_hi_hi_lo_hi_lo_lo_lo_5 = _GEN_103;
  wire [63:0]        regroupV0_hi_hi_lo_hi_lo_lo_lo_10;
  assign regroupV0_hi_hi_lo_hi_lo_lo_lo_10 = _GEN_103;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_lo_hi_lo_lo_lo;
  assign slideAddressGen_slideMaskInput_hi_hi_lo_hi_lo_lo_lo = _GEN_103;
  wire [63:0]        selectReadStageMask_hi_hi_lo_hi_lo_lo_lo;
  assign selectReadStageMask_hi_hi_lo_hi_lo_lo_lo = _GEN_103;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_lo_lo_lo;
  assign maskSplit_maskSelect_hi_hi_lo_hi_lo_lo_lo = _GEN_103;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_lo_lo_lo_1;
  assign maskSplit_maskSelect_hi_hi_lo_hi_lo_lo_lo_1 = _GEN_103;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_lo_lo_lo_2;
  assign maskSplit_maskSelect_hi_hi_lo_hi_lo_lo_lo_2 = _GEN_103;
  wire [63:0]        maskForDestination_hi_hi_lo_hi_lo_lo_lo;
  assign maskForDestination_hi_hi_lo_hi_lo_lo_lo = _GEN_103;
  wire [63:0]        _GEN_104 = {v0_211, v0_210};
  wire [63:0]        regroupV0_hi_hi_lo_hi_lo_lo_hi;
  assign regroupV0_hi_hi_lo_hi_lo_lo_hi = _GEN_104;
  wire [63:0]        regroupV0_hi_hi_lo_hi_lo_lo_hi_5;
  assign regroupV0_hi_hi_lo_hi_lo_lo_hi_5 = _GEN_104;
  wire [63:0]        regroupV0_hi_hi_lo_hi_lo_lo_hi_10;
  assign regroupV0_hi_hi_lo_hi_lo_lo_hi_10 = _GEN_104;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_lo_hi_lo_lo_hi;
  assign slideAddressGen_slideMaskInput_hi_hi_lo_hi_lo_lo_hi = _GEN_104;
  wire [63:0]        selectReadStageMask_hi_hi_lo_hi_lo_lo_hi;
  assign selectReadStageMask_hi_hi_lo_hi_lo_lo_hi = _GEN_104;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_lo_lo_hi;
  assign maskSplit_maskSelect_hi_hi_lo_hi_lo_lo_hi = _GEN_104;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_lo_lo_hi_1;
  assign maskSplit_maskSelect_hi_hi_lo_hi_lo_lo_hi_1 = _GEN_104;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_lo_lo_hi_2;
  assign maskSplit_maskSelect_hi_hi_lo_hi_lo_lo_hi_2 = _GEN_104;
  wire [63:0]        maskForDestination_hi_hi_lo_hi_lo_lo_hi;
  assign maskForDestination_hi_hi_lo_hi_lo_lo_hi = _GEN_104;
  wire [127:0]       regroupV0_hi_hi_lo_hi_lo_lo = {regroupV0_hi_hi_lo_hi_lo_lo_hi, regroupV0_hi_hi_lo_hi_lo_lo_lo};
  wire [63:0]        _GEN_105 = {v0_213, v0_212};
  wire [63:0]        regroupV0_hi_hi_lo_hi_lo_hi_lo;
  assign regroupV0_hi_hi_lo_hi_lo_hi_lo = _GEN_105;
  wire [63:0]        regroupV0_hi_hi_lo_hi_lo_hi_lo_5;
  assign regroupV0_hi_hi_lo_hi_lo_hi_lo_5 = _GEN_105;
  wire [63:0]        regroupV0_hi_hi_lo_hi_lo_hi_lo_10;
  assign regroupV0_hi_hi_lo_hi_lo_hi_lo_10 = _GEN_105;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_lo_hi_lo_hi_lo;
  assign slideAddressGen_slideMaskInput_hi_hi_lo_hi_lo_hi_lo = _GEN_105;
  wire [63:0]        selectReadStageMask_hi_hi_lo_hi_lo_hi_lo;
  assign selectReadStageMask_hi_hi_lo_hi_lo_hi_lo = _GEN_105;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_lo_hi_lo;
  assign maskSplit_maskSelect_hi_hi_lo_hi_lo_hi_lo = _GEN_105;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_lo_hi_lo_1;
  assign maskSplit_maskSelect_hi_hi_lo_hi_lo_hi_lo_1 = _GEN_105;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_lo_hi_lo_2;
  assign maskSplit_maskSelect_hi_hi_lo_hi_lo_hi_lo_2 = _GEN_105;
  wire [63:0]        maskForDestination_hi_hi_lo_hi_lo_hi_lo;
  assign maskForDestination_hi_hi_lo_hi_lo_hi_lo = _GEN_105;
  wire [63:0]        _GEN_106 = {v0_215, v0_214};
  wire [63:0]        regroupV0_hi_hi_lo_hi_lo_hi_hi;
  assign regroupV0_hi_hi_lo_hi_lo_hi_hi = _GEN_106;
  wire [63:0]        regroupV0_hi_hi_lo_hi_lo_hi_hi_5;
  assign regroupV0_hi_hi_lo_hi_lo_hi_hi_5 = _GEN_106;
  wire [63:0]        regroupV0_hi_hi_lo_hi_lo_hi_hi_10;
  assign regroupV0_hi_hi_lo_hi_lo_hi_hi_10 = _GEN_106;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_lo_hi_lo_hi_hi;
  assign slideAddressGen_slideMaskInput_hi_hi_lo_hi_lo_hi_hi = _GEN_106;
  wire [63:0]        selectReadStageMask_hi_hi_lo_hi_lo_hi_hi;
  assign selectReadStageMask_hi_hi_lo_hi_lo_hi_hi = _GEN_106;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_lo_hi_hi;
  assign maskSplit_maskSelect_hi_hi_lo_hi_lo_hi_hi = _GEN_106;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_lo_hi_hi_1;
  assign maskSplit_maskSelect_hi_hi_lo_hi_lo_hi_hi_1 = _GEN_106;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_lo_hi_hi_2;
  assign maskSplit_maskSelect_hi_hi_lo_hi_lo_hi_hi_2 = _GEN_106;
  wire [63:0]        maskForDestination_hi_hi_lo_hi_lo_hi_hi;
  assign maskForDestination_hi_hi_lo_hi_lo_hi_hi = _GEN_106;
  wire [127:0]       regroupV0_hi_hi_lo_hi_lo_hi = {regroupV0_hi_hi_lo_hi_lo_hi_hi, regroupV0_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]       regroupV0_hi_hi_lo_hi_lo = {regroupV0_hi_hi_lo_hi_lo_hi, regroupV0_hi_hi_lo_hi_lo_lo};
  wire [63:0]        _GEN_107 = {v0_217, v0_216};
  wire [63:0]        regroupV0_hi_hi_lo_hi_hi_lo_lo;
  assign regroupV0_hi_hi_lo_hi_hi_lo_lo = _GEN_107;
  wire [63:0]        regroupV0_hi_hi_lo_hi_hi_lo_lo_5;
  assign regroupV0_hi_hi_lo_hi_hi_lo_lo_5 = _GEN_107;
  wire [63:0]        regroupV0_hi_hi_lo_hi_hi_lo_lo_10;
  assign regroupV0_hi_hi_lo_hi_hi_lo_lo_10 = _GEN_107;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_lo_hi_hi_lo_lo;
  assign slideAddressGen_slideMaskInput_hi_hi_lo_hi_hi_lo_lo = _GEN_107;
  wire [63:0]        selectReadStageMask_hi_hi_lo_hi_hi_lo_lo;
  assign selectReadStageMask_hi_hi_lo_hi_hi_lo_lo = _GEN_107;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_hi_lo_lo;
  assign maskSplit_maskSelect_hi_hi_lo_hi_hi_lo_lo = _GEN_107;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_hi_lo_lo_1;
  assign maskSplit_maskSelect_hi_hi_lo_hi_hi_lo_lo_1 = _GEN_107;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_hi_lo_lo_2;
  assign maskSplit_maskSelect_hi_hi_lo_hi_hi_lo_lo_2 = _GEN_107;
  wire [63:0]        maskForDestination_hi_hi_lo_hi_hi_lo_lo;
  assign maskForDestination_hi_hi_lo_hi_hi_lo_lo = _GEN_107;
  wire [63:0]        _GEN_108 = {v0_219, v0_218};
  wire [63:0]        regroupV0_hi_hi_lo_hi_hi_lo_hi;
  assign regroupV0_hi_hi_lo_hi_hi_lo_hi = _GEN_108;
  wire [63:0]        regroupV0_hi_hi_lo_hi_hi_lo_hi_5;
  assign regroupV0_hi_hi_lo_hi_hi_lo_hi_5 = _GEN_108;
  wire [63:0]        regroupV0_hi_hi_lo_hi_hi_lo_hi_10;
  assign regroupV0_hi_hi_lo_hi_hi_lo_hi_10 = _GEN_108;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_lo_hi_hi_lo_hi;
  assign slideAddressGen_slideMaskInput_hi_hi_lo_hi_hi_lo_hi = _GEN_108;
  wire [63:0]        selectReadStageMask_hi_hi_lo_hi_hi_lo_hi;
  assign selectReadStageMask_hi_hi_lo_hi_hi_lo_hi = _GEN_108;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_hi_lo_hi;
  assign maskSplit_maskSelect_hi_hi_lo_hi_hi_lo_hi = _GEN_108;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_hi_lo_hi_1;
  assign maskSplit_maskSelect_hi_hi_lo_hi_hi_lo_hi_1 = _GEN_108;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_hi_lo_hi_2;
  assign maskSplit_maskSelect_hi_hi_lo_hi_hi_lo_hi_2 = _GEN_108;
  wire [63:0]        maskForDestination_hi_hi_lo_hi_hi_lo_hi;
  assign maskForDestination_hi_hi_lo_hi_hi_lo_hi = _GEN_108;
  wire [127:0]       regroupV0_hi_hi_lo_hi_hi_lo = {regroupV0_hi_hi_lo_hi_hi_lo_hi, regroupV0_hi_hi_lo_hi_hi_lo_lo};
  wire [63:0]        _GEN_109 = {v0_221, v0_220};
  wire [63:0]        regroupV0_hi_hi_lo_hi_hi_hi_lo;
  assign regroupV0_hi_hi_lo_hi_hi_hi_lo = _GEN_109;
  wire [63:0]        regroupV0_hi_hi_lo_hi_hi_hi_lo_5;
  assign regroupV0_hi_hi_lo_hi_hi_hi_lo_5 = _GEN_109;
  wire [63:0]        regroupV0_hi_hi_lo_hi_hi_hi_lo_10;
  assign regroupV0_hi_hi_lo_hi_hi_hi_lo_10 = _GEN_109;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_lo_hi_hi_hi_lo;
  assign slideAddressGen_slideMaskInput_hi_hi_lo_hi_hi_hi_lo = _GEN_109;
  wire [63:0]        selectReadStageMask_hi_hi_lo_hi_hi_hi_lo;
  assign selectReadStageMask_hi_hi_lo_hi_hi_hi_lo = _GEN_109;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_hi_hi_lo;
  assign maskSplit_maskSelect_hi_hi_lo_hi_hi_hi_lo = _GEN_109;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_hi_hi_lo_1;
  assign maskSplit_maskSelect_hi_hi_lo_hi_hi_hi_lo_1 = _GEN_109;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_hi_hi_lo_2;
  assign maskSplit_maskSelect_hi_hi_lo_hi_hi_hi_lo_2 = _GEN_109;
  wire [63:0]        maskForDestination_hi_hi_lo_hi_hi_hi_lo;
  assign maskForDestination_hi_hi_lo_hi_hi_hi_lo = _GEN_109;
  wire [63:0]        _GEN_110 = {v0_223, v0_222};
  wire [63:0]        regroupV0_hi_hi_lo_hi_hi_hi_hi;
  assign regroupV0_hi_hi_lo_hi_hi_hi_hi = _GEN_110;
  wire [63:0]        regroupV0_hi_hi_lo_hi_hi_hi_hi_5;
  assign regroupV0_hi_hi_lo_hi_hi_hi_hi_5 = _GEN_110;
  wire [63:0]        regroupV0_hi_hi_lo_hi_hi_hi_hi_10;
  assign regroupV0_hi_hi_lo_hi_hi_hi_hi_10 = _GEN_110;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_lo_hi_hi_hi_hi;
  assign slideAddressGen_slideMaskInput_hi_hi_lo_hi_hi_hi_hi = _GEN_110;
  wire [63:0]        selectReadStageMask_hi_hi_lo_hi_hi_hi_hi;
  assign selectReadStageMask_hi_hi_lo_hi_hi_hi_hi = _GEN_110;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_hi_hi_hi;
  assign maskSplit_maskSelect_hi_hi_lo_hi_hi_hi_hi = _GEN_110;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_hi_hi_hi_1;
  assign maskSplit_maskSelect_hi_hi_lo_hi_hi_hi_hi_1 = _GEN_110;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_hi_hi_hi_2;
  assign maskSplit_maskSelect_hi_hi_lo_hi_hi_hi_hi_2 = _GEN_110;
  wire [63:0]        maskForDestination_hi_hi_lo_hi_hi_hi_hi;
  assign maskForDestination_hi_hi_lo_hi_hi_hi_hi = _GEN_110;
  wire [127:0]       regroupV0_hi_hi_lo_hi_hi_hi = {regroupV0_hi_hi_lo_hi_hi_hi_hi, regroupV0_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]       regroupV0_hi_hi_lo_hi_hi = {regroupV0_hi_hi_lo_hi_hi_hi, regroupV0_hi_hi_lo_hi_hi_lo};
  wire [511:0]       regroupV0_hi_hi_lo_hi = {regroupV0_hi_hi_lo_hi_hi, regroupV0_hi_hi_lo_hi_lo};
  wire [1023:0]      regroupV0_hi_hi_lo = {regroupV0_hi_hi_lo_hi, regroupV0_hi_hi_lo_lo};
  wire [63:0]        _GEN_111 = {v0_225, v0_224};
  wire [63:0]        regroupV0_hi_hi_hi_lo_lo_lo_lo;
  assign regroupV0_hi_hi_hi_lo_lo_lo_lo = _GEN_111;
  wire [63:0]        regroupV0_hi_hi_hi_lo_lo_lo_lo_5;
  assign regroupV0_hi_hi_hi_lo_lo_lo_lo_5 = _GEN_111;
  wire [63:0]        regroupV0_hi_hi_hi_lo_lo_lo_lo_10;
  assign regroupV0_hi_hi_hi_lo_lo_lo_lo_10 = _GEN_111;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_hi_lo_lo_lo_lo;
  assign slideAddressGen_slideMaskInput_hi_hi_hi_lo_lo_lo_lo = _GEN_111;
  wire [63:0]        selectReadStageMask_hi_hi_hi_lo_lo_lo_lo;
  assign selectReadStageMask_hi_hi_hi_lo_lo_lo_lo = _GEN_111;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_lo_lo_lo;
  assign maskSplit_maskSelect_hi_hi_hi_lo_lo_lo_lo = _GEN_111;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_lo_lo_lo_1;
  assign maskSplit_maskSelect_hi_hi_hi_lo_lo_lo_lo_1 = _GEN_111;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_lo_lo_lo_2;
  assign maskSplit_maskSelect_hi_hi_hi_lo_lo_lo_lo_2 = _GEN_111;
  wire [63:0]        maskForDestination_hi_hi_hi_lo_lo_lo_lo;
  assign maskForDestination_hi_hi_hi_lo_lo_lo_lo = _GEN_111;
  wire [63:0]        _GEN_112 = {v0_227, v0_226};
  wire [63:0]        regroupV0_hi_hi_hi_lo_lo_lo_hi;
  assign regroupV0_hi_hi_hi_lo_lo_lo_hi = _GEN_112;
  wire [63:0]        regroupV0_hi_hi_hi_lo_lo_lo_hi_5;
  assign regroupV0_hi_hi_hi_lo_lo_lo_hi_5 = _GEN_112;
  wire [63:0]        regroupV0_hi_hi_hi_lo_lo_lo_hi_10;
  assign regroupV0_hi_hi_hi_lo_lo_lo_hi_10 = _GEN_112;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_hi_lo_lo_lo_hi;
  assign slideAddressGen_slideMaskInput_hi_hi_hi_lo_lo_lo_hi = _GEN_112;
  wire [63:0]        selectReadStageMask_hi_hi_hi_lo_lo_lo_hi;
  assign selectReadStageMask_hi_hi_hi_lo_lo_lo_hi = _GEN_112;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_lo_lo_hi;
  assign maskSplit_maskSelect_hi_hi_hi_lo_lo_lo_hi = _GEN_112;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_lo_lo_hi_1;
  assign maskSplit_maskSelect_hi_hi_hi_lo_lo_lo_hi_1 = _GEN_112;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_lo_lo_hi_2;
  assign maskSplit_maskSelect_hi_hi_hi_lo_lo_lo_hi_2 = _GEN_112;
  wire [63:0]        maskForDestination_hi_hi_hi_lo_lo_lo_hi;
  assign maskForDestination_hi_hi_hi_lo_lo_lo_hi = _GEN_112;
  wire [127:0]       regroupV0_hi_hi_hi_lo_lo_lo = {regroupV0_hi_hi_hi_lo_lo_lo_hi, regroupV0_hi_hi_hi_lo_lo_lo_lo};
  wire [63:0]        _GEN_113 = {v0_229, v0_228};
  wire [63:0]        regroupV0_hi_hi_hi_lo_lo_hi_lo;
  assign regroupV0_hi_hi_hi_lo_lo_hi_lo = _GEN_113;
  wire [63:0]        regroupV0_hi_hi_hi_lo_lo_hi_lo_5;
  assign regroupV0_hi_hi_hi_lo_lo_hi_lo_5 = _GEN_113;
  wire [63:0]        regroupV0_hi_hi_hi_lo_lo_hi_lo_10;
  assign regroupV0_hi_hi_hi_lo_lo_hi_lo_10 = _GEN_113;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_hi_lo_lo_hi_lo;
  assign slideAddressGen_slideMaskInput_hi_hi_hi_lo_lo_hi_lo = _GEN_113;
  wire [63:0]        selectReadStageMask_hi_hi_hi_lo_lo_hi_lo;
  assign selectReadStageMask_hi_hi_hi_lo_lo_hi_lo = _GEN_113;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_lo_hi_lo;
  assign maskSplit_maskSelect_hi_hi_hi_lo_lo_hi_lo = _GEN_113;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_lo_hi_lo_1;
  assign maskSplit_maskSelect_hi_hi_hi_lo_lo_hi_lo_1 = _GEN_113;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_lo_hi_lo_2;
  assign maskSplit_maskSelect_hi_hi_hi_lo_lo_hi_lo_2 = _GEN_113;
  wire [63:0]        maskForDestination_hi_hi_hi_lo_lo_hi_lo;
  assign maskForDestination_hi_hi_hi_lo_lo_hi_lo = _GEN_113;
  wire [63:0]        _GEN_114 = {v0_231, v0_230};
  wire [63:0]        regroupV0_hi_hi_hi_lo_lo_hi_hi;
  assign regroupV0_hi_hi_hi_lo_lo_hi_hi = _GEN_114;
  wire [63:0]        regroupV0_hi_hi_hi_lo_lo_hi_hi_5;
  assign regroupV0_hi_hi_hi_lo_lo_hi_hi_5 = _GEN_114;
  wire [63:0]        regroupV0_hi_hi_hi_lo_lo_hi_hi_10;
  assign regroupV0_hi_hi_hi_lo_lo_hi_hi_10 = _GEN_114;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_hi_lo_lo_hi_hi;
  assign slideAddressGen_slideMaskInput_hi_hi_hi_lo_lo_hi_hi = _GEN_114;
  wire [63:0]        selectReadStageMask_hi_hi_hi_lo_lo_hi_hi;
  assign selectReadStageMask_hi_hi_hi_lo_lo_hi_hi = _GEN_114;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_lo_hi_hi;
  assign maskSplit_maskSelect_hi_hi_hi_lo_lo_hi_hi = _GEN_114;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_lo_hi_hi_1;
  assign maskSplit_maskSelect_hi_hi_hi_lo_lo_hi_hi_1 = _GEN_114;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_lo_hi_hi_2;
  assign maskSplit_maskSelect_hi_hi_hi_lo_lo_hi_hi_2 = _GEN_114;
  wire [63:0]        maskForDestination_hi_hi_hi_lo_lo_hi_hi;
  assign maskForDestination_hi_hi_hi_lo_lo_hi_hi = _GEN_114;
  wire [127:0]       regroupV0_hi_hi_hi_lo_lo_hi = {regroupV0_hi_hi_hi_lo_lo_hi_hi, regroupV0_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]       regroupV0_hi_hi_hi_lo_lo = {regroupV0_hi_hi_hi_lo_lo_hi, regroupV0_hi_hi_hi_lo_lo_lo};
  wire [63:0]        _GEN_115 = {v0_233, v0_232};
  wire [63:0]        regroupV0_hi_hi_hi_lo_hi_lo_lo;
  assign regroupV0_hi_hi_hi_lo_hi_lo_lo = _GEN_115;
  wire [63:0]        regroupV0_hi_hi_hi_lo_hi_lo_lo_5;
  assign regroupV0_hi_hi_hi_lo_hi_lo_lo_5 = _GEN_115;
  wire [63:0]        regroupV0_hi_hi_hi_lo_hi_lo_lo_10;
  assign regroupV0_hi_hi_hi_lo_hi_lo_lo_10 = _GEN_115;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_hi_lo_hi_lo_lo;
  assign slideAddressGen_slideMaskInput_hi_hi_hi_lo_hi_lo_lo = _GEN_115;
  wire [63:0]        selectReadStageMask_hi_hi_hi_lo_hi_lo_lo;
  assign selectReadStageMask_hi_hi_hi_lo_hi_lo_lo = _GEN_115;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_hi_lo_lo;
  assign maskSplit_maskSelect_hi_hi_hi_lo_hi_lo_lo = _GEN_115;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_hi_lo_lo_1;
  assign maskSplit_maskSelect_hi_hi_hi_lo_hi_lo_lo_1 = _GEN_115;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_hi_lo_lo_2;
  assign maskSplit_maskSelect_hi_hi_hi_lo_hi_lo_lo_2 = _GEN_115;
  wire [63:0]        maskForDestination_hi_hi_hi_lo_hi_lo_lo;
  assign maskForDestination_hi_hi_hi_lo_hi_lo_lo = _GEN_115;
  wire [63:0]        _GEN_116 = {v0_235, v0_234};
  wire [63:0]        regroupV0_hi_hi_hi_lo_hi_lo_hi;
  assign regroupV0_hi_hi_hi_lo_hi_lo_hi = _GEN_116;
  wire [63:0]        regroupV0_hi_hi_hi_lo_hi_lo_hi_5;
  assign regroupV0_hi_hi_hi_lo_hi_lo_hi_5 = _GEN_116;
  wire [63:0]        regroupV0_hi_hi_hi_lo_hi_lo_hi_10;
  assign regroupV0_hi_hi_hi_lo_hi_lo_hi_10 = _GEN_116;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_hi_lo_hi_lo_hi;
  assign slideAddressGen_slideMaskInput_hi_hi_hi_lo_hi_lo_hi = _GEN_116;
  wire [63:0]        selectReadStageMask_hi_hi_hi_lo_hi_lo_hi;
  assign selectReadStageMask_hi_hi_hi_lo_hi_lo_hi = _GEN_116;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_hi_lo_hi;
  assign maskSplit_maskSelect_hi_hi_hi_lo_hi_lo_hi = _GEN_116;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_hi_lo_hi_1;
  assign maskSplit_maskSelect_hi_hi_hi_lo_hi_lo_hi_1 = _GEN_116;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_hi_lo_hi_2;
  assign maskSplit_maskSelect_hi_hi_hi_lo_hi_lo_hi_2 = _GEN_116;
  wire [63:0]        maskForDestination_hi_hi_hi_lo_hi_lo_hi;
  assign maskForDestination_hi_hi_hi_lo_hi_lo_hi = _GEN_116;
  wire [127:0]       regroupV0_hi_hi_hi_lo_hi_lo = {regroupV0_hi_hi_hi_lo_hi_lo_hi, regroupV0_hi_hi_hi_lo_hi_lo_lo};
  wire [63:0]        _GEN_117 = {v0_237, v0_236};
  wire [63:0]        regroupV0_hi_hi_hi_lo_hi_hi_lo;
  assign regroupV0_hi_hi_hi_lo_hi_hi_lo = _GEN_117;
  wire [63:0]        regroupV0_hi_hi_hi_lo_hi_hi_lo_5;
  assign regroupV0_hi_hi_hi_lo_hi_hi_lo_5 = _GEN_117;
  wire [63:0]        regroupV0_hi_hi_hi_lo_hi_hi_lo_10;
  assign regroupV0_hi_hi_hi_lo_hi_hi_lo_10 = _GEN_117;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_hi_lo_hi_hi_lo;
  assign slideAddressGen_slideMaskInput_hi_hi_hi_lo_hi_hi_lo = _GEN_117;
  wire [63:0]        selectReadStageMask_hi_hi_hi_lo_hi_hi_lo;
  assign selectReadStageMask_hi_hi_hi_lo_hi_hi_lo = _GEN_117;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_hi_hi_lo;
  assign maskSplit_maskSelect_hi_hi_hi_lo_hi_hi_lo = _GEN_117;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_hi_hi_lo_1;
  assign maskSplit_maskSelect_hi_hi_hi_lo_hi_hi_lo_1 = _GEN_117;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_hi_hi_lo_2;
  assign maskSplit_maskSelect_hi_hi_hi_lo_hi_hi_lo_2 = _GEN_117;
  wire [63:0]        maskForDestination_hi_hi_hi_lo_hi_hi_lo;
  assign maskForDestination_hi_hi_hi_lo_hi_hi_lo = _GEN_117;
  wire [63:0]        _GEN_118 = {v0_239, v0_238};
  wire [63:0]        regroupV0_hi_hi_hi_lo_hi_hi_hi;
  assign regroupV0_hi_hi_hi_lo_hi_hi_hi = _GEN_118;
  wire [63:0]        regroupV0_hi_hi_hi_lo_hi_hi_hi_5;
  assign regroupV0_hi_hi_hi_lo_hi_hi_hi_5 = _GEN_118;
  wire [63:0]        regroupV0_hi_hi_hi_lo_hi_hi_hi_10;
  assign regroupV0_hi_hi_hi_lo_hi_hi_hi_10 = _GEN_118;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_hi_lo_hi_hi_hi;
  assign slideAddressGen_slideMaskInput_hi_hi_hi_lo_hi_hi_hi = _GEN_118;
  wire [63:0]        selectReadStageMask_hi_hi_hi_lo_hi_hi_hi;
  assign selectReadStageMask_hi_hi_hi_lo_hi_hi_hi = _GEN_118;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_hi_hi_hi;
  assign maskSplit_maskSelect_hi_hi_hi_lo_hi_hi_hi = _GEN_118;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_hi_hi_hi_1;
  assign maskSplit_maskSelect_hi_hi_hi_lo_hi_hi_hi_1 = _GEN_118;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_hi_hi_hi_2;
  assign maskSplit_maskSelect_hi_hi_hi_lo_hi_hi_hi_2 = _GEN_118;
  wire [63:0]        maskForDestination_hi_hi_hi_lo_hi_hi_hi;
  assign maskForDestination_hi_hi_hi_lo_hi_hi_hi = _GEN_118;
  wire [127:0]       regroupV0_hi_hi_hi_lo_hi_hi = {regroupV0_hi_hi_hi_lo_hi_hi_hi, regroupV0_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]       regroupV0_hi_hi_hi_lo_hi = {regroupV0_hi_hi_hi_lo_hi_hi, regroupV0_hi_hi_hi_lo_hi_lo};
  wire [511:0]       regroupV0_hi_hi_hi_lo = {regroupV0_hi_hi_hi_lo_hi, regroupV0_hi_hi_hi_lo_lo};
  wire [63:0]        _GEN_119 = {v0_241, v0_240};
  wire [63:0]        regroupV0_hi_hi_hi_hi_lo_lo_lo;
  assign regroupV0_hi_hi_hi_hi_lo_lo_lo = _GEN_119;
  wire [63:0]        regroupV0_hi_hi_hi_hi_lo_lo_lo_5;
  assign regroupV0_hi_hi_hi_hi_lo_lo_lo_5 = _GEN_119;
  wire [63:0]        regroupV0_hi_hi_hi_hi_lo_lo_lo_10;
  assign regroupV0_hi_hi_hi_hi_lo_lo_lo_10 = _GEN_119;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_hi_hi_lo_lo_lo;
  assign slideAddressGen_slideMaskInput_hi_hi_hi_hi_lo_lo_lo = _GEN_119;
  wire [63:0]        selectReadStageMask_hi_hi_hi_hi_lo_lo_lo;
  assign selectReadStageMask_hi_hi_hi_hi_lo_lo_lo = _GEN_119;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_lo_lo_lo;
  assign maskSplit_maskSelect_hi_hi_hi_hi_lo_lo_lo = _GEN_119;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_lo_lo_lo_1;
  assign maskSplit_maskSelect_hi_hi_hi_hi_lo_lo_lo_1 = _GEN_119;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_lo_lo_lo_2;
  assign maskSplit_maskSelect_hi_hi_hi_hi_lo_lo_lo_2 = _GEN_119;
  wire [63:0]        maskForDestination_hi_hi_hi_hi_lo_lo_lo;
  assign maskForDestination_hi_hi_hi_hi_lo_lo_lo = _GEN_119;
  wire [63:0]        _GEN_120 = {v0_243, v0_242};
  wire [63:0]        regroupV0_hi_hi_hi_hi_lo_lo_hi;
  assign regroupV0_hi_hi_hi_hi_lo_lo_hi = _GEN_120;
  wire [63:0]        regroupV0_hi_hi_hi_hi_lo_lo_hi_5;
  assign regroupV0_hi_hi_hi_hi_lo_lo_hi_5 = _GEN_120;
  wire [63:0]        regroupV0_hi_hi_hi_hi_lo_lo_hi_10;
  assign regroupV0_hi_hi_hi_hi_lo_lo_hi_10 = _GEN_120;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_hi_hi_lo_lo_hi;
  assign slideAddressGen_slideMaskInput_hi_hi_hi_hi_lo_lo_hi = _GEN_120;
  wire [63:0]        selectReadStageMask_hi_hi_hi_hi_lo_lo_hi;
  assign selectReadStageMask_hi_hi_hi_hi_lo_lo_hi = _GEN_120;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_lo_lo_hi;
  assign maskSplit_maskSelect_hi_hi_hi_hi_lo_lo_hi = _GEN_120;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_lo_lo_hi_1;
  assign maskSplit_maskSelect_hi_hi_hi_hi_lo_lo_hi_1 = _GEN_120;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_lo_lo_hi_2;
  assign maskSplit_maskSelect_hi_hi_hi_hi_lo_lo_hi_2 = _GEN_120;
  wire [63:0]        maskForDestination_hi_hi_hi_hi_lo_lo_hi;
  assign maskForDestination_hi_hi_hi_hi_lo_lo_hi = _GEN_120;
  wire [127:0]       regroupV0_hi_hi_hi_hi_lo_lo = {regroupV0_hi_hi_hi_hi_lo_lo_hi, regroupV0_hi_hi_hi_hi_lo_lo_lo};
  wire [63:0]        _GEN_121 = {v0_245, v0_244};
  wire [63:0]        regroupV0_hi_hi_hi_hi_lo_hi_lo;
  assign regroupV0_hi_hi_hi_hi_lo_hi_lo = _GEN_121;
  wire [63:0]        regroupV0_hi_hi_hi_hi_lo_hi_lo_5;
  assign regroupV0_hi_hi_hi_hi_lo_hi_lo_5 = _GEN_121;
  wire [63:0]        regroupV0_hi_hi_hi_hi_lo_hi_lo_10;
  assign regroupV0_hi_hi_hi_hi_lo_hi_lo_10 = _GEN_121;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_hi_hi_lo_hi_lo;
  assign slideAddressGen_slideMaskInput_hi_hi_hi_hi_lo_hi_lo = _GEN_121;
  wire [63:0]        selectReadStageMask_hi_hi_hi_hi_lo_hi_lo;
  assign selectReadStageMask_hi_hi_hi_hi_lo_hi_lo = _GEN_121;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_lo_hi_lo;
  assign maskSplit_maskSelect_hi_hi_hi_hi_lo_hi_lo = _GEN_121;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_lo_hi_lo_1;
  assign maskSplit_maskSelect_hi_hi_hi_hi_lo_hi_lo_1 = _GEN_121;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_lo_hi_lo_2;
  assign maskSplit_maskSelect_hi_hi_hi_hi_lo_hi_lo_2 = _GEN_121;
  wire [63:0]        maskForDestination_hi_hi_hi_hi_lo_hi_lo;
  assign maskForDestination_hi_hi_hi_hi_lo_hi_lo = _GEN_121;
  wire [63:0]        _GEN_122 = {v0_247, v0_246};
  wire [63:0]        regroupV0_hi_hi_hi_hi_lo_hi_hi;
  assign regroupV0_hi_hi_hi_hi_lo_hi_hi = _GEN_122;
  wire [63:0]        regroupV0_hi_hi_hi_hi_lo_hi_hi_5;
  assign regroupV0_hi_hi_hi_hi_lo_hi_hi_5 = _GEN_122;
  wire [63:0]        regroupV0_hi_hi_hi_hi_lo_hi_hi_10;
  assign regroupV0_hi_hi_hi_hi_lo_hi_hi_10 = _GEN_122;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_hi_hi_lo_hi_hi;
  assign slideAddressGen_slideMaskInput_hi_hi_hi_hi_lo_hi_hi = _GEN_122;
  wire [63:0]        selectReadStageMask_hi_hi_hi_hi_lo_hi_hi;
  assign selectReadStageMask_hi_hi_hi_hi_lo_hi_hi = _GEN_122;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_lo_hi_hi;
  assign maskSplit_maskSelect_hi_hi_hi_hi_lo_hi_hi = _GEN_122;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_lo_hi_hi_1;
  assign maskSplit_maskSelect_hi_hi_hi_hi_lo_hi_hi_1 = _GEN_122;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_lo_hi_hi_2;
  assign maskSplit_maskSelect_hi_hi_hi_hi_lo_hi_hi_2 = _GEN_122;
  wire [63:0]        maskForDestination_hi_hi_hi_hi_lo_hi_hi;
  assign maskForDestination_hi_hi_hi_hi_lo_hi_hi = _GEN_122;
  wire [127:0]       regroupV0_hi_hi_hi_hi_lo_hi = {regroupV0_hi_hi_hi_hi_lo_hi_hi, regroupV0_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]       regroupV0_hi_hi_hi_hi_lo = {regroupV0_hi_hi_hi_hi_lo_hi, regroupV0_hi_hi_hi_hi_lo_lo};
  wire [63:0]        _GEN_123 = {v0_249, v0_248};
  wire [63:0]        regroupV0_hi_hi_hi_hi_hi_lo_lo;
  assign regroupV0_hi_hi_hi_hi_hi_lo_lo = _GEN_123;
  wire [63:0]        regroupV0_hi_hi_hi_hi_hi_lo_lo_5;
  assign regroupV0_hi_hi_hi_hi_hi_lo_lo_5 = _GEN_123;
  wire [63:0]        regroupV0_hi_hi_hi_hi_hi_lo_lo_10;
  assign regroupV0_hi_hi_hi_hi_hi_lo_lo_10 = _GEN_123;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_hi_hi_hi_lo_lo;
  assign slideAddressGen_slideMaskInput_hi_hi_hi_hi_hi_lo_lo = _GEN_123;
  wire [63:0]        selectReadStageMask_hi_hi_hi_hi_hi_lo_lo;
  assign selectReadStageMask_hi_hi_hi_hi_hi_lo_lo = _GEN_123;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_hi_lo_lo;
  assign maskSplit_maskSelect_hi_hi_hi_hi_hi_lo_lo = _GEN_123;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_hi_lo_lo_1;
  assign maskSplit_maskSelect_hi_hi_hi_hi_hi_lo_lo_1 = _GEN_123;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_hi_lo_lo_2;
  assign maskSplit_maskSelect_hi_hi_hi_hi_hi_lo_lo_2 = _GEN_123;
  wire [63:0]        maskForDestination_hi_hi_hi_hi_hi_lo_lo;
  assign maskForDestination_hi_hi_hi_hi_hi_lo_lo = _GEN_123;
  wire [63:0]        _GEN_124 = {v0_251, v0_250};
  wire [63:0]        regroupV0_hi_hi_hi_hi_hi_lo_hi;
  assign regroupV0_hi_hi_hi_hi_hi_lo_hi = _GEN_124;
  wire [63:0]        regroupV0_hi_hi_hi_hi_hi_lo_hi_5;
  assign regroupV0_hi_hi_hi_hi_hi_lo_hi_5 = _GEN_124;
  wire [63:0]        regroupV0_hi_hi_hi_hi_hi_lo_hi_10;
  assign regroupV0_hi_hi_hi_hi_hi_lo_hi_10 = _GEN_124;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_hi_hi_hi_lo_hi;
  assign slideAddressGen_slideMaskInput_hi_hi_hi_hi_hi_lo_hi = _GEN_124;
  wire [63:0]        selectReadStageMask_hi_hi_hi_hi_hi_lo_hi;
  assign selectReadStageMask_hi_hi_hi_hi_hi_lo_hi = _GEN_124;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_hi_lo_hi;
  assign maskSplit_maskSelect_hi_hi_hi_hi_hi_lo_hi = _GEN_124;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_hi_lo_hi_1;
  assign maskSplit_maskSelect_hi_hi_hi_hi_hi_lo_hi_1 = _GEN_124;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_hi_lo_hi_2;
  assign maskSplit_maskSelect_hi_hi_hi_hi_hi_lo_hi_2 = _GEN_124;
  wire [63:0]        maskForDestination_hi_hi_hi_hi_hi_lo_hi;
  assign maskForDestination_hi_hi_hi_hi_hi_lo_hi = _GEN_124;
  wire [127:0]       regroupV0_hi_hi_hi_hi_hi_lo = {regroupV0_hi_hi_hi_hi_hi_lo_hi, regroupV0_hi_hi_hi_hi_hi_lo_lo};
  wire [63:0]        _GEN_125 = {v0_253, v0_252};
  wire [63:0]        regroupV0_hi_hi_hi_hi_hi_hi_lo;
  assign regroupV0_hi_hi_hi_hi_hi_hi_lo = _GEN_125;
  wire [63:0]        regroupV0_hi_hi_hi_hi_hi_hi_lo_5;
  assign regroupV0_hi_hi_hi_hi_hi_hi_lo_5 = _GEN_125;
  wire [63:0]        regroupV0_hi_hi_hi_hi_hi_hi_lo_10;
  assign regroupV0_hi_hi_hi_hi_hi_hi_lo_10 = _GEN_125;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_hi_hi_hi_hi_lo;
  assign slideAddressGen_slideMaskInput_hi_hi_hi_hi_hi_hi_lo = _GEN_125;
  wire [63:0]        selectReadStageMask_hi_hi_hi_hi_hi_hi_lo;
  assign selectReadStageMask_hi_hi_hi_hi_hi_hi_lo = _GEN_125;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_hi_hi_lo;
  assign maskSplit_maskSelect_hi_hi_hi_hi_hi_hi_lo = _GEN_125;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_hi_hi_lo_1;
  assign maskSplit_maskSelect_hi_hi_hi_hi_hi_hi_lo_1 = _GEN_125;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_hi_hi_lo_2;
  assign maskSplit_maskSelect_hi_hi_hi_hi_hi_hi_lo_2 = _GEN_125;
  wire [63:0]        maskForDestination_hi_hi_hi_hi_hi_hi_lo;
  assign maskForDestination_hi_hi_hi_hi_hi_hi_lo = _GEN_125;
  wire [63:0]        _GEN_126 = {v0_255, v0_254};
  wire [63:0]        regroupV0_hi_hi_hi_hi_hi_hi_hi;
  assign regroupV0_hi_hi_hi_hi_hi_hi_hi = _GEN_126;
  wire [63:0]        regroupV0_hi_hi_hi_hi_hi_hi_hi_5;
  assign regroupV0_hi_hi_hi_hi_hi_hi_hi_5 = _GEN_126;
  wire [63:0]        regroupV0_hi_hi_hi_hi_hi_hi_hi_10;
  assign regroupV0_hi_hi_hi_hi_hi_hi_hi_10 = _GEN_126;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_hi_hi_hi_hi_hi;
  assign slideAddressGen_slideMaskInput_hi_hi_hi_hi_hi_hi_hi = _GEN_126;
  wire [63:0]        selectReadStageMask_hi_hi_hi_hi_hi_hi_hi;
  assign selectReadStageMask_hi_hi_hi_hi_hi_hi_hi = _GEN_126;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_hi_hi_hi;
  assign maskSplit_maskSelect_hi_hi_hi_hi_hi_hi_hi = _GEN_126;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_hi_hi_hi_1;
  assign maskSplit_maskSelect_hi_hi_hi_hi_hi_hi_hi_1 = _GEN_126;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_hi_hi_hi_2;
  assign maskSplit_maskSelect_hi_hi_hi_hi_hi_hi_hi_2 = _GEN_126;
  wire [63:0]        maskForDestination_hi_hi_hi_hi_hi_hi_hi;
  assign maskForDestination_hi_hi_hi_hi_hi_hi_hi = _GEN_126;
  wire [127:0]       regroupV0_hi_hi_hi_hi_hi_hi = {regroupV0_hi_hi_hi_hi_hi_hi_hi, regroupV0_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]       regroupV0_hi_hi_hi_hi_hi = {regroupV0_hi_hi_hi_hi_hi_hi, regroupV0_hi_hi_hi_hi_hi_lo};
  wire [511:0]       regroupV0_hi_hi_hi_hi = {regroupV0_hi_hi_hi_hi_hi, regroupV0_hi_hi_hi_hi_lo};
  wire [1023:0]      regroupV0_hi_hi_hi = {regroupV0_hi_hi_hi_hi, regroupV0_hi_hi_hi_lo};
  wire [2047:0]      regroupV0_hi_hi = {regroupV0_hi_hi_hi, regroupV0_hi_hi_lo};
  wire [4095:0]      regroupV0_hi = {regroupV0_hi_hi, regroupV0_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo = {regroupV0_lo[19:16], regroupV0_lo[3:0]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi = {regroupV0_lo[51:48], regroupV0_lo[35:32]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_lo_lo_1 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo = {regroupV0_lo[83:80], regroupV0_lo[67:64]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi = {regroupV0_lo[115:112], regroupV0_lo[99:96]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_lo_hi_1 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [31:0]        regroupV0_lo_lo_lo_lo_lo_lo_1 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo = {regroupV0_lo[147:144], regroupV0_lo[131:128]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi = {regroupV0_lo[179:176], regroupV0_lo[163:160]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_hi_lo_1 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo = {regroupV0_lo[211:208], regroupV0_lo[195:192]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi = {regroupV0_lo[243:240], regroupV0_lo[227:224]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_hi_hi_1 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [31:0]        regroupV0_lo_lo_lo_lo_lo_hi_1 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_1, regroupV0_lo_lo_lo_lo_lo_hi_lo_1};
  wire [63:0]        regroupV0_lo_lo_lo_lo_lo_1 = {regroupV0_lo_lo_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo = {regroupV0_lo[275:272], regroupV0_lo[259:256]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi = {regroupV0_lo[307:304], regroupV0_lo[291:288]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_lo_lo_1 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo = {regroupV0_lo[339:336], regroupV0_lo[323:320]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi = {regroupV0_lo[371:368], regroupV0_lo[355:352]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_lo_hi_1 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [31:0]        regroupV0_lo_lo_lo_lo_hi_lo_1 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_1, regroupV0_lo_lo_lo_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo = {regroupV0_lo[403:400], regroupV0_lo[387:384]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi = {regroupV0_lo[435:432], regroupV0_lo[419:416]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_hi_lo_1 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo = {regroupV0_lo[467:464], regroupV0_lo[451:448]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi = {regroupV0_lo[499:496], regroupV0_lo[483:480]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_hi_hi_1 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [31:0]        regroupV0_lo_lo_lo_lo_hi_hi_1 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_1, regroupV0_lo_lo_lo_lo_hi_hi_lo_1};
  wire [63:0]        regroupV0_lo_lo_lo_lo_hi_1 = {regroupV0_lo_lo_lo_lo_hi_hi_1, regroupV0_lo_lo_lo_lo_hi_lo_1};
  wire [127:0]       regroupV0_lo_lo_lo_lo_1 = {regroupV0_lo_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo = {regroupV0_lo[531:528], regroupV0_lo[515:512]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi = {regroupV0_lo[563:560], regroupV0_lo[547:544]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_lo_lo_1 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo = {regroupV0_lo[595:592], regroupV0_lo[579:576]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi = {regroupV0_lo[627:624], regroupV0_lo[611:608]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_lo_hi_1 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [31:0]        regroupV0_lo_lo_lo_hi_lo_lo_1 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_1, regroupV0_lo_lo_lo_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo = {regroupV0_lo[659:656], regroupV0_lo[643:640]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi = {regroupV0_lo[691:688], regroupV0_lo[675:672]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_hi_lo_1 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo = {regroupV0_lo[723:720], regroupV0_lo[707:704]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi = {regroupV0_lo[755:752], regroupV0_lo[739:736]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_hi_hi_1 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [31:0]        regroupV0_lo_lo_lo_hi_lo_hi_1 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_1, regroupV0_lo_lo_lo_hi_lo_hi_lo_1};
  wire [63:0]        regroupV0_lo_lo_lo_hi_lo_1 = {regroupV0_lo_lo_lo_hi_lo_hi_1, regroupV0_lo_lo_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo = {regroupV0_lo[787:784], regroupV0_lo[771:768]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi = {regroupV0_lo[819:816], regroupV0_lo[803:800]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_lo_lo_1 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo = {regroupV0_lo[851:848], regroupV0_lo[835:832]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi = {regroupV0_lo[883:880], regroupV0_lo[867:864]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_lo_hi_1 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [31:0]        regroupV0_lo_lo_lo_hi_hi_lo_1 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_1, regroupV0_lo_lo_lo_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo = {regroupV0_lo[915:912], regroupV0_lo[899:896]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi = {regroupV0_lo[947:944], regroupV0_lo[931:928]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_hi_lo_1 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo = {regroupV0_lo[979:976], regroupV0_lo[963:960]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi = {regroupV0_lo[1011:1008], regroupV0_lo[995:992]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_hi_hi_1 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [31:0]        regroupV0_lo_lo_lo_hi_hi_hi_1 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_1, regroupV0_lo_lo_lo_hi_hi_hi_lo_1};
  wire [63:0]        regroupV0_lo_lo_lo_hi_hi_1 = {regroupV0_lo_lo_lo_hi_hi_hi_1, regroupV0_lo_lo_lo_hi_hi_lo_1};
  wire [127:0]       regroupV0_lo_lo_lo_hi_1 = {regroupV0_lo_lo_lo_hi_hi_1, regroupV0_lo_lo_lo_hi_lo_1};
  wire [255:0]       regroupV0_lo_lo_lo_1 = {regroupV0_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo = {regroupV0_lo[1043:1040], regroupV0_lo[1027:1024]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi = {regroupV0_lo[1075:1072], regroupV0_lo[1059:1056]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_lo_lo_1 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo = {regroupV0_lo[1107:1104], regroupV0_lo[1091:1088]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi = {regroupV0_lo[1139:1136], regroupV0_lo[1123:1120]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_lo_hi_1 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [31:0]        regroupV0_lo_lo_hi_lo_lo_lo_1 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_1, regroupV0_lo_lo_hi_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo = {regroupV0_lo[1171:1168], regroupV0_lo[1155:1152]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi = {regroupV0_lo[1203:1200], regroupV0_lo[1187:1184]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_hi_lo_1 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo = {regroupV0_lo[1235:1232], regroupV0_lo[1219:1216]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi = {regroupV0_lo[1267:1264], regroupV0_lo[1251:1248]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_hi_hi_1 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [31:0]        regroupV0_lo_lo_hi_lo_lo_hi_1 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_1, regroupV0_lo_lo_hi_lo_lo_hi_lo_1};
  wire [63:0]        regroupV0_lo_lo_hi_lo_lo_1 = {regroupV0_lo_lo_hi_lo_lo_hi_1, regroupV0_lo_lo_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo = {regroupV0_lo[1299:1296], regroupV0_lo[1283:1280]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi = {regroupV0_lo[1331:1328], regroupV0_lo[1315:1312]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_lo_lo_1 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo = {regroupV0_lo[1363:1360], regroupV0_lo[1347:1344]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi = {regroupV0_lo[1395:1392], regroupV0_lo[1379:1376]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_lo_hi_1 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [31:0]        regroupV0_lo_lo_hi_lo_hi_lo_1 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_1, regroupV0_lo_lo_hi_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo = {regroupV0_lo[1427:1424], regroupV0_lo[1411:1408]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi = {regroupV0_lo[1459:1456], regroupV0_lo[1443:1440]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_hi_lo_1 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo = {regroupV0_lo[1491:1488], regroupV0_lo[1475:1472]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi = {regroupV0_lo[1523:1520], regroupV0_lo[1507:1504]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_hi_hi_1 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [31:0]        regroupV0_lo_lo_hi_lo_hi_hi_1 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_1, regroupV0_lo_lo_hi_lo_hi_hi_lo_1};
  wire [63:0]        regroupV0_lo_lo_hi_lo_hi_1 = {regroupV0_lo_lo_hi_lo_hi_hi_1, regroupV0_lo_lo_hi_lo_hi_lo_1};
  wire [127:0]       regroupV0_lo_lo_hi_lo_1 = {regroupV0_lo_lo_hi_lo_hi_1, regroupV0_lo_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo = {regroupV0_lo[1555:1552], regroupV0_lo[1539:1536]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi = {regroupV0_lo[1587:1584], regroupV0_lo[1571:1568]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_lo_lo_1 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo = {regroupV0_lo[1619:1616], regroupV0_lo[1603:1600]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi = {regroupV0_lo[1651:1648], regroupV0_lo[1635:1632]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_lo_hi_1 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [31:0]        regroupV0_lo_lo_hi_hi_lo_lo_1 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_1, regroupV0_lo_lo_hi_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo = {regroupV0_lo[1683:1680], regroupV0_lo[1667:1664]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi = {regroupV0_lo[1715:1712], regroupV0_lo[1699:1696]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_hi_lo_1 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo = {regroupV0_lo[1747:1744], regroupV0_lo[1731:1728]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi = {regroupV0_lo[1779:1776], regroupV0_lo[1763:1760]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_hi_hi_1 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [31:0]        regroupV0_lo_lo_hi_hi_lo_hi_1 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_1, regroupV0_lo_lo_hi_hi_lo_hi_lo_1};
  wire [63:0]        regroupV0_lo_lo_hi_hi_lo_1 = {regroupV0_lo_lo_hi_hi_lo_hi_1, regroupV0_lo_lo_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo = {regroupV0_lo[1811:1808], regroupV0_lo[1795:1792]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi = {regroupV0_lo[1843:1840], regroupV0_lo[1827:1824]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_lo_lo_1 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo = {regroupV0_lo[1875:1872], regroupV0_lo[1859:1856]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi = {regroupV0_lo[1907:1904], regroupV0_lo[1891:1888]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_lo_hi_1 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [31:0]        regroupV0_lo_lo_hi_hi_hi_lo_1 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_1, regroupV0_lo_lo_hi_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo = {regroupV0_lo[1939:1936], regroupV0_lo[1923:1920]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi = {regroupV0_lo[1971:1968], regroupV0_lo[1955:1952]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_hi_lo_1 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo = {regroupV0_lo[2003:2000], regroupV0_lo[1987:1984]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi = {regroupV0_lo[2035:2032], regroupV0_lo[2019:2016]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_hi_hi_1 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [31:0]        regroupV0_lo_lo_hi_hi_hi_hi_1 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_1, regroupV0_lo_lo_hi_hi_hi_hi_lo_1};
  wire [63:0]        regroupV0_lo_lo_hi_hi_hi_1 = {regroupV0_lo_lo_hi_hi_hi_hi_1, regroupV0_lo_lo_hi_hi_hi_lo_1};
  wire [127:0]       regroupV0_lo_lo_hi_hi_1 = {regroupV0_lo_lo_hi_hi_hi_1, regroupV0_lo_lo_hi_hi_lo_1};
  wire [255:0]       regroupV0_lo_lo_hi_1 = {regroupV0_lo_lo_hi_hi_1, regroupV0_lo_lo_hi_lo_1};
  wire [511:0]       regroupV0_lo_lo_1 = {regroupV0_lo_lo_hi_1, regroupV0_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo = {regroupV0_lo[2067:2064], regroupV0_lo[2051:2048]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi = {regroupV0_lo[2099:2096], regroupV0_lo[2083:2080]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_lo_lo_1 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo = {regroupV0_lo[2131:2128], regroupV0_lo[2115:2112]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi = {regroupV0_lo[2163:2160], regroupV0_lo[2147:2144]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_lo_hi_1 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [31:0]        regroupV0_lo_hi_lo_lo_lo_lo_1 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_1, regroupV0_lo_hi_lo_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo = {regroupV0_lo[2195:2192], regroupV0_lo[2179:2176]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi = {regroupV0_lo[2227:2224], regroupV0_lo[2211:2208]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_hi_lo_1 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo = {regroupV0_lo[2259:2256], regroupV0_lo[2243:2240]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi = {regroupV0_lo[2291:2288], regroupV0_lo[2275:2272]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_hi_hi_1 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [31:0]        regroupV0_lo_hi_lo_lo_lo_hi_1 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_1, regroupV0_lo_hi_lo_lo_lo_hi_lo_1};
  wire [63:0]        regroupV0_lo_hi_lo_lo_lo_1 = {regroupV0_lo_hi_lo_lo_lo_hi_1, regroupV0_lo_hi_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo = {regroupV0_lo[2323:2320], regroupV0_lo[2307:2304]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi = {regroupV0_lo[2355:2352], regroupV0_lo[2339:2336]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_lo_lo_1 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo = {regroupV0_lo[2387:2384], regroupV0_lo[2371:2368]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi = {regroupV0_lo[2419:2416], regroupV0_lo[2403:2400]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_lo_hi_1 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [31:0]        regroupV0_lo_hi_lo_lo_hi_lo_1 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_1, regroupV0_lo_hi_lo_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo = {regroupV0_lo[2451:2448], regroupV0_lo[2435:2432]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi = {regroupV0_lo[2483:2480], regroupV0_lo[2467:2464]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_hi_lo_1 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo = {regroupV0_lo[2515:2512], regroupV0_lo[2499:2496]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi = {regroupV0_lo[2547:2544], regroupV0_lo[2531:2528]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_hi_hi_1 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [31:0]        regroupV0_lo_hi_lo_lo_hi_hi_1 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_1, regroupV0_lo_hi_lo_lo_hi_hi_lo_1};
  wire [63:0]        regroupV0_lo_hi_lo_lo_hi_1 = {regroupV0_lo_hi_lo_lo_hi_hi_1, regroupV0_lo_hi_lo_lo_hi_lo_1};
  wire [127:0]       regroupV0_lo_hi_lo_lo_1 = {regroupV0_lo_hi_lo_lo_hi_1, regroupV0_lo_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo = {regroupV0_lo[2579:2576], regroupV0_lo[2563:2560]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi = {regroupV0_lo[2611:2608], regroupV0_lo[2595:2592]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_lo_lo_1 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo = {regroupV0_lo[2643:2640], regroupV0_lo[2627:2624]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi = {regroupV0_lo[2675:2672], regroupV0_lo[2659:2656]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_lo_hi_1 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [31:0]        regroupV0_lo_hi_lo_hi_lo_lo_1 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_1, regroupV0_lo_hi_lo_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo = {regroupV0_lo[2707:2704], regroupV0_lo[2691:2688]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi = {regroupV0_lo[2739:2736], regroupV0_lo[2723:2720]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_hi_lo_1 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo = {regroupV0_lo[2771:2768], regroupV0_lo[2755:2752]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi = {regroupV0_lo[2803:2800], regroupV0_lo[2787:2784]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_hi_hi_1 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [31:0]        regroupV0_lo_hi_lo_hi_lo_hi_1 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_1, regroupV0_lo_hi_lo_hi_lo_hi_lo_1};
  wire [63:0]        regroupV0_lo_hi_lo_hi_lo_1 = {regroupV0_lo_hi_lo_hi_lo_hi_1, regroupV0_lo_hi_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo = {regroupV0_lo[2835:2832], regroupV0_lo[2819:2816]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi = {regroupV0_lo[2867:2864], regroupV0_lo[2851:2848]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_lo_lo_1 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo = {regroupV0_lo[2899:2896], regroupV0_lo[2883:2880]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi = {regroupV0_lo[2931:2928], regroupV0_lo[2915:2912]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_lo_hi_1 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [31:0]        regroupV0_lo_hi_lo_hi_hi_lo_1 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_1, regroupV0_lo_hi_lo_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo = {regroupV0_lo[2963:2960], regroupV0_lo[2947:2944]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi = {regroupV0_lo[2995:2992], regroupV0_lo[2979:2976]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_hi_lo_1 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo = {regroupV0_lo[3027:3024], regroupV0_lo[3011:3008]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi = {regroupV0_lo[3059:3056], regroupV0_lo[3043:3040]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_hi_hi_1 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [31:0]        regroupV0_lo_hi_lo_hi_hi_hi_1 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_1, regroupV0_lo_hi_lo_hi_hi_hi_lo_1};
  wire [63:0]        regroupV0_lo_hi_lo_hi_hi_1 = {regroupV0_lo_hi_lo_hi_hi_hi_1, regroupV0_lo_hi_lo_hi_hi_lo_1};
  wire [127:0]       regroupV0_lo_hi_lo_hi_1 = {regroupV0_lo_hi_lo_hi_hi_1, regroupV0_lo_hi_lo_hi_lo_1};
  wire [255:0]       regroupV0_lo_hi_lo_1 = {regroupV0_lo_hi_lo_hi_1, regroupV0_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo = {regroupV0_lo[3091:3088], regroupV0_lo[3075:3072]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi = {regroupV0_lo[3123:3120], regroupV0_lo[3107:3104]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_lo_lo_1 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo = {regroupV0_lo[3155:3152], regroupV0_lo[3139:3136]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi = {regroupV0_lo[3187:3184], regroupV0_lo[3171:3168]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_lo_hi_1 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [31:0]        regroupV0_lo_hi_hi_lo_lo_lo_1 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_1, regroupV0_lo_hi_hi_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo = {regroupV0_lo[3219:3216], regroupV0_lo[3203:3200]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi = {regroupV0_lo[3251:3248], regroupV0_lo[3235:3232]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_hi_lo_1 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo = {regroupV0_lo[3283:3280], regroupV0_lo[3267:3264]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi = {regroupV0_lo[3315:3312], regroupV0_lo[3299:3296]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_hi_hi_1 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [31:0]        regroupV0_lo_hi_hi_lo_lo_hi_1 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_1, regroupV0_lo_hi_hi_lo_lo_hi_lo_1};
  wire [63:0]        regroupV0_lo_hi_hi_lo_lo_1 = {regroupV0_lo_hi_hi_lo_lo_hi_1, regroupV0_lo_hi_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo = {regroupV0_lo[3347:3344], regroupV0_lo[3331:3328]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi = {regroupV0_lo[3379:3376], regroupV0_lo[3363:3360]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_lo_lo_1 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo = {regroupV0_lo[3411:3408], regroupV0_lo[3395:3392]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi = {regroupV0_lo[3443:3440], regroupV0_lo[3427:3424]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_lo_hi_1 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [31:0]        regroupV0_lo_hi_hi_lo_hi_lo_1 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_1, regroupV0_lo_hi_hi_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo = {regroupV0_lo[3475:3472], regroupV0_lo[3459:3456]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi = {regroupV0_lo[3507:3504], regroupV0_lo[3491:3488]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_hi_lo_1 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo = {regroupV0_lo[3539:3536], regroupV0_lo[3523:3520]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi = {regroupV0_lo[3571:3568], regroupV0_lo[3555:3552]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_hi_hi_1 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [31:0]        regroupV0_lo_hi_hi_lo_hi_hi_1 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_1, regroupV0_lo_hi_hi_lo_hi_hi_lo_1};
  wire [63:0]        regroupV0_lo_hi_hi_lo_hi_1 = {regroupV0_lo_hi_hi_lo_hi_hi_1, regroupV0_lo_hi_hi_lo_hi_lo_1};
  wire [127:0]       regroupV0_lo_hi_hi_lo_1 = {regroupV0_lo_hi_hi_lo_hi_1, regroupV0_lo_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo = {regroupV0_lo[3603:3600], regroupV0_lo[3587:3584]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi = {regroupV0_lo[3635:3632], regroupV0_lo[3619:3616]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_lo_lo_1 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo = {regroupV0_lo[3667:3664], regroupV0_lo[3651:3648]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi = {regroupV0_lo[3699:3696], regroupV0_lo[3683:3680]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_lo_hi_1 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [31:0]        regroupV0_lo_hi_hi_hi_lo_lo_1 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_1, regroupV0_lo_hi_hi_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo = {regroupV0_lo[3731:3728], regroupV0_lo[3715:3712]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi = {regroupV0_lo[3763:3760], regroupV0_lo[3747:3744]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_hi_lo_1 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo = {regroupV0_lo[3795:3792], regroupV0_lo[3779:3776]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi = {regroupV0_lo[3827:3824], regroupV0_lo[3811:3808]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_hi_hi_1 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [31:0]        regroupV0_lo_hi_hi_hi_lo_hi_1 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_1, regroupV0_lo_hi_hi_hi_lo_hi_lo_1};
  wire [63:0]        regroupV0_lo_hi_hi_hi_lo_1 = {regroupV0_lo_hi_hi_hi_lo_hi_1, regroupV0_lo_hi_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo = {regroupV0_lo[3859:3856], regroupV0_lo[3843:3840]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi = {regroupV0_lo[3891:3888], regroupV0_lo[3875:3872]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_lo_lo_1 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo = {regroupV0_lo[3923:3920], regroupV0_lo[3907:3904]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi = {regroupV0_lo[3955:3952], regroupV0_lo[3939:3936]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_lo_hi_1 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [31:0]        regroupV0_lo_hi_hi_hi_hi_lo_1 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_1, regroupV0_lo_hi_hi_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo = {regroupV0_lo[3987:3984], regroupV0_lo[3971:3968]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi = {regroupV0_lo[4019:4016], regroupV0_lo[4003:4000]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_hi_lo_1 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo = {regroupV0_lo[4051:4048], regroupV0_lo[4035:4032]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi = {regroupV0_lo[4083:4080], regroupV0_lo[4067:4064]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_hi_hi_1 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [31:0]        regroupV0_lo_hi_hi_hi_hi_hi_1 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_1, regroupV0_lo_hi_hi_hi_hi_hi_lo_1};
  wire [63:0]        regroupV0_lo_hi_hi_hi_hi_1 = {regroupV0_lo_hi_hi_hi_hi_hi_1, regroupV0_lo_hi_hi_hi_hi_lo_1};
  wire [127:0]       regroupV0_lo_hi_hi_hi_1 = {regroupV0_lo_hi_hi_hi_hi_1, regroupV0_lo_hi_hi_hi_lo_1};
  wire [255:0]       regroupV0_lo_hi_hi_1 = {regroupV0_lo_hi_hi_hi_1, regroupV0_lo_hi_hi_lo_1};
  wire [511:0]       regroupV0_lo_hi_1 = {regroupV0_lo_hi_hi_1, regroupV0_lo_hi_lo_1};
  wire [1023:0]      regroupV0_lo_1 = {regroupV0_lo_hi_1, regroupV0_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo = {regroupV0_hi[19:16], regroupV0_hi[3:0]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi = {regroupV0_hi[51:48], regroupV0_hi[35:32]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_lo_lo_1 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo = {regroupV0_hi[83:80], regroupV0_hi[67:64]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi = {regroupV0_hi[115:112], regroupV0_hi[99:96]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_lo_hi_1 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [31:0]        regroupV0_hi_lo_lo_lo_lo_lo_1 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo = {regroupV0_hi[147:144], regroupV0_hi[131:128]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi = {regroupV0_hi[179:176], regroupV0_hi[163:160]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_hi_lo_1 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo = {regroupV0_hi[211:208], regroupV0_hi[195:192]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi = {regroupV0_hi[243:240], regroupV0_hi[227:224]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_hi_hi_1 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [31:0]        regroupV0_hi_lo_lo_lo_lo_hi_1 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_1, regroupV0_hi_lo_lo_lo_lo_hi_lo_1};
  wire [63:0]        regroupV0_hi_lo_lo_lo_lo_1 = {regroupV0_hi_lo_lo_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo = {regroupV0_hi[275:272], regroupV0_hi[259:256]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi = {regroupV0_hi[307:304], regroupV0_hi[291:288]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_lo_lo_1 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo = {regroupV0_hi[339:336], regroupV0_hi[323:320]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi = {regroupV0_hi[371:368], regroupV0_hi[355:352]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_lo_hi_1 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [31:0]        regroupV0_hi_lo_lo_lo_hi_lo_1 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_1, regroupV0_hi_lo_lo_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo = {regroupV0_hi[403:400], regroupV0_hi[387:384]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi = {regroupV0_hi[435:432], regroupV0_hi[419:416]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_hi_lo_1 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo = {regroupV0_hi[467:464], regroupV0_hi[451:448]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi = {regroupV0_hi[499:496], regroupV0_hi[483:480]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_hi_hi_1 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [31:0]        regroupV0_hi_lo_lo_lo_hi_hi_1 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_1, regroupV0_hi_lo_lo_lo_hi_hi_lo_1};
  wire [63:0]        regroupV0_hi_lo_lo_lo_hi_1 = {regroupV0_hi_lo_lo_lo_hi_hi_1, regroupV0_hi_lo_lo_lo_hi_lo_1};
  wire [127:0]       regroupV0_hi_lo_lo_lo_1 = {regroupV0_hi_lo_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo = {regroupV0_hi[531:528], regroupV0_hi[515:512]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi = {regroupV0_hi[563:560], regroupV0_hi[547:544]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_lo_lo_1 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo = {regroupV0_hi[595:592], regroupV0_hi[579:576]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi = {regroupV0_hi[627:624], regroupV0_hi[611:608]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_lo_hi_1 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [31:0]        regroupV0_hi_lo_lo_hi_lo_lo_1 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_1, regroupV0_hi_lo_lo_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo = {regroupV0_hi[659:656], regroupV0_hi[643:640]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi = {regroupV0_hi[691:688], regroupV0_hi[675:672]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_hi_lo_1 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo = {regroupV0_hi[723:720], regroupV0_hi[707:704]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi = {regroupV0_hi[755:752], regroupV0_hi[739:736]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_hi_hi_1 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [31:0]        regroupV0_hi_lo_lo_hi_lo_hi_1 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_1, regroupV0_hi_lo_lo_hi_lo_hi_lo_1};
  wire [63:0]        regroupV0_hi_lo_lo_hi_lo_1 = {regroupV0_hi_lo_lo_hi_lo_hi_1, regroupV0_hi_lo_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo = {regroupV0_hi[787:784], regroupV0_hi[771:768]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi = {regroupV0_hi[819:816], regroupV0_hi[803:800]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_lo_lo_1 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo = {regroupV0_hi[851:848], regroupV0_hi[835:832]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi = {regroupV0_hi[883:880], regroupV0_hi[867:864]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_lo_hi_1 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [31:0]        regroupV0_hi_lo_lo_hi_hi_lo_1 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_1, regroupV0_hi_lo_lo_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo = {regroupV0_hi[915:912], regroupV0_hi[899:896]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi = {regroupV0_hi[947:944], regroupV0_hi[931:928]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_hi_lo_1 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo = {regroupV0_hi[979:976], regroupV0_hi[963:960]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi = {regroupV0_hi[1011:1008], regroupV0_hi[995:992]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_hi_hi_1 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [31:0]        regroupV0_hi_lo_lo_hi_hi_hi_1 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_1, regroupV0_hi_lo_lo_hi_hi_hi_lo_1};
  wire [63:0]        regroupV0_hi_lo_lo_hi_hi_1 = {regroupV0_hi_lo_lo_hi_hi_hi_1, regroupV0_hi_lo_lo_hi_hi_lo_1};
  wire [127:0]       regroupV0_hi_lo_lo_hi_1 = {regroupV0_hi_lo_lo_hi_hi_1, regroupV0_hi_lo_lo_hi_lo_1};
  wire [255:0]       regroupV0_hi_lo_lo_1 = {regroupV0_hi_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo = {regroupV0_hi[1043:1040], regroupV0_hi[1027:1024]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi = {regroupV0_hi[1075:1072], regroupV0_hi[1059:1056]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_lo_lo_1 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo = {regroupV0_hi[1107:1104], regroupV0_hi[1091:1088]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi = {regroupV0_hi[1139:1136], regroupV0_hi[1123:1120]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_lo_hi_1 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [31:0]        regroupV0_hi_lo_hi_lo_lo_lo_1 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_1, regroupV0_hi_lo_hi_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo = {regroupV0_hi[1171:1168], regroupV0_hi[1155:1152]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi = {regroupV0_hi[1203:1200], regroupV0_hi[1187:1184]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_hi_lo_1 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo = {regroupV0_hi[1235:1232], regroupV0_hi[1219:1216]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi = {regroupV0_hi[1267:1264], regroupV0_hi[1251:1248]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_hi_hi_1 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [31:0]        regroupV0_hi_lo_hi_lo_lo_hi_1 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_1, regroupV0_hi_lo_hi_lo_lo_hi_lo_1};
  wire [63:0]        regroupV0_hi_lo_hi_lo_lo_1 = {regroupV0_hi_lo_hi_lo_lo_hi_1, regroupV0_hi_lo_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo = {regroupV0_hi[1299:1296], regroupV0_hi[1283:1280]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi = {regroupV0_hi[1331:1328], regroupV0_hi[1315:1312]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_lo_lo_1 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo = {regroupV0_hi[1363:1360], regroupV0_hi[1347:1344]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi = {regroupV0_hi[1395:1392], regroupV0_hi[1379:1376]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_lo_hi_1 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [31:0]        regroupV0_hi_lo_hi_lo_hi_lo_1 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_1, regroupV0_hi_lo_hi_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo = {regroupV0_hi[1427:1424], regroupV0_hi[1411:1408]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi = {regroupV0_hi[1459:1456], regroupV0_hi[1443:1440]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_hi_lo_1 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo = {regroupV0_hi[1491:1488], regroupV0_hi[1475:1472]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi = {regroupV0_hi[1523:1520], regroupV0_hi[1507:1504]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_hi_hi_1 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [31:0]        regroupV0_hi_lo_hi_lo_hi_hi_1 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_1, regroupV0_hi_lo_hi_lo_hi_hi_lo_1};
  wire [63:0]        regroupV0_hi_lo_hi_lo_hi_1 = {regroupV0_hi_lo_hi_lo_hi_hi_1, regroupV0_hi_lo_hi_lo_hi_lo_1};
  wire [127:0]       regroupV0_hi_lo_hi_lo_1 = {regroupV0_hi_lo_hi_lo_hi_1, regroupV0_hi_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo = {regroupV0_hi[1555:1552], regroupV0_hi[1539:1536]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi = {regroupV0_hi[1587:1584], regroupV0_hi[1571:1568]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_lo_lo_1 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo = {regroupV0_hi[1619:1616], regroupV0_hi[1603:1600]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi = {regroupV0_hi[1651:1648], regroupV0_hi[1635:1632]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_lo_hi_1 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [31:0]        regroupV0_hi_lo_hi_hi_lo_lo_1 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_1, regroupV0_hi_lo_hi_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo = {regroupV0_hi[1683:1680], regroupV0_hi[1667:1664]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi = {regroupV0_hi[1715:1712], regroupV0_hi[1699:1696]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_hi_lo_1 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo = {regroupV0_hi[1747:1744], regroupV0_hi[1731:1728]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi = {regroupV0_hi[1779:1776], regroupV0_hi[1763:1760]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_hi_hi_1 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [31:0]        regroupV0_hi_lo_hi_hi_lo_hi_1 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_1, regroupV0_hi_lo_hi_hi_lo_hi_lo_1};
  wire [63:0]        regroupV0_hi_lo_hi_hi_lo_1 = {regroupV0_hi_lo_hi_hi_lo_hi_1, regroupV0_hi_lo_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo = {regroupV0_hi[1811:1808], regroupV0_hi[1795:1792]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi = {regroupV0_hi[1843:1840], regroupV0_hi[1827:1824]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_lo_lo_1 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo = {regroupV0_hi[1875:1872], regroupV0_hi[1859:1856]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi = {regroupV0_hi[1907:1904], regroupV0_hi[1891:1888]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_lo_hi_1 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [31:0]        regroupV0_hi_lo_hi_hi_hi_lo_1 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_1, regroupV0_hi_lo_hi_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo = {regroupV0_hi[1939:1936], regroupV0_hi[1923:1920]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi = {regroupV0_hi[1971:1968], regroupV0_hi[1955:1952]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_hi_lo_1 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo = {regroupV0_hi[2003:2000], regroupV0_hi[1987:1984]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi = {regroupV0_hi[2035:2032], regroupV0_hi[2019:2016]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_hi_hi_1 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [31:0]        regroupV0_hi_lo_hi_hi_hi_hi_1 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_1, regroupV0_hi_lo_hi_hi_hi_hi_lo_1};
  wire [63:0]        regroupV0_hi_lo_hi_hi_hi_1 = {regroupV0_hi_lo_hi_hi_hi_hi_1, regroupV0_hi_lo_hi_hi_hi_lo_1};
  wire [127:0]       regroupV0_hi_lo_hi_hi_1 = {regroupV0_hi_lo_hi_hi_hi_1, regroupV0_hi_lo_hi_hi_lo_1};
  wire [255:0]       regroupV0_hi_lo_hi_1 = {regroupV0_hi_lo_hi_hi_1, regroupV0_hi_lo_hi_lo_1};
  wire [511:0]       regroupV0_hi_lo_1 = {regroupV0_hi_lo_hi_1, regroupV0_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo = {regroupV0_hi[2067:2064], regroupV0_hi[2051:2048]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi = {regroupV0_hi[2099:2096], regroupV0_hi[2083:2080]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_lo_lo_1 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo = {regroupV0_hi[2131:2128], regroupV0_hi[2115:2112]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi = {regroupV0_hi[2163:2160], regroupV0_hi[2147:2144]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_lo_hi_1 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [31:0]        regroupV0_hi_hi_lo_lo_lo_lo_1 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_1, regroupV0_hi_hi_lo_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo = {regroupV0_hi[2195:2192], regroupV0_hi[2179:2176]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi = {regroupV0_hi[2227:2224], regroupV0_hi[2211:2208]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_hi_lo_1 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo = {regroupV0_hi[2259:2256], regroupV0_hi[2243:2240]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi = {regroupV0_hi[2291:2288], regroupV0_hi[2275:2272]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_hi_hi_1 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [31:0]        regroupV0_hi_hi_lo_lo_lo_hi_1 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_1, regroupV0_hi_hi_lo_lo_lo_hi_lo_1};
  wire [63:0]        regroupV0_hi_hi_lo_lo_lo_1 = {regroupV0_hi_hi_lo_lo_lo_hi_1, regroupV0_hi_hi_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo = {regroupV0_hi[2323:2320], regroupV0_hi[2307:2304]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi = {regroupV0_hi[2355:2352], regroupV0_hi[2339:2336]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_lo_lo_1 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo = {regroupV0_hi[2387:2384], regroupV0_hi[2371:2368]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi = {regroupV0_hi[2419:2416], regroupV0_hi[2403:2400]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_lo_hi_1 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [31:0]        regroupV0_hi_hi_lo_lo_hi_lo_1 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_1, regroupV0_hi_hi_lo_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo = {regroupV0_hi[2451:2448], regroupV0_hi[2435:2432]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi = {regroupV0_hi[2483:2480], regroupV0_hi[2467:2464]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_hi_lo_1 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo = {regroupV0_hi[2515:2512], regroupV0_hi[2499:2496]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi = {regroupV0_hi[2547:2544], regroupV0_hi[2531:2528]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_hi_hi_1 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [31:0]        regroupV0_hi_hi_lo_lo_hi_hi_1 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_1, regroupV0_hi_hi_lo_lo_hi_hi_lo_1};
  wire [63:0]        regroupV0_hi_hi_lo_lo_hi_1 = {regroupV0_hi_hi_lo_lo_hi_hi_1, regroupV0_hi_hi_lo_lo_hi_lo_1};
  wire [127:0]       regroupV0_hi_hi_lo_lo_1 = {regroupV0_hi_hi_lo_lo_hi_1, regroupV0_hi_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo = {regroupV0_hi[2579:2576], regroupV0_hi[2563:2560]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi = {regroupV0_hi[2611:2608], regroupV0_hi[2595:2592]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_lo_lo_1 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo = {regroupV0_hi[2643:2640], regroupV0_hi[2627:2624]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi = {regroupV0_hi[2675:2672], regroupV0_hi[2659:2656]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_lo_hi_1 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [31:0]        regroupV0_hi_hi_lo_hi_lo_lo_1 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_1, regroupV0_hi_hi_lo_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo = {regroupV0_hi[2707:2704], regroupV0_hi[2691:2688]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi = {regroupV0_hi[2739:2736], regroupV0_hi[2723:2720]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_hi_lo_1 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo = {regroupV0_hi[2771:2768], regroupV0_hi[2755:2752]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi = {regroupV0_hi[2803:2800], regroupV0_hi[2787:2784]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_hi_hi_1 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [31:0]        regroupV0_hi_hi_lo_hi_lo_hi_1 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_1, regroupV0_hi_hi_lo_hi_lo_hi_lo_1};
  wire [63:0]        regroupV0_hi_hi_lo_hi_lo_1 = {regroupV0_hi_hi_lo_hi_lo_hi_1, regroupV0_hi_hi_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo = {regroupV0_hi[2835:2832], regroupV0_hi[2819:2816]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi = {regroupV0_hi[2867:2864], regroupV0_hi[2851:2848]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_lo_lo_1 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo = {regroupV0_hi[2899:2896], regroupV0_hi[2883:2880]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi = {regroupV0_hi[2931:2928], regroupV0_hi[2915:2912]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_lo_hi_1 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [31:0]        regroupV0_hi_hi_lo_hi_hi_lo_1 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_1, regroupV0_hi_hi_lo_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo = {regroupV0_hi[2963:2960], regroupV0_hi[2947:2944]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi = {regroupV0_hi[2995:2992], regroupV0_hi[2979:2976]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_hi_lo_1 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo = {regroupV0_hi[3027:3024], regroupV0_hi[3011:3008]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi = {regroupV0_hi[3059:3056], regroupV0_hi[3043:3040]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_hi_hi_1 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [31:0]        regroupV0_hi_hi_lo_hi_hi_hi_1 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_1, regroupV0_hi_hi_lo_hi_hi_hi_lo_1};
  wire [63:0]        regroupV0_hi_hi_lo_hi_hi_1 = {regroupV0_hi_hi_lo_hi_hi_hi_1, regroupV0_hi_hi_lo_hi_hi_lo_1};
  wire [127:0]       regroupV0_hi_hi_lo_hi_1 = {regroupV0_hi_hi_lo_hi_hi_1, regroupV0_hi_hi_lo_hi_lo_1};
  wire [255:0]       regroupV0_hi_hi_lo_1 = {regroupV0_hi_hi_lo_hi_1, regroupV0_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo = {regroupV0_hi[3091:3088], regroupV0_hi[3075:3072]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi = {regroupV0_hi[3123:3120], regroupV0_hi[3107:3104]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_lo_lo_1 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo = {regroupV0_hi[3155:3152], regroupV0_hi[3139:3136]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi = {regroupV0_hi[3187:3184], regroupV0_hi[3171:3168]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_lo_hi_1 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [31:0]        regroupV0_hi_hi_hi_lo_lo_lo_1 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_1, regroupV0_hi_hi_hi_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo = {regroupV0_hi[3219:3216], regroupV0_hi[3203:3200]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi = {regroupV0_hi[3251:3248], regroupV0_hi[3235:3232]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_hi_lo_1 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo = {regroupV0_hi[3283:3280], regroupV0_hi[3267:3264]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi = {regroupV0_hi[3315:3312], regroupV0_hi[3299:3296]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_hi_hi_1 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [31:0]        regroupV0_hi_hi_hi_lo_lo_hi_1 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_1, regroupV0_hi_hi_hi_lo_lo_hi_lo_1};
  wire [63:0]        regroupV0_hi_hi_hi_lo_lo_1 = {regroupV0_hi_hi_hi_lo_lo_hi_1, regroupV0_hi_hi_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo = {regroupV0_hi[3347:3344], regroupV0_hi[3331:3328]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi = {regroupV0_hi[3379:3376], regroupV0_hi[3363:3360]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_lo_lo_1 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo = {regroupV0_hi[3411:3408], regroupV0_hi[3395:3392]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi = {regroupV0_hi[3443:3440], regroupV0_hi[3427:3424]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_lo_hi_1 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [31:0]        regroupV0_hi_hi_hi_lo_hi_lo_1 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_1, regroupV0_hi_hi_hi_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo = {regroupV0_hi[3475:3472], regroupV0_hi[3459:3456]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi = {regroupV0_hi[3507:3504], regroupV0_hi[3491:3488]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_hi_lo_1 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo = {regroupV0_hi[3539:3536], regroupV0_hi[3523:3520]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi = {regroupV0_hi[3571:3568], regroupV0_hi[3555:3552]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_hi_hi_1 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [31:0]        regroupV0_hi_hi_hi_lo_hi_hi_1 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_1, regroupV0_hi_hi_hi_lo_hi_hi_lo_1};
  wire [63:0]        regroupV0_hi_hi_hi_lo_hi_1 = {regroupV0_hi_hi_hi_lo_hi_hi_1, regroupV0_hi_hi_hi_lo_hi_lo_1};
  wire [127:0]       regroupV0_hi_hi_hi_lo_1 = {regroupV0_hi_hi_hi_lo_hi_1, regroupV0_hi_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo = {regroupV0_hi[3603:3600], regroupV0_hi[3587:3584]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi = {regroupV0_hi[3635:3632], regroupV0_hi[3619:3616]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_lo_lo_1 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo = {regroupV0_hi[3667:3664], regroupV0_hi[3651:3648]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi = {regroupV0_hi[3699:3696], regroupV0_hi[3683:3680]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_lo_hi_1 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [31:0]        regroupV0_hi_hi_hi_hi_lo_lo_1 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_1, regroupV0_hi_hi_hi_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo = {regroupV0_hi[3731:3728], regroupV0_hi[3715:3712]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi = {regroupV0_hi[3763:3760], regroupV0_hi[3747:3744]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_hi_lo_1 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo = {regroupV0_hi[3795:3792], regroupV0_hi[3779:3776]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi = {regroupV0_hi[3827:3824], regroupV0_hi[3811:3808]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_hi_hi_1 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [31:0]        regroupV0_hi_hi_hi_hi_lo_hi_1 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_1, regroupV0_hi_hi_hi_hi_lo_hi_lo_1};
  wire [63:0]        regroupV0_hi_hi_hi_hi_lo_1 = {regroupV0_hi_hi_hi_hi_lo_hi_1, regroupV0_hi_hi_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo = {regroupV0_hi[3859:3856], regroupV0_hi[3843:3840]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi = {regroupV0_hi[3891:3888], regroupV0_hi[3875:3872]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_lo_lo_1 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo = {regroupV0_hi[3923:3920], regroupV0_hi[3907:3904]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi = {regroupV0_hi[3955:3952], regroupV0_hi[3939:3936]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_lo_hi_1 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [31:0]        regroupV0_hi_hi_hi_hi_hi_lo_1 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_1, regroupV0_hi_hi_hi_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo = {regroupV0_hi[3987:3984], regroupV0_hi[3971:3968]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi = {regroupV0_hi[4019:4016], regroupV0_hi[4003:4000]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_hi_lo_1 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo = {regroupV0_hi[4051:4048], regroupV0_hi[4035:4032]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi = {regroupV0_hi[4083:4080], regroupV0_hi[4067:4064]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_hi_hi_1 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [31:0]        regroupV0_hi_hi_hi_hi_hi_hi_1 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_hi_hi_hi_lo_1};
  wire [63:0]        regroupV0_hi_hi_hi_hi_hi_1 = {regroupV0_hi_hi_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_hi_hi_lo_1};
  wire [127:0]       regroupV0_hi_hi_hi_hi_1 = {regroupV0_hi_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_hi_lo_1};
  wire [255:0]       regroupV0_hi_hi_hi_1 = {regroupV0_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_lo_1};
  wire [511:0]       regroupV0_hi_hi_1 = {regroupV0_hi_hi_hi_1, regroupV0_hi_hi_lo_1};
  wire [1023:0]      regroupV0_hi_1 = {regroupV0_hi_hi_1, regroupV0_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_1 = {regroupV0_lo[23:20], regroupV0_lo[7:4]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_1 = {regroupV0_lo[55:52], regroupV0_lo[39:36]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_lo_lo_2 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_1 = {regroupV0_lo[87:84], regroupV0_lo[71:68]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_1 = {regroupV0_lo[119:116], regroupV0_lo[103:100]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_lo_hi_2 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_1, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_1};
  wire [31:0]        regroupV0_lo_lo_lo_lo_lo_lo_2 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_1 = {regroupV0_lo[151:148], regroupV0_lo[135:132]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_1 = {regroupV0_lo[183:180], regroupV0_lo[167:164]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_hi_lo_2 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_1, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_1 = {regroupV0_lo[215:212], regroupV0_lo[199:196]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_1 = {regroupV0_lo[247:244], regroupV0_lo[231:228]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_hi_hi_2 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_1, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_1};
  wire [31:0]        regroupV0_lo_lo_lo_lo_lo_hi_2 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_2, regroupV0_lo_lo_lo_lo_lo_hi_lo_2};
  wire [63:0]        regroupV0_lo_lo_lo_lo_lo_2 = {regroupV0_lo_lo_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_1 = {regroupV0_lo[279:276], regroupV0_lo[263:260]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_1 = {regroupV0_lo[311:308], regroupV0_lo[295:292]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_lo_lo_2 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_1 = {regroupV0_lo[343:340], regroupV0_lo[327:324]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_1 = {regroupV0_lo[375:372], regroupV0_lo[359:356]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_lo_hi_2 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_1, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_1};
  wire [31:0]        regroupV0_lo_lo_lo_lo_hi_lo_2 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_2, regroupV0_lo_lo_lo_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_1 = {regroupV0_lo[407:404], regroupV0_lo[391:388]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_1 = {regroupV0_lo[439:436], regroupV0_lo[423:420]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_hi_lo_2 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_1, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_1 = {regroupV0_lo[471:468], regroupV0_lo[455:452]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_1 = {regroupV0_lo[503:500], regroupV0_lo[487:484]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_hi_hi_2 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_1, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_1};
  wire [31:0]        regroupV0_lo_lo_lo_lo_hi_hi_2 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_2, regroupV0_lo_lo_lo_lo_hi_hi_lo_2};
  wire [63:0]        regroupV0_lo_lo_lo_lo_hi_2 = {regroupV0_lo_lo_lo_lo_hi_hi_2, regroupV0_lo_lo_lo_lo_hi_lo_2};
  wire [127:0]       regroupV0_lo_lo_lo_lo_2 = {regroupV0_lo_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_1 = {regroupV0_lo[535:532], regroupV0_lo[519:516]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_1 = {regroupV0_lo[567:564], regroupV0_lo[551:548]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_lo_lo_2 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_1 = {regroupV0_lo[599:596], regroupV0_lo[583:580]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_1 = {regroupV0_lo[631:628], regroupV0_lo[615:612]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_lo_hi_2 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_1, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_1};
  wire [31:0]        regroupV0_lo_lo_lo_hi_lo_lo_2 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_2, regroupV0_lo_lo_lo_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_1 = {regroupV0_lo[663:660], regroupV0_lo[647:644]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_1 = {regroupV0_lo[695:692], regroupV0_lo[679:676]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_hi_lo_2 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_1, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_1 = {regroupV0_lo[727:724], regroupV0_lo[711:708]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_1 = {regroupV0_lo[759:756], regroupV0_lo[743:740]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_hi_hi_2 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_1, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_1};
  wire [31:0]        regroupV0_lo_lo_lo_hi_lo_hi_2 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_2, regroupV0_lo_lo_lo_hi_lo_hi_lo_2};
  wire [63:0]        regroupV0_lo_lo_lo_hi_lo_2 = {regroupV0_lo_lo_lo_hi_lo_hi_2, regroupV0_lo_lo_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_1 = {regroupV0_lo[791:788], regroupV0_lo[775:772]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_1 = {regroupV0_lo[823:820], regroupV0_lo[807:804]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_lo_lo_2 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_1, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_1 = {regroupV0_lo[855:852], regroupV0_lo[839:836]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_1 = {regroupV0_lo[887:884], regroupV0_lo[871:868]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_lo_hi_2 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_1, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_1};
  wire [31:0]        regroupV0_lo_lo_lo_hi_hi_lo_2 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_2, regroupV0_lo_lo_lo_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_1 = {regroupV0_lo[919:916], regroupV0_lo[903:900]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_1 = {regroupV0_lo[951:948], regroupV0_lo[935:932]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_hi_lo_2 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_1, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_1 = {regroupV0_lo[983:980], regroupV0_lo[967:964]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_1 = {regroupV0_lo[1015:1012], regroupV0_lo[999:996]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_hi_hi_2 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_1, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_1};
  wire [31:0]        regroupV0_lo_lo_lo_hi_hi_hi_2 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_2, regroupV0_lo_lo_lo_hi_hi_hi_lo_2};
  wire [63:0]        regroupV0_lo_lo_lo_hi_hi_2 = {regroupV0_lo_lo_lo_hi_hi_hi_2, regroupV0_lo_lo_lo_hi_hi_lo_2};
  wire [127:0]       regroupV0_lo_lo_lo_hi_2 = {regroupV0_lo_lo_lo_hi_hi_2, regroupV0_lo_lo_lo_hi_lo_2};
  wire [255:0]       regroupV0_lo_lo_lo_2 = {regroupV0_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_1 = {regroupV0_lo[1047:1044], regroupV0_lo[1031:1028]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_1 = {regroupV0_lo[1079:1076], regroupV0_lo[1063:1060]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_lo_lo_2 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_1, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_1 = {regroupV0_lo[1111:1108], regroupV0_lo[1095:1092]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_1 = {regroupV0_lo[1143:1140], regroupV0_lo[1127:1124]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_lo_hi_2 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_1, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_1};
  wire [31:0]        regroupV0_lo_lo_hi_lo_lo_lo_2 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_2, regroupV0_lo_lo_hi_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_1 = {regroupV0_lo[1175:1172], regroupV0_lo[1159:1156]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_1 = {regroupV0_lo[1207:1204], regroupV0_lo[1191:1188]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_hi_lo_2 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_1, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_1 = {regroupV0_lo[1239:1236], regroupV0_lo[1223:1220]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_1 = {regroupV0_lo[1271:1268], regroupV0_lo[1255:1252]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_hi_hi_2 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_1, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_1};
  wire [31:0]        regroupV0_lo_lo_hi_lo_lo_hi_2 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_2, regroupV0_lo_lo_hi_lo_lo_hi_lo_2};
  wire [63:0]        regroupV0_lo_lo_hi_lo_lo_2 = {regroupV0_lo_lo_hi_lo_lo_hi_2, regroupV0_lo_lo_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_1 = {regroupV0_lo[1303:1300], regroupV0_lo[1287:1284]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_1 = {regroupV0_lo[1335:1332], regroupV0_lo[1319:1316]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_lo_lo_2 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_1, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_1 = {regroupV0_lo[1367:1364], regroupV0_lo[1351:1348]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_1 = {regroupV0_lo[1399:1396], regroupV0_lo[1383:1380]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_lo_hi_2 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_1, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_1};
  wire [31:0]        regroupV0_lo_lo_hi_lo_hi_lo_2 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_2, regroupV0_lo_lo_hi_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_1 = {regroupV0_lo[1431:1428], regroupV0_lo[1415:1412]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_1 = {regroupV0_lo[1463:1460], regroupV0_lo[1447:1444]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_hi_lo_2 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_1, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_1 = {regroupV0_lo[1495:1492], regroupV0_lo[1479:1476]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_1 = {regroupV0_lo[1527:1524], regroupV0_lo[1511:1508]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_hi_hi_2 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_1, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_1};
  wire [31:0]        regroupV0_lo_lo_hi_lo_hi_hi_2 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_2, regroupV0_lo_lo_hi_lo_hi_hi_lo_2};
  wire [63:0]        regroupV0_lo_lo_hi_lo_hi_2 = {regroupV0_lo_lo_hi_lo_hi_hi_2, regroupV0_lo_lo_hi_lo_hi_lo_2};
  wire [127:0]       regroupV0_lo_lo_hi_lo_2 = {regroupV0_lo_lo_hi_lo_hi_2, regroupV0_lo_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_1 = {regroupV0_lo[1559:1556], regroupV0_lo[1543:1540]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_1 = {regroupV0_lo[1591:1588], regroupV0_lo[1575:1572]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_lo_lo_2 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_1, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_1 = {regroupV0_lo[1623:1620], regroupV0_lo[1607:1604]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_1 = {regroupV0_lo[1655:1652], regroupV0_lo[1639:1636]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_lo_hi_2 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_1, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_1};
  wire [31:0]        regroupV0_lo_lo_hi_hi_lo_lo_2 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_2, regroupV0_lo_lo_hi_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_1 = {regroupV0_lo[1687:1684], regroupV0_lo[1671:1668]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_1 = {regroupV0_lo[1719:1716], regroupV0_lo[1703:1700]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_hi_lo_2 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_1, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_1 = {regroupV0_lo[1751:1748], regroupV0_lo[1735:1732]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_1 = {regroupV0_lo[1783:1780], regroupV0_lo[1767:1764]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_hi_hi_2 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_1, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_1};
  wire [31:0]        regroupV0_lo_lo_hi_hi_lo_hi_2 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_2, regroupV0_lo_lo_hi_hi_lo_hi_lo_2};
  wire [63:0]        regroupV0_lo_lo_hi_hi_lo_2 = {regroupV0_lo_lo_hi_hi_lo_hi_2, regroupV0_lo_lo_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_1 = {regroupV0_lo[1815:1812], regroupV0_lo[1799:1796]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_1 = {regroupV0_lo[1847:1844], regroupV0_lo[1831:1828]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_lo_lo_2 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_1, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_1 = {regroupV0_lo[1879:1876], regroupV0_lo[1863:1860]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_1 = {regroupV0_lo[1911:1908], regroupV0_lo[1895:1892]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_lo_hi_2 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_1, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_1};
  wire [31:0]        regroupV0_lo_lo_hi_hi_hi_lo_2 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_2, regroupV0_lo_lo_hi_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_1 = {regroupV0_lo[1943:1940], regroupV0_lo[1927:1924]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_1 = {regroupV0_lo[1975:1972], regroupV0_lo[1959:1956]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_hi_lo_2 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_1, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_1 = {regroupV0_lo[2007:2004], regroupV0_lo[1991:1988]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_1 = {regroupV0_lo[2039:2036], regroupV0_lo[2023:2020]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_hi_hi_2 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_1, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_1};
  wire [31:0]        regroupV0_lo_lo_hi_hi_hi_hi_2 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_2, regroupV0_lo_lo_hi_hi_hi_hi_lo_2};
  wire [63:0]        regroupV0_lo_lo_hi_hi_hi_2 = {regroupV0_lo_lo_hi_hi_hi_hi_2, regroupV0_lo_lo_hi_hi_hi_lo_2};
  wire [127:0]       regroupV0_lo_lo_hi_hi_2 = {regroupV0_lo_lo_hi_hi_hi_2, regroupV0_lo_lo_hi_hi_lo_2};
  wire [255:0]       regroupV0_lo_lo_hi_2 = {regroupV0_lo_lo_hi_hi_2, regroupV0_lo_lo_hi_lo_2};
  wire [511:0]       regroupV0_lo_lo_2 = {regroupV0_lo_lo_hi_2, regroupV0_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_1 = {regroupV0_lo[2071:2068], regroupV0_lo[2055:2052]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_1 = {regroupV0_lo[2103:2100], regroupV0_lo[2087:2084]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_lo_lo_2 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_1, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_1 = {regroupV0_lo[2135:2132], regroupV0_lo[2119:2116]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_1 = {regroupV0_lo[2167:2164], regroupV0_lo[2151:2148]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_lo_hi_2 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_1, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_1};
  wire [31:0]        regroupV0_lo_hi_lo_lo_lo_lo_2 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_2, regroupV0_lo_hi_lo_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_1 = {regroupV0_lo[2199:2196], regroupV0_lo[2183:2180]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_1 = {regroupV0_lo[2231:2228], regroupV0_lo[2215:2212]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_hi_lo_2 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_1, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_1 = {regroupV0_lo[2263:2260], regroupV0_lo[2247:2244]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_1 = {regroupV0_lo[2295:2292], regroupV0_lo[2279:2276]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_hi_hi_2 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_1, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_1};
  wire [31:0]        regroupV0_lo_hi_lo_lo_lo_hi_2 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_2, regroupV0_lo_hi_lo_lo_lo_hi_lo_2};
  wire [63:0]        regroupV0_lo_hi_lo_lo_lo_2 = {regroupV0_lo_hi_lo_lo_lo_hi_2, regroupV0_lo_hi_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_1 = {regroupV0_lo[2327:2324], regroupV0_lo[2311:2308]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_1 = {regroupV0_lo[2359:2356], regroupV0_lo[2343:2340]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_lo_lo_2 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_1, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_1 = {regroupV0_lo[2391:2388], regroupV0_lo[2375:2372]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_1 = {regroupV0_lo[2423:2420], regroupV0_lo[2407:2404]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_lo_hi_2 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_1, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_1};
  wire [31:0]        regroupV0_lo_hi_lo_lo_hi_lo_2 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_2, regroupV0_lo_hi_lo_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_1 = {regroupV0_lo[2455:2452], regroupV0_lo[2439:2436]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_1 = {regroupV0_lo[2487:2484], regroupV0_lo[2471:2468]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_hi_lo_2 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_1, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_1 = {regroupV0_lo[2519:2516], regroupV0_lo[2503:2500]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_1 = {regroupV0_lo[2551:2548], regroupV0_lo[2535:2532]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_hi_hi_2 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_1, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_1};
  wire [31:0]        regroupV0_lo_hi_lo_lo_hi_hi_2 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_2, regroupV0_lo_hi_lo_lo_hi_hi_lo_2};
  wire [63:0]        regroupV0_lo_hi_lo_lo_hi_2 = {regroupV0_lo_hi_lo_lo_hi_hi_2, regroupV0_lo_hi_lo_lo_hi_lo_2};
  wire [127:0]       regroupV0_lo_hi_lo_lo_2 = {regroupV0_lo_hi_lo_lo_hi_2, regroupV0_lo_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_1 = {regroupV0_lo[2583:2580], regroupV0_lo[2567:2564]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_1 = {regroupV0_lo[2615:2612], regroupV0_lo[2599:2596]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_lo_lo_2 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_1, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_1 = {regroupV0_lo[2647:2644], regroupV0_lo[2631:2628]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_1 = {regroupV0_lo[2679:2676], regroupV0_lo[2663:2660]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_lo_hi_2 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_1, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_1};
  wire [31:0]        regroupV0_lo_hi_lo_hi_lo_lo_2 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_2, regroupV0_lo_hi_lo_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_1 = {regroupV0_lo[2711:2708], regroupV0_lo[2695:2692]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_1 = {regroupV0_lo[2743:2740], regroupV0_lo[2727:2724]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_hi_lo_2 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_1, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_1 = {regroupV0_lo[2775:2772], regroupV0_lo[2759:2756]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_1 = {regroupV0_lo[2807:2804], regroupV0_lo[2791:2788]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_hi_hi_2 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_1, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_1};
  wire [31:0]        regroupV0_lo_hi_lo_hi_lo_hi_2 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_2, regroupV0_lo_hi_lo_hi_lo_hi_lo_2};
  wire [63:0]        regroupV0_lo_hi_lo_hi_lo_2 = {regroupV0_lo_hi_lo_hi_lo_hi_2, regroupV0_lo_hi_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_1 = {regroupV0_lo[2839:2836], regroupV0_lo[2823:2820]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_1 = {regroupV0_lo[2871:2868], regroupV0_lo[2855:2852]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_lo_lo_2 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_1, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_1 = {regroupV0_lo[2903:2900], regroupV0_lo[2887:2884]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_1 = {regroupV0_lo[2935:2932], regroupV0_lo[2919:2916]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_lo_hi_2 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_1, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_1};
  wire [31:0]        regroupV0_lo_hi_lo_hi_hi_lo_2 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_2, regroupV0_lo_hi_lo_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_1 = {regroupV0_lo[2967:2964], regroupV0_lo[2951:2948]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_1 = {regroupV0_lo[2999:2996], regroupV0_lo[2983:2980]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_hi_lo_2 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_1, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_1 = {regroupV0_lo[3031:3028], regroupV0_lo[3015:3012]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_1 = {regroupV0_lo[3063:3060], regroupV0_lo[3047:3044]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_hi_hi_2 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_1, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_1};
  wire [31:0]        regroupV0_lo_hi_lo_hi_hi_hi_2 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_2, regroupV0_lo_hi_lo_hi_hi_hi_lo_2};
  wire [63:0]        regroupV0_lo_hi_lo_hi_hi_2 = {regroupV0_lo_hi_lo_hi_hi_hi_2, regroupV0_lo_hi_lo_hi_hi_lo_2};
  wire [127:0]       regroupV0_lo_hi_lo_hi_2 = {regroupV0_lo_hi_lo_hi_hi_2, regroupV0_lo_hi_lo_hi_lo_2};
  wire [255:0]       regroupV0_lo_hi_lo_2 = {regroupV0_lo_hi_lo_hi_2, regroupV0_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_1 = {regroupV0_lo[3095:3092], regroupV0_lo[3079:3076]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_1 = {regroupV0_lo[3127:3124], regroupV0_lo[3111:3108]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_lo_lo_2 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_1, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_1 = {regroupV0_lo[3159:3156], regroupV0_lo[3143:3140]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_1 = {regroupV0_lo[3191:3188], regroupV0_lo[3175:3172]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_lo_hi_2 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_1, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_1};
  wire [31:0]        regroupV0_lo_hi_hi_lo_lo_lo_2 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_2, regroupV0_lo_hi_hi_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_1 = {regroupV0_lo[3223:3220], regroupV0_lo[3207:3204]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_1 = {regroupV0_lo[3255:3252], regroupV0_lo[3239:3236]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_hi_lo_2 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_1, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_1 = {regroupV0_lo[3287:3284], regroupV0_lo[3271:3268]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_1 = {regroupV0_lo[3319:3316], regroupV0_lo[3303:3300]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_hi_hi_2 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_1, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_1};
  wire [31:0]        regroupV0_lo_hi_hi_lo_lo_hi_2 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_2, regroupV0_lo_hi_hi_lo_lo_hi_lo_2};
  wire [63:0]        regroupV0_lo_hi_hi_lo_lo_2 = {regroupV0_lo_hi_hi_lo_lo_hi_2, regroupV0_lo_hi_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_1 = {regroupV0_lo[3351:3348], regroupV0_lo[3335:3332]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_1 = {regroupV0_lo[3383:3380], regroupV0_lo[3367:3364]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_lo_lo_2 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_1, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_1 = {regroupV0_lo[3415:3412], regroupV0_lo[3399:3396]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_1 = {regroupV0_lo[3447:3444], regroupV0_lo[3431:3428]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_lo_hi_2 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_1, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_1};
  wire [31:0]        regroupV0_lo_hi_hi_lo_hi_lo_2 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_2, regroupV0_lo_hi_hi_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_1 = {regroupV0_lo[3479:3476], regroupV0_lo[3463:3460]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_1 = {regroupV0_lo[3511:3508], regroupV0_lo[3495:3492]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_hi_lo_2 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_1, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_1 = {regroupV0_lo[3543:3540], regroupV0_lo[3527:3524]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_1 = {regroupV0_lo[3575:3572], regroupV0_lo[3559:3556]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_hi_hi_2 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_1, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_1};
  wire [31:0]        regroupV0_lo_hi_hi_lo_hi_hi_2 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_2, regroupV0_lo_hi_hi_lo_hi_hi_lo_2};
  wire [63:0]        regroupV0_lo_hi_hi_lo_hi_2 = {regroupV0_lo_hi_hi_lo_hi_hi_2, regroupV0_lo_hi_hi_lo_hi_lo_2};
  wire [127:0]       regroupV0_lo_hi_hi_lo_2 = {regroupV0_lo_hi_hi_lo_hi_2, regroupV0_lo_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_1 = {regroupV0_lo[3607:3604], regroupV0_lo[3591:3588]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_1 = {regroupV0_lo[3639:3636], regroupV0_lo[3623:3620]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_lo_lo_2 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_1, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_1 = {regroupV0_lo[3671:3668], regroupV0_lo[3655:3652]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_1 = {regroupV0_lo[3703:3700], regroupV0_lo[3687:3684]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_lo_hi_2 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_1, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_1};
  wire [31:0]        regroupV0_lo_hi_hi_hi_lo_lo_2 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_2, regroupV0_lo_hi_hi_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_1 = {regroupV0_lo[3735:3732], regroupV0_lo[3719:3716]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_1 = {regroupV0_lo[3767:3764], regroupV0_lo[3751:3748]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_hi_lo_2 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_1, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_1 = {regroupV0_lo[3799:3796], regroupV0_lo[3783:3780]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_1 = {regroupV0_lo[3831:3828], regroupV0_lo[3815:3812]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_hi_hi_2 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_1, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_1};
  wire [31:0]        regroupV0_lo_hi_hi_hi_lo_hi_2 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_2, regroupV0_lo_hi_hi_hi_lo_hi_lo_2};
  wire [63:0]        regroupV0_lo_hi_hi_hi_lo_2 = {regroupV0_lo_hi_hi_hi_lo_hi_2, regroupV0_lo_hi_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_1 = {regroupV0_lo[3863:3860], regroupV0_lo[3847:3844]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_1 = {regroupV0_lo[3895:3892], regroupV0_lo[3879:3876]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_lo_lo_2 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_1, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_1 = {regroupV0_lo[3927:3924], regroupV0_lo[3911:3908]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_1 = {regroupV0_lo[3959:3956], regroupV0_lo[3943:3940]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_lo_hi_2 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_1, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_1};
  wire [31:0]        regroupV0_lo_hi_hi_hi_hi_lo_2 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_2, regroupV0_lo_hi_hi_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_1 = {regroupV0_lo[3991:3988], regroupV0_lo[3975:3972]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_1 = {regroupV0_lo[4023:4020], regroupV0_lo[4007:4004]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_hi_lo_2 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_1, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_1 = {regroupV0_lo[4055:4052], regroupV0_lo[4039:4036]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_1 = {regroupV0_lo[4087:4084], regroupV0_lo[4071:4068]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_hi_hi_2 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_1, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_1};
  wire [31:0]        regroupV0_lo_hi_hi_hi_hi_hi_2 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_2, regroupV0_lo_hi_hi_hi_hi_hi_lo_2};
  wire [63:0]        regroupV0_lo_hi_hi_hi_hi_2 = {regroupV0_lo_hi_hi_hi_hi_hi_2, regroupV0_lo_hi_hi_hi_hi_lo_2};
  wire [127:0]       regroupV0_lo_hi_hi_hi_2 = {regroupV0_lo_hi_hi_hi_hi_2, regroupV0_lo_hi_hi_hi_lo_2};
  wire [255:0]       regroupV0_lo_hi_hi_2 = {regroupV0_lo_hi_hi_hi_2, regroupV0_lo_hi_hi_lo_2};
  wire [511:0]       regroupV0_lo_hi_2 = {regroupV0_lo_hi_hi_2, regroupV0_lo_hi_lo_2};
  wire [1023:0]      regroupV0_lo_2 = {regroupV0_lo_hi_2, regroupV0_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_1 = {regroupV0_hi[23:20], regroupV0_hi[7:4]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_1 = {regroupV0_hi[55:52], regroupV0_hi[39:36]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_lo_lo_2 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_1 = {regroupV0_hi[87:84], regroupV0_hi[71:68]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_1 = {regroupV0_hi[119:116], regroupV0_hi[103:100]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_lo_hi_2 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_1, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_1};
  wire [31:0]        regroupV0_hi_lo_lo_lo_lo_lo_2 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_1 = {regroupV0_hi[151:148], regroupV0_hi[135:132]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_1 = {regroupV0_hi[183:180], regroupV0_hi[167:164]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_hi_lo_2 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_1, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_1 = {regroupV0_hi[215:212], regroupV0_hi[199:196]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_1 = {regroupV0_hi[247:244], regroupV0_hi[231:228]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_hi_hi_2 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_1, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_1};
  wire [31:0]        regroupV0_hi_lo_lo_lo_lo_hi_2 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_2, regroupV0_hi_lo_lo_lo_lo_hi_lo_2};
  wire [63:0]        regroupV0_hi_lo_lo_lo_lo_2 = {regroupV0_hi_lo_lo_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_1 = {regroupV0_hi[279:276], regroupV0_hi[263:260]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_1 = {regroupV0_hi[311:308], regroupV0_hi[295:292]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_lo_lo_2 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_1 = {regroupV0_hi[343:340], regroupV0_hi[327:324]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_1 = {regroupV0_hi[375:372], regroupV0_hi[359:356]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_lo_hi_2 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_1, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_1};
  wire [31:0]        regroupV0_hi_lo_lo_lo_hi_lo_2 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_2, regroupV0_hi_lo_lo_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_1 = {regroupV0_hi[407:404], regroupV0_hi[391:388]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_1 = {regroupV0_hi[439:436], regroupV0_hi[423:420]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_hi_lo_2 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_1, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_1 = {regroupV0_hi[471:468], regroupV0_hi[455:452]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_1 = {regroupV0_hi[503:500], regroupV0_hi[487:484]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_hi_hi_2 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_1, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_1};
  wire [31:0]        regroupV0_hi_lo_lo_lo_hi_hi_2 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_2, regroupV0_hi_lo_lo_lo_hi_hi_lo_2};
  wire [63:0]        regroupV0_hi_lo_lo_lo_hi_2 = {regroupV0_hi_lo_lo_lo_hi_hi_2, regroupV0_hi_lo_lo_lo_hi_lo_2};
  wire [127:0]       regroupV0_hi_lo_lo_lo_2 = {regroupV0_hi_lo_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_1 = {regroupV0_hi[535:532], regroupV0_hi[519:516]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_1 = {regroupV0_hi[567:564], regroupV0_hi[551:548]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_lo_lo_2 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_1, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_1 = {regroupV0_hi[599:596], regroupV0_hi[583:580]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_1 = {regroupV0_hi[631:628], regroupV0_hi[615:612]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_lo_hi_2 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_1, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_1};
  wire [31:0]        regroupV0_hi_lo_lo_hi_lo_lo_2 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_2, regroupV0_hi_lo_lo_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_1 = {regroupV0_hi[663:660], regroupV0_hi[647:644]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_1 = {regroupV0_hi[695:692], regroupV0_hi[679:676]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_hi_lo_2 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_1, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_1 = {regroupV0_hi[727:724], regroupV0_hi[711:708]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_1 = {regroupV0_hi[759:756], regroupV0_hi[743:740]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_hi_hi_2 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_1, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_1};
  wire [31:0]        regroupV0_hi_lo_lo_hi_lo_hi_2 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_2, regroupV0_hi_lo_lo_hi_lo_hi_lo_2};
  wire [63:0]        regroupV0_hi_lo_lo_hi_lo_2 = {regroupV0_hi_lo_lo_hi_lo_hi_2, regroupV0_hi_lo_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_1 = {regroupV0_hi[791:788], regroupV0_hi[775:772]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_1 = {regroupV0_hi[823:820], regroupV0_hi[807:804]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_lo_lo_2 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_1, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_1 = {regroupV0_hi[855:852], regroupV0_hi[839:836]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_1 = {regroupV0_hi[887:884], regroupV0_hi[871:868]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_lo_hi_2 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_1, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_1};
  wire [31:0]        regroupV0_hi_lo_lo_hi_hi_lo_2 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_2, regroupV0_hi_lo_lo_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_1 = {regroupV0_hi[919:916], regroupV0_hi[903:900]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_1 = {regroupV0_hi[951:948], regroupV0_hi[935:932]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_hi_lo_2 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_1, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_1 = {regroupV0_hi[983:980], regroupV0_hi[967:964]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_1 = {regroupV0_hi[1015:1012], regroupV0_hi[999:996]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_hi_hi_2 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_1, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_1};
  wire [31:0]        regroupV0_hi_lo_lo_hi_hi_hi_2 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_2, regroupV0_hi_lo_lo_hi_hi_hi_lo_2};
  wire [63:0]        regroupV0_hi_lo_lo_hi_hi_2 = {regroupV0_hi_lo_lo_hi_hi_hi_2, regroupV0_hi_lo_lo_hi_hi_lo_2};
  wire [127:0]       regroupV0_hi_lo_lo_hi_2 = {regroupV0_hi_lo_lo_hi_hi_2, regroupV0_hi_lo_lo_hi_lo_2};
  wire [255:0]       regroupV0_hi_lo_lo_2 = {regroupV0_hi_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_1 = {regroupV0_hi[1047:1044], regroupV0_hi[1031:1028]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_1 = {regroupV0_hi[1079:1076], regroupV0_hi[1063:1060]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_lo_lo_2 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_1, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_1 = {regroupV0_hi[1111:1108], regroupV0_hi[1095:1092]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_1 = {regroupV0_hi[1143:1140], regroupV0_hi[1127:1124]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_lo_hi_2 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_1, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_1};
  wire [31:0]        regroupV0_hi_lo_hi_lo_lo_lo_2 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_2, regroupV0_hi_lo_hi_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_1 = {regroupV0_hi[1175:1172], regroupV0_hi[1159:1156]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_1 = {regroupV0_hi[1207:1204], regroupV0_hi[1191:1188]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_hi_lo_2 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_1, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_1 = {regroupV0_hi[1239:1236], regroupV0_hi[1223:1220]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_1 = {regroupV0_hi[1271:1268], regroupV0_hi[1255:1252]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_hi_hi_2 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_1, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_1};
  wire [31:0]        regroupV0_hi_lo_hi_lo_lo_hi_2 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_2, regroupV0_hi_lo_hi_lo_lo_hi_lo_2};
  wire [63:0]        regroupV0_hi_lo_hi_lo_lo_2 = {regroupV0_hi_lo_hi_lo_lo_hi_2, regroupV0_hi_lo_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_1 = {regroupV0_hi[1303:1300], regroupV0_hi[1287:1284]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_1 = {regroupV0_hi[1335:1332], regroupV0_hi[1319:1316]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_lo_lo_2 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_1, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_1 = {regroupV0_hi[1367:1364], regroupV0_hi[1351:1348]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_1 = {regroupV0_hi[1399:1396], regroupV0_hi[1383:1380]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_lo_hi_2 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_1, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_1};
  wire [31:0]        regroupV0_hi_lo_hi_lo_hi_lo_2 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_2, regroupV0_hi_lo_hi_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_1 = {regroupV0_hi[1431:1428], regroupV0_hi[1415:1412]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_1 = {regroupV0_hi[1463:1460], regroupV0_hi[1447:1444]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_hi_lo_2 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_1, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_1 = {regroupV0_hi[1495:1492], regroupV0_hi[1479:1476]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_1 = {regroupV0_hi[1527:1524], regroupV0_hi[1511:1508]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_hi_hi_2 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_1, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_1};
  wire [31:0]        regroupV0_hi_lo_hi_lo_hi_hi_2 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_2, regroupV0_hi_lo_hi_lo_hi_hi_lo_2};
  wire [63:0]        regroupV0_hi_lo_hi_lo_hi_2 = {regroupV0_hi_lo_hi_lo_hi_hi_2, regroupV0_hi_lo_hi_lo_hi_lo_2};
  wire [127:0]       regroupV0_hi_lo_hi_lo_2 = {regroupV0_hi_lo_hi_lo_hi_2, regroupV0_hi_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_1 = {regroupV0_hi[1559:1556], regroupV0_hi[1543:1540]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_1 = {regroupV0_hi[1591:1588], regroupV0_hi[1575:1572]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_lo_lo_2 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_1, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_1 = {regroupV0_hi[1623:1620], regroupV0_hi[1607:1604]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_1 = {regroupV0_hi[1655:1652], regroupV0_hi[1639:1636]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_lo_hi_2 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_1, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_1};
  wire [31:0]        regroupV0_hi_lo_hi_hi_lo_lo_2 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_2, regroupV0_hi_lo_hi_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_1 = {regroupV0_hi[1687:1684], regroupV0_hi[1671:1668]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_1 = {regroupV0_hi[1719:1716], regroupV0_hi[1703:1700]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_hi_lo_2 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_1, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_1 = {regroupV0_hi[1751:1748], regroupV0_hi[1735:1732]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_1 = {regroupV0_hi[1783:1780], regroupV0_hi[1767:1764]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_hi_hi_2 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_1, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_1};
  wire [31:0]        regroupV0_hi_lo_hi_hi_lo_hi_2 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_2, regroupV0_hi_lo_hi_hi_lo_hi_lo_2};
  wire [63:0]        regroupV0_hi_lo_hi_hi_lo_2 = {regroupV0_hi_lo_hi_hi_lo_hi_2, regroupV0_hi_lo_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_1 = {regroupV0_hi[1815:1812], regroupV0_hi[1799:1796]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_1 = {regroupV0_hi[1847:1844], regroupV0_hi[1831:1828]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_lo_lo_2 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_1, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_1 = {regroupV0_hi[1879:1876], regroupV0_hi[1863:1860]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_1 = {regroupV0_hi[1911:1908], regroupV0_hi[1895:1892]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_lo_hi_2 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_1, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_1};
  wire [31:0]        regroupV0_hi_lo_hi_hi_hi_lo_2 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_2, regroupV0_hi_lo_hi_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_1 = {regroupV0_hi[1943:1940], regroupV0_hi[1927:1924]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_1 = {regroupV0_hi[1975:1972], regroupV0_hi[1959:1956]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_hi_lo_2 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_1, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_1 = {regroupV0_hi[2007:2004], regroupV0_hi[1991:1988]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_1 = {regroupV0_hi[2039:2036], regroupV0_hi[2023:2020]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_hi_hi_2 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_1, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_1};
  wire [31:0]        regroupV0_hi_lo_hi_hi_hi_hi_2 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_2, regroupV0_hi_lo_hi_hi_hi_hi_lo_2};
  wire [63:0]        regroupV0_hi_lo_hi_hi_hi_2 = {regroupV0_hi_lo_hi_hi_hi_hi_2, regroupV0_hi_lo_hi_hi_hi_lo_2};
  wire [127:0]       regroupV0_hi_lo_hi_hi_2 = {regroupV0_hi_lo_hi_hi_hi_2, regroupV0_hi_lo_hi_hi_lo_2};
  wire [255:0]       regroupV0_hi_lo_hi_2 = {regroupV0_hi_lo_hi_hi_2, regroupV0_hi_lo_hi_lo_2};
  wire [511:0]       regroupV0_hi_lo_2 = {regroupV0_hi_lo_hi_2, regroupV0_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_1 = {regroupV0_hi[2071:2068], regroupV0_hi[2055:2052]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_1 = {regroupV0_hi[2103:2100], regroupV0_hi[2087:2084]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_lo_lo_2 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_1, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_1 = {regroupV0_hi[2135:2132], regroupV0_hi[2119:2116]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_1 = {regroupV0_hi[2167:2164], regroupV0_hi[2151:2148]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_lo_hi_2 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_1, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_1};
  wire [31:0]        regroupV0_hi_hi_lo_lo_lo_lo_2 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_2, regroupV0_hi_hi_lo_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_1 = {regroupV0_hi[2199:2196], regroupV0_hi[2183:2180]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_1 = {regroupV0_hi[2231:2228], regroupV0_hi[2215:2212]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_hi_lo_2 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_1, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_1 = {regroupV0_hi[2263:2260], regroupV0_hi[2247:2244]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_1 = {regroupV0_hi[2295:2292], regroupV0_hi[2279:2276]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_hi_hi_2 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_1, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_1};
  wire [31:0]        regroupV0_hi_hi_lo_lo_lo_hi_2 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_2, regroupV0_hi_hi_lo_lo_lo_hi_lo_2};
  wire [63:0]        regroupV0_hi_hi_lo_lo_lo_2 = {regroupV0_hi_hi_lo_lo_lo_hi_2, regroupV0_hi_hi_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_1 = {regroupV0_hi[2327:2324], regroupV0_hi[2311:2308]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_1 = {regroupV0_hi[2359:2356], regroupV0_hi[2343:2340]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_lo_lo_2 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_1, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_1 = {regroupV0_hi[2391:2388], regroupV0_hi[2375:2372]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_1 = {regroupV0_hi[2423:2420], regroupV0_hi[2407:2404]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_lo_hi_2 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_1, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_1};
  wire [31:0]        regroupV0_hi_hi_lo_lo_hi_lo_2 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_2, regroupV0_hi_hi_lo_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_1 = {regroupV0_hi[2455:2452], regroupV0_hi[2439:2436]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_1 = {regroupV0_hi[2487:2484], regroupV0_hi[2471:2468]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_hi_lo_2 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_1, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_1 = {regroupV0_hi[2519:2516], regroupV0_hi[2503:2500]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_1 = {regroupV0_hi[2551:2548], regroupV0_hi[2535:2532]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_hi_hi_2 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_1, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_1};
  wire [31:0]        regroupV0_hi_hi_lo_lo_hi_hi_2 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_2, regroupV0_hi_hi_lo_lo_hi_hi_lo_2};
  wire [63:0]        regroupV0_hi_hi_lo_lo_hi_2 = {regroupV0_hi_hi_lo_lo_hi_hi_2, regroupV0_hi_hi_lo_lo_hi_lo_2};
  wire [127:0]       regroupV0_hi_hi_lo_lo_2 = {regroupV0_hi_hi_lo_lo_hi_2, regroupV0_hi_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_1 = {regroupV0_hi[2583:2580], regroupV0_hi[2567:2564]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_1 = {regroupV0_hi[2615:2612], regroupV0_hi[2599:2596]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_lo_lo_2 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_1, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_1 = {regroupV0_hi[2647:2644], regroupV0_hi[2631:2628]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_1 = {regroupV0_hi[2679:2676], regroupV0_hi[2663:2660]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_lo_hi_2 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_1, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_1};
  wire [31:0]        regroupV0_hi_hi_lo_hi_lo_lo_2 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_2, regroupV0_hi_hi_lo_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_1 = {regroupV0_hi[2711:2708], regroupV0_hi[2695:2692]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_1 = {regroupV0_hi[2743:2740], regroupV0_hi[2727:2724]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_hi_lo_2 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_1, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_1 = {regroupV0_hi[2775:2772], regroupV0_hi[2759:2756]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_1 = {regroupV0_hi[2807:2804], regroupV0_hi[2791:2788]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_hi_hi_2 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_1, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_1};
  wire [31:0]        regroupV0_hi_hi_lo_hi_lo_hi_2 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_2, regroupV0_hi_hi_lo_hi_lo_hi_lo_2};
  wire [63:0]        regroupV0_hi_hi_lo_hi_lo_2 = {regroupV0_hi_hi_lo_hi_lo_hi_2, regroupV0_hi_hi_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_1 = {regroupV0_hi[2839:2836], regroupV0_hi[2823:2820]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_1 = {regroupV0_hi[2871:2868], regroupV0_hi[2855:2852]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_lo_lo_2 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_1, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_1 = {regroupV0_hi[2903:2900], regroupV0_hi[2887:2884]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_1 = {regroupV0_hi[2935:2932], regroupV0_hi[2919:2916]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_lo_hi_2 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_1, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_1};
  wire [31:0]        regroupV0_hi_hi_lo_hi_hi_lo_2 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_2, regroupV0_hi_hi_lo_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_1 = {regroupV0_hi[2967:2964], regroupV0_hi[2951:2948]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_1 = {regroupV0_hi[2999:2996], regroupV0_hi[2983:2980]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_hi_lo_2 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_1, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_1 = {regroupV0_hi[3031:3028], regroupV0_hi[3015:3012]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_1 = {regroupV0_hi[3063:3060], regroupV0_hi[3047:3044]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_hi_hi_2 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_1, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_1};
  wire [31:0]        regroupV0_hi_hi_lo_hi_hi_hi_2 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_2, regroupV0_hi_hi_lo_hi_hi_hi_lo_2};
  wire [63:0]        regroupV0_hi_hi_lo_hi_hi_2 = {regroupV0_hi_hi_lo_hi_hi_hi_2, regroupV0_hi_hi_lo_hi_hi_lo_2};
  wire [127:0]       regroupV0_hi_hi_lo_hi_2 = {regroupV0_hi_hi_lo_hi_hi_2, regroupV0_hi_hi_lo_hi_lo_2};
  wire [255:0]       regroupV0_hi_hi_lo_2 = {regroupV0_hi_hi_lo_hi_2, regroupV0_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_1 = {regroupV0_hi[3095:3092], regroupV0_hi[3079:3076]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_1 = {regroupV0_hi[3127:3124], regroupV0_hi[3111:3108]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_lo_lo_2 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_1, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_1 = {regroupV0_hi[3159:3156], regroupV0_hi[3143:3140]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_1 = {regroupV0_hi[3191:3188], regroupV0_hi[3175:3172]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_lo_hi_2 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_1, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_1};
  wire [31:0]        regroupV0_hi_hi_hi_lo_lo_lo_2 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_2, regroupV0_hi_hi_hi_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_1 = {regroupV0_hi[3223:3220], regroupV0_hi[3207:3204]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_1 = {regroupV0_hi[3255:3252], regroupV0_hi[3239:3236]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_hi_lo_2 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_1, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_1 = {regroupV0_hi[3287:3284], regroupV0_hi[3271:3268]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_1 = {regroupV0_hi[3319:3316], regroupV0_hi[3303:3300]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_hi_hi_2 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_1, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_1};
  wire [31:0]        regroupV0_hi_hi_hi_lo_lo_hi_2 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_2, regroupV0_hi_hi_hi_lo_lo_hi_lo_2};
  wire [63:0]        regroupV0_hi_hi_hi_lo_lo_2 = {regroupV0_hi_hi_hi_lo_lo_hi_2, regroupV0_hi_hi_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_1 = {regroupV0_hi[3351:3348], regroupV0_hi[3335:3332]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_1 = {regroupV0_hi[3383:3380], regroupV0_hi[3367:3364]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_lo_lo_2 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_1, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_1 = {regroupV0_hi[3415:3412], regroupV0_hi[3399:3396]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_1 = {regroupV0_hi[3447:3444], regroupV0_hi[3431:3428]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_lo_hi_2 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_1, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_1};
  wire [31:0]        regroupV0_hi_hi_hi_lo_hi_lo_2 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_2, regroupV0_hi_hi_hi_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_1 = {regroupV0_hi[3479:3476], regroupV0_hi[3463:3460]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_1 = {regroupV0_hi[3511:3508], regroupV0_hi[3495:3492]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_hi_lo_2 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_1, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_1 = {regroupV0_hi[3543:3540], regroupV0_hi[3527:3524]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_1 = {regroupV0_hi[3575:3572], regroupV0_hi[3559:3556]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_hi_hi_2 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_1};
  wire [31:0]        regroupV0_hi_hi_hi_lo_hi_hi_2 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_2, regroupV0_hi_hi_hi_lo_hi_hi_lo_2};
  wire [63:0]        regroupV0_hi_hi_hi_lo_hi_2 = {regroupV0_hi_hi_hi_lo_hi_hi_2, regroupV0_hi_hi_hi_lo_hi_lo_2};
  wire [127:0]       regroupV0_hi_hi_hi_lo_2 = {regroupV0_hi_hi_hi_lo_hi_2, regroupV0_hi_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_1 = {regroupV0_hi[3607:3604], regroupV0_hi[3591:3588]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_1 = {regroupV0_hi[3639:3636], regroupV0_hi[3623:3620]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_lo_lo_2 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_1, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_1 = {regroupV0_hi[3671:3668], regroupV0_hi[3655:3652]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_1 = {regroupV0_hi[3703:3700], regroupV0_hi[3687:3684]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_lo_hi_2 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_1, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_1};
  wire [31:0]        regroupV0_hi_hi_hi_hi_lo_lo_2 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_2, regroupV0_hi_hi_hi_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_1 = {regroupV0_hi[3735:3732], regroupV0_hi[3719:3716]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_1 = {regroupV0_hi[3767:3764], regroupV0_hi[3751:3748]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_hi_lo_2 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_1, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_1 = {regroupV0_hi[3799:3796], regroupV0_hi[3783:3780]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_1 = {regroupV0_hi[3831:3828], regroupV0_hi[3815:3812]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_hi_hi_2 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_1, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_1};
  wire [31:0]        regroupV0_hi_hi_hi_hi_lo_hi_2 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_2, regroupV0_hi_hi_hi_hi_lo_hi_lo_2};
  wire [63:0]        regroupV0_hi_hi_hi_hi_lo_2 = {regroupV0_hi_hi_hi_hi_lo_hi_2, regroupV0_hi_hi_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_1 = {regroupV0_hi[3863:3860], regroupV0_hi[3847:3844]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_1 = {regroupV0_hi[3895:3892], regroupV0_hi[3879:3876]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_lo_lo_2 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_1, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_1 = {regroupV0_hi[3927:3924], regroupV0_hi[3911:3908]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_1 = {regroupV0_hi[3959:3956], regroupV0_hi[3943:3940]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_lo_hi_2 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_1, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_1};
  wire [31:0]        regroupV0_hi_hi_hi_hi_hi_lo_2 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_2, regroupV0_hi_hi_hi_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_1 = {regroupV0_hi[3991:3988], regroupV0_hi[3975:3972]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_1 = {regroupV0_hi[4023:4020], regroupV0_hi[4007:4004]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_hi_lo_2 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_1, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_1 = {regroupV0_hi[4055:4052], regroupV0_hi[4039:4036]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_1 = {regroupV0_hi[4087:4084], regroupV0_hi[4071:4068]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_hi_hi_2 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_1};
  wire [31:0]        regroupV0_hi_hi_hi_hi_hi_hi_2 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_hi_hi_hi_lo_2};
  wire [63:0]        regroupV0_hi_hi_hi_hi_hi_2 = {regroupV0_hi_hi_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_hi_hi_lo_2};
  wire [127:0]       regroupV0_hi_hi_hi_hi_2 = {regroupV0_hi_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_hi_lo_2};
  wire [255:0]       regroupV0_hi_hi_hi_2 = {regroupV0_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_lo_2};
  wire [511:0]       regroupV0_hi_hi_2 = {regroupV0_hi_hi_hi_2, regroupV0_hi_hi_lo_2};
  wire [1023:0]      regroupV0_hi_2 = {regroupV0_hi_hi_2, regroupV0_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_2 = {regroupV0_lo[27:24], regroupV0_lo[11:8]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_2 = {regroupV0_lo[59:56], regroupV0_lo[43:40]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_lo_lo_3 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_2 = {regroupV0_lo[91:88], regroupV0_lo[75:72]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_2 = {regroupV0_lo[123:120], regroupV0_lo[107:104]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_lo_hi_3 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_2, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_2};
  wire [31:0]        regroupV0_lo_lo_lo_lo_lo_lo_3 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_2 = {regroupV0_lo[155:152], regroupV0_lo[139:136]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_2 = {regroupV0_lo[187:184], regroupV0_lo[171:168]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_hi_lo_3 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_2, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_2 = {regroupV0_lo[219:216], regroupV0_lo[203:200]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_2 = {regroupV0_lo[251:248], regroupV0_lo[235:232]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_hi_hi_3 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_2, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_2};
  wire [31:0]        regroupV0_lo_lo_lo_lo_lo_hi_3 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_3, regroupV0_lo_lo_lo_lo_lo_hi_lo_3};
  wire [63:0]        regroupV0_lo_lo_lo_lo_lo_3 = {regroupV0_lo_lo_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_2 = {regroupV0_lo[283:280], regroupV0_lo[267:264]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_2 = {regroupV0_lo[315:312], regroupV0_lo[299:296]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_lo_lo_3 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_2 = {regroupV0_lo[347:344], regroupV0_lo[331:328]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_2 = {regroupV0_lo[379:376], regroupV0_lo[363:360]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_lo_hi_3 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_2, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_2};
  wire [31:0]        regroupV0_lo_lo_lo_lo_hi_lo_3 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_3, regroupV0_lo_lo_lo_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_2 = {regroupV0_lo[411:408], regroupV0_lo[395:392]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_2 = {regroupV0_lo[443:440], regroupV0_lo[427:424]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_hi_lo_3 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_2, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_2 = {regroupV0_lo[475:472], regroupV0_lo[459:456]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_2 = {regroupV0_lo[507:504], regroupV0_lo[491:488]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_hi_hi_3 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_2, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_2};
  wire [31:0]        regroupV0_lo_lo_lo_lo_hi_hi_3 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_3, regroupV0_lo_lo_lo_lo_hi_hi_lo_3};
  wire [63:0]        regroupV0_lo_lo_lo_lo_hi_3 = {regroupV0_lo_lo_lo_lo_hi_hi_3, regroupV0_lo_lo_lo_lo_hi_lo_3};
  wire [127:0]       regroupV0_lo_lo_lo_lo_3 = {regroupV0_lo_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_2 = {regroupV0_lo[539:536], regroupV0_lo[523:520]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_2 = {regroupV0_lo[571:568], regroupV0_lo[555:552]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_lo_lo_3 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_2 = {regroupV0_lo[603:600], regroupV0_lo[587:584]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_2 = {regroupV0_lo[635:632], regroupV0_lo[619:616]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_lo_hi_3 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_2, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_2};
  wire [31:0]        regroupV0_lo_lo_lo_hi_lo_lo_3 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_3, regroupV0_lo_lo_lo_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_2 = {regroupV0_lo[667:664], regroupV0_lo[651:648]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_2 = {regroupV0_lo[699:696], regroupV0_lo[683:680]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_hi_lo_3 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_2, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_2 = {regroupV0_lo[731:728], regroupV0_lo[715:712]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_2 = {regroupV0_lo[763:760], regroupV0_lo[747:744]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_hi_hi_3 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_2, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_2};
  wire [31:0]        regroupV0_lo_lo_lo_hi_lo_hi_3 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_3, regroupV0_lo_lo_lo_hi_lo_hi_lo_3};
  wire [63:0]        regroupV0_lo_lo_lo_hi_lo_3 = {regroupV0_lo_lo_lo_hi_lo_hi_3, regroupV0_lo_lo_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_2 = {regroupV0_lo[795:792], regroupV0_lo[779:776]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_2 = {regroupV0_lo[827:824], regroupV0_lo[811:808]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_lo_lo_3 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_2, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_2 = {regroupV0_lo[859:856], regroupV0_lo[843:840]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_2 = {regroupV0_lo[891:888], regroupV0_lo[875:872]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_lo_hi_3 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_2, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_2};
  wire [31:0]        regroupV0_lo_lo_lo_hi_hi_lo_3 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_3, regroupV0_lo_lo_lo_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_2 = {regroupV0_lo[923:920], regroupV0_lo[907:904]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_2 = {regroupV0_lo[955:952], regroupV0_lo[939:936]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_hi_lo_3 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_2, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_2 = {regroupV0_lo[987:984], regroupV0_lo[971:968]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_2 = {regroupV0_lo[1019:1016], regroupV0_lo[1003:1000]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_hi_hi_3 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_2, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_2};
  wire [31:0]        regroupV0_lo_lo_lo_hi_hi_hi_3 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_3, regroupV0_lo_lo_lo_hi_hi_hi_lo_3};
  wire [63:0]        regroupV0_lo_lo_lo_hi_hi_3 = {regroupV0_lo_lo_lo_hi_hi_hi_3, regroupV0_lo_lo_lo_hi_hi_lo_3};
  wire [127:0]       regroupV0_lo_lo_lo_hi_3 = {regroupV0_lo_lo_lo_hi_hi_3, regroupV0_lo_lo_lo_hi_lo_3};
  wire [255:0]       regroupV0_lo_lo_lo_3 = {regroupV0_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_2 = {regroupV0_lo[1051:1048], regroupV0_lo[1035:1032]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_2 = {regroupV0_lo[1083:1080], regroupV0_lo[1067:1064]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_lo_lo_3 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_2, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_2 = {regroupV0_lo[1115:1112], regroupV0_lo[1099:1096]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_2 = {regroupV0_lo[1147:1144], regroupV0_lo[1131:1128]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_lo_hi_3 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_2, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_2};
  wire [31:0]        regroupV0_lo_lo_hi_lo_lo_lo_3 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_3, regroupV0_lo_lo_hi_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_2 = {regroupV0_lo[1179:1176], regroupV0_lo[1163:1160]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_2 = {regroupV0_lo[1211:1208], regroupV0_lo[1195:1192]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_hi_lo_3 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_2, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_2 = {regroupV0_lo[1243:1240], regroupV0_lo[1227:1224]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_2 = {regroupV0_lo[1275:1272], regroupV0_lo[1259:1256]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_hi_hi_3 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_2, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_2};
  wire [31:0]        regroupV0_lo_lo_hi_lo_lo_hi_3 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_3, regroupV0_lo_lo_hi_lo_lo_hi_lo_3};
  wire [63:0]        regroupV0_lo_lo_hi_lo_lo_3 = {regroupV0_lo_lo_hi_lo_lo_hi_3, regroupV0_lo_lo_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_2 = {regroupV0_lo[1307:1304], regroupV0_lo[1291:1288]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_2 = {regroupV0_lo[1339:1336], regroupV0_lo[1323:1320]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_lo_lo_3 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_2, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_2 = {regroupV0_lo[1371:1368], regroupV0_lo[1355:1352]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_2 = {regroupV0_lo[1403:1400], regroupV0_lo[1387:1384]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_lo_hi_3 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_2, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_2};
  wire [31:0]        regroupV0_lo_lo_hi_lo_hi_lo_3 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_3, regroupV0_lo_lo_hi_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_2 = {regroupV0_lo[1435:1432], regroupV0_lo[1419:1416]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_2 = {regroupV0_lo[1467:1464], regroupV0_lo[1451:1448]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_hi_lo_3 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_2, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_2 = {regroupV0_lo[1499:1496], regroupV0_lo[1483:1480]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_2 = {regroupV0_lo[1531:1528], regroupV0_lo[1515:1512]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_hi_hi_3 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_2, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_2};
  wire [31:0]        regroupV0_lo_lo_hi_lo_hi_hi_3 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_3, regroupV0_lo_lo_hi_lo_hi_hi_lo_3};
  wire [63:0]        regroupV0_lo_lo_hi_lo_hi_3 = {regroupV0_lo_lo_hi_lo_hi_hi_3, regroupV0_lo_lo_hi_lo_hi_lo_3};
  wire [127:0]       regroupV0_lo_lo_hi_lo_3 = {regroupV0_lo_lo_hi_lo_hi_3, regroupV0_lo_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_2 = {regroupV0_lo[1563:1560], regroupV0_lo[1547:1544]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_2 = {regroupV0_lo[1595:1592], regroupV0_lo[1579:1576]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_lo_lo_3 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_2, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_2 = {regroupV0_lo[1627:1624], regroupV0_lo[1611:1608]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_2 = {regroupV0_lo[1659:1656], regroupV0_lo[1643:1640]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_lo_hi_3 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_2, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_2};
  wire [31:0]        regroupV0_lo_lo_hi_hi_lo_lo_3 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_3, regroupV0_lo_lo_hi_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_2 = {regroupV0_lo[1691:1688], regroupV0_lo[1675:1672]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_2 = {regroupV0_lo[1723:1720], regroupV0_lo[1707:1704]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_hi_lo_3 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_2, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_2 = {regroupV0_lo[1755:1752], regroupV0_lo[1739:1736]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_2 = {regroupV0_lo[1787:1784], regroupV0_lo[1771:1768]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_hi_hi_3 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_2, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_2};
  wire [31:0]        regroupV0_lo_lo_hi_hi_lo_hi_3 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_3, regroupV0_lo_lo_hi_hi_lo_hi_lo_3};
  wire [63:0]        regroupV0_lo_lo_hi_hi_lo_3 = {regroupV0_lo_lo_hi_hi_lo_hi_3, regroupV0_lo_lo_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_2 = {regroupV0_lo[1819:1816], regroupV0_lo[1803:1800]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_2 = {regroupV0_lo[1851:1848], regroupV0_lo[1835:1832]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_lo_lo_3 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_2, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_2 = {regroupV0_lo[1883:1880], regroupV0_lo[1867:1864]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_2 = {regroupV0_lo[1915:1912], regroupV0_lo[1899:1896]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_lo_hi_3 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_2, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_2};
  wire [31:0]        regroupV0_lo_lo_hi_hi_hi_lo_3 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_3, regroupV0_lo_lo_hi_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_2 = {regroupV0_lo[1947:1944], regroupV0_lo[1931:1928]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_2 = {regroupV0_lo[1979:1976], regroupV0_lo[1963:1960]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_hi_lo_3 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_2, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_2 = {regroupV0_lo[2011:2008], regroupV0_lo[1995:1992]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_2 = {regroupV0_lo[2043:2040], regroupV0_lo[2027:2024]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_hi_hi_3 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_2, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_2};
  wire [31:0]        regroupV0_lo_lo_hi_hi_hi_hi_3 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_3, regroupV0_lo_lo_hi_hi_hi_hi_lo_3};
  wire [63:0]        regroupV0_lo_lo_hi_hi_hi_3 = {regroupV0_lo_lo_hi_hi_hi_hi_3, regroupV0_lo_lo_hi_hi_hi_lo_3};
  wire [127:0]       regroupV0_lo_lo_hi_hi_3 = {regroupV0_lo_lo_hi_hi_hi_3, regroupV0_lo_lo_hi_hi_lo_3};
  wire [255:0]       regroupV0_lo_lo_hi_3 = {regroupV0_lo_lo_hi_hi_3, regroupV0_lo_lo_hi_lo_3};
  wire [511:0]       regroupV0_lo_lo_3 = {regroupV0_lo_lo_hi_3, regroupV0_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_2 = {regroupV0_lo[2075:2072], regroupV0_lo[2059:2056]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_2 = {regroupV0_lo[2107:2104], regroupV0_lo[2091:2088]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_lo_lo_3 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_2, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_2 = {regroupV0_lo[2139:2136], regroupV0_lo[2123:2120]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_2 = {regroupV0_lo[2171:2168], regroupV0_lo[2155:2152]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_lo_hi_3 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_2, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_2};
  wire [31:0]        regroupV0_lo_hi_lo_lo_lo_lo_3 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_3, regroupV0_lo_hi_lo_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_2 = {regroupV0_lo[2203:2200], regroupV0_lo[2187:2184]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_2 = {regroupV0_lo[2235:2232], regroupV0_lo[2219:2216]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_hi_lo_3 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_2, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_2 = {regroupV0_lo[2267:2264], regroupV0_lo[2251:2248]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_2 = {regroupV0_lo[2299:2296], regroupV0_lo[2283:2280]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_hi_hi_3 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_2, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_2};
  wire [31:0]        regroupV0_lo_hi_lo_lo_lo_hi_3 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_3, regroupV0_lo_hi_lo_lo_lo_hi_lo_3};
  wire [63:0]        regroupV0_lo_hi_lo_lo_lo_3 = {regroupV0_lo_hi_lo_lo_lo_hi_3, regroupV0_lo_hi_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_2 = {regroupV0_lo[2331:2328], regroupV0_lo[2315:2312]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_2 = {regroupV0_lo[2363:2360], regroupV0_lo[2347:2344]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_lo_lo_3 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_2, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_2 = {regroupV0_lo[2395:2392], regroupV0_lo[2379:2376]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_2 = {regroupV0_lo[2427:2424], regroupV0_lo[2411:2408]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_lo_hi_3 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_2, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_2};
  wire [31:0]        regroupV0_lo_hi_lo_lo_hi_lo_3 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_3, regroupV0_lo_hi_lo_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_2 = {regroupV0_lo[2459:2456], regroupV0_lo[2443:2440]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_2 = {regroupV0_lo[2491:2488], regroupV0_lo[2475:2472]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_hi_lo_3 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_2, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_2 = {regroupV0_lo[2523:2520], regroupV0_lo[2507:2504]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_2 = {regroupV0_lo[2555:2552], regroupV0_lo[2539:2536]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_hi_hi_3 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_2, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_2};
  wire [31:0]        regroupV0_lo_hi_lo_lo_hi_hi_3 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_3, regroupV0_lo_hi_lo_lo_hi_hi_lo_3};
  wire [63:0]        regroupV0_lo_hi_lo_lo_hi_3 = {regroupV0_lo_hi_lo_lo_hi_hi_3, regroupV0_lo_hi_lo_lo_hi_lo_3};
  wire [127:0]       regroupV0_lo_hi_lo_lo_3 = {regroupV0_lo_hi_lo_lo_hi_3, regroupV0_lo_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_2 = {regroupV0_lo[2587:2584], regroupV0_lo[2571:2568]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_2 = {regroupV0_lo[2619:2616], regroupV0_lo[2603:2600]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_lo_lo_3 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_2, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_2 = {regroupV0_lo[2651:2648], regroupV0_lo[2635:2632]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_2 = {regroupV0_lo[2683:2680], regroupV0_lo[2667:2664]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_lo_hi_3 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_2, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_2};
  wire [31:0]        regroupV0_lo_hi_lo_hi_lo_lo_3 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_3, regroupV0_lo_hi_lo_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_2 = {regroupV0_lo[2715:2712], regroupV0_lo[2699:2696]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_2 = {regroupV0_lo[2747:2744], regroupV0_lo[2731:2728]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_hi_lo_3 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_2, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_2 = {regroupV0_lo[2779:2776], regroupV0_lo[2763:2760]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_2 = {regroupV0_lo[2811:2808], regroupV0_lo[2795:2792]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_hi_hi_3 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_2, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_2};
  wire [31:0]        regroupV0_lo_hi_lo_hi_lo_hi_3 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_3, regroupV0_lo_hi_lo_hi_lo_hi_lo_3};
  wire [63:0]        regroupV0_lo_hi_lo_hi_lo_3 = {regroupV0_lo_hi_lo_hi_lo_hi_3, regroupV0_lo_hi_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_2 = {regroupV0_lo[2843:2840], regroupV0_lo[2827:2824]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_2 = {regroupV0_lo[2875:2872], regroupV0_lo[2859:2856]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_lo_lo_3 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_2, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_2 = {regroupV0_lo[2907:2904], regroupV0_lo[2891:2888]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_2 = {regroupV0_lo[2939:2936], regroupV0_lo[2923:2920]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_lo_hi_3 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_2, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_2};
  wire [31:0]        regroupV0_lo_hi_lo_hi_hi_lo_3 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_3, regroupV0_lo_hi_lo_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_2 = {regroupV0_lo[2971:2968], regroupV0_lo[2955:2952]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_2 = {regroupV0_lo[3003:3000], regroupV0_lo[2987:2984]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_hi_lo_3 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_2, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_2 = {regroupV0_lo[3035:3032], regroupV0_lo[3019:3016]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_2 = {regroupV0_lo[3067:3064], regroupV0_lo[3051:3048]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_hi_hi_3 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_2, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_2};
  wire [31:0]        regroupV0_lo_hi_lo_hi_hi_hi_3 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_3, regroupV0_lo_hi_lo_hi_hi_hi_lo_3};
  wire [63:0]        regroupV0_lo_hi_lo_hi_hi_3 = {regroupV0_lo_hi_lo_hi_hi_hi_3, regroupV0_lo_hi_lo_hi_hi_lo_3};
  wire [127:0]       regroupV0_lo_hi_lo_hi_3 = {regroupV0_lo_hi_lo_hi_hi_3, regroupV0_lo_hi_lo_hi_lo_3};
  wire [255:0]       regroupV0_lo_hi_lo_3 = {regroupV0_lo_hi_lo_hi_3, regroupV0_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_2 = {regroupV0_lo[3099:3096], regroupV0_lo[3083:3080]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_2 = {regroupV0_lo[3131:3128], regroupV0_lo[3115:3112]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_lo_lo_3 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_2, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_2 = {regroupV0_lo[3163:3160], regroupV0_lo[3147:3144]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_2 = {regroupV0_lo[3195:3192], regroupV0_lo[3179:3176]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_lo_hi_3 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_2, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_2};
  wire [31:0]        regroupV0_lo_hi_hi_lo_lo_lo_3 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_3, regroupV0_lo_hi_hi_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_2 = {regroupV0_lo[3227:3224], regroupV0_lo[3211:3208]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_2 = {regroupV0_lo[3259:3256], regroupV0_lo[3243:3240]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_hi_lo_3 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_2, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_2 = {regroupV0_lo[3291:3288], regroupV0_lo[3275:3272]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_2 = {regroupV0_lo[3323:3320], regroupV0_lo[3307:3304]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_hi_hi_3 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_2, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_2};
  wire [31:0]        regroupV0_lo_hi_hi_lo_lo_hi_3 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_3, regroupV0_lo_hi_hi_lo_lo_hi_lo_3};
  wire [63:0]        regroupV0_lo_hi_hi_lo_lo_3 = {regroupV0_lo_hi_hi_lo_lo_hi_3, regroupV0_lo_hi_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_2 = {regroupV0_lo[3355:3352], regroupV0_lo[3339:3336]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_2 = {regroupV0_lo[3387:3384], regroupV0_lo[3371:3368]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_lo_lo_3 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_2, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_2 = {regroupV0_lo[3419:3416], regroupV0_lo[3403:3400]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_2 = {regroupV0_lo[3451:3448], regroupV0_lo[3435:3432]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_lo_hi_3 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_2, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_2};
  wire [31:0]        regroupV0_lo_hi_hi_lo_hi_lo_3 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_3, regroupV0_lo_hi_hi_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_2 = {regroupV0_lo[3483:3480], regroupV0_lo[3467:3464]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_2 = {regroupV0_lo[3515:3512], regroupV0_lo[3499:3496]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_hi_lo_3 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_2, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_2 = {regroupV0_lo[3547:3544], regroupV0_lo[3531:3528]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_2 = {regroupV0_lo[3579:3576], regroupV0_lo[3563:3560]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_hi_hi_3 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_2, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_2};
  wire [31:0]        regroupV0_lo_hi_hi_lo_hi_hi_3 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_3, regroupV0_lo_hi_hi_lo_hi_hi_lo_3};
  wire [63:0]        regroupV0_lo_hi_hi_lo_hi_3 = {regroupV0_lo_hi_hi_lo_hi_hi_3, regroupV0_lo_hi_hi_lo_hi_lo_3};
  wire [127:0]       regroupV0_lo_hi_hi_lo_3 = {regroupV0_lo_hi_hi_lo_hi_3, regroupV0_lo_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_2 = {regroupV0_lo[3611:3608], regroupV0_lo[3595:3592]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_2 = {regroupV0_lo[3643:3640], regroupV0_lo[3627:3624]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_lo_lo_3 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_2, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_2 = {regroupV0_lo[3675:3672], regroupV0_lo[3659:3656]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_2 = {regroupV0_lo[3707:3704], regroupV0_lo[3691:3688]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_lo_hi_3 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_2, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_2};
  wire [31:0]        regroupV0_lo_hi_hi_hi_lo_lo_3 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_3, regroupV0_lo_hi_hi_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_2 = {regroupV0_lo[3739:3736], regroupV0_lo[3723:3720]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_2 = {regroupV0_lo[3771:3768], regroupV0_lo[3755:3752]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_hi_lo_3 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_2, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_2 = {regroupV0_lo[3803:3800], regroupV0_lo[3787:3784]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_2 = {regroupV0_lo[3835:3832], regroupV0_lo[3819:3816]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_hi_hi_3 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_2, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_2};
  wire [31:0]        regroupV0_lo_hi_hi_hi_lo_hi_3 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_3, regroupV0_lo_hi_hi_hi_lo_hi_lo_3};
  wire [63:0]        regroupV0_lo_hi_hi_hi_lo_3 = {regroupV0_lo_hi_hi_hi_lo_hi_3, regroupV0_lo_hi_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_2 = {regroupV0_lo[3867:3864], regroupV0_lo[3851:3848]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_2 = {regroupV0_lo[3899:3896], regroupV0_lo[3883:3880]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_lo_lo_3 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_2, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_2 = {regroupV0_lo[3931:3928], regroupV0_lo[3915:3912]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_2 = {regroupV0_lo[3963:3960], regroupV0_lo[3947:3944]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_lo_hi_3 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_2, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_2};
  wire [31:0]        regroupV0_lo_hi_hi_hi_hi_lo_3 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_3, regroupV0_lo_hi_hi_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_2 = {regroupV0_lo[3995:3992], regroupV0_lo[3979:3976]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_2 = {regroupV0_lo[4027:4024], regroupV0_lo[4011:4008]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_hi_lo_3 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_2, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_2 = {regroupV0_lo[4059:4056], regroupV0_lo[4043:4040]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_2 = {regroupV0_lo[4091:4088], regroupV0_lo[4075:4072]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_hi_hi_3 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_2, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_2};
  wire [31:0]        regroupV0_lo_hi_hi_hi_hi_hi_3 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_3, regroupV0_lo_hi_hi_hi_hi_hi_lo_3};
  wire [63:0]        regroupV0_lo_hi_hi_hi_hi_3 = {regroupV0_lo_hi_hi_hi_hi_hi_3, regroupV0_lo_hi_hi_hi_hi_lo_3};
  wire [127:0]       regroupV0_lo_hi_hi_hi_3 = {regroupV0_lo_hi_hi_hi_hi_3, regroupV0_lo_hi_hi_hi_lo_3};
  wire [255:0]       regroupV0_lo_hi_hi_3 = {regroupV0_lo_hi_hi_hi_3, regroupV0_lo_hi_hi_lo_3};
  wire [511:0]       regroupV0_lo_hi_3 = {regroupV0_lo_hi_hi_3, regroupV0_lo_hi_lo_3};
  wire [1023:0]      regroupV0_lo_3 = {regroupV0_lo_hi_3, regroupV0_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_2 = {regroupV0_hi[27:24], regroupV0_hi[11:8]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_2 = {regroupV0_hi[59:56], regroupV0_hi[43:40]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_lo_lo_3 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_2 = {regroupV0_hi[91:88], regroupV0_hi[75:72]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_2 = {regroupV0_hi[123:120], regroupV0_hi[107:104]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_lo_hi_3 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_2, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_2};
  wire [31:0]        regroupV0_hi_lo_lo_lo_lo_lo_3 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_2 = {regroupV0_hi[155:152], regroupV0_hi[139:136]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_2 = {regroupV0_hi[187:184], regroupV0_hi[171:168]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_hi_lo_3 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_2, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_2 = {regroupV0_hi[219:216], regroupV0_hi[203:200]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_2 = {regroupV0_hi[251:248], regroupV0_hi[235:232]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_hi_hi_3 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_2, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_2};
  wire [31:0]        regroupV0_hi_lo_lo_lo_lo_hi_3 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_3, regroupV0_hi_lo_lo_lo_lo_hi_lo_3};
  wire [63:0]        regroupV0_hi_lo_lo_lo_lo_3 = {regroupV0_hi_lo_lo_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_2 = {regroupV0_hi[283:280], regroupV0_hi[267:264]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_2 = {regroupV0_hi[315:312], regroupV0_hi[299:296]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_lo_lo_3 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_2 = {regroupV0_hi[347:344], regroupV0_hi[331:328]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_2 = {regroupV0_hi[379:376], regroupV0_hi[363:360]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_lo_hi_3 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_2, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_2};
  wire [31:0]        regroupV0_hi_lo_lo_lo_hi_lo_3 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_3, regroupV0_hi_lo_lo_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_2 = {regroupV0_hi[411:408], regroupV0_hi[395:392]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_2 = {regroupV0_hi[443:440], regroupV0_hi[427:424]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_hi_lo_3 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_2, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_2 = {regroupV0_hi[475:472], regroupV0_hi[459:456]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_2 = {regroupV0_hi[507:504], regroupV0_hi[491:488]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_hi_hi_3 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_2, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_2};
  wire [31:0]        regroupV0_hi_lo_lo_lo_hi_hi_3 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_3, regroupV0_hi_lo_lo_lo_hi_hi_lo_3};
  wire [63:0]        regroupV0_hi_lo_lo_lo_hi_3 = {regroupV0_hi_lo_lo_lo_hi_hi_3, regroupV0_hi_lo_lo_lo_hi_lo_3};
  wire [127:0]       regroupV0_hi_lo_lo_lo_3 = {regroupV0_hi_lo_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_2 = {regroupV0_hi[539:536], regroupV0_hi[523:520]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_2 = {regroupV0_hi[571:568], regroupV0_hi[555:552]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_lo_lo_3 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_2, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_2 = {regroupV0_hi[603:600], regroupV0_hi[587:584]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_2 = {regroupV0_hi[635:632], regroupV0_hi[619:616]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_lo_hi_3 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_2, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_2};
  wire [31:0]        regroupV0_hi_lo_lo_hi_lo_lo_3 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_3, regroupV0_hi_lo_lo_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_2 = {regroupV0_hi[667:664], regroupV0_hi[651:648]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_2 = {regroupV0_hi[699:696], regroupV0_hi[683:680]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_hi_lo_3 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_2, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_2 = {regroupV0_hi[731:728], regroupV0_hi[715:712]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_2 = {regroupV0_hi[763:760], regroupV0_hi[747:744]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_hi_hi_3 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_2, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_2};
  wire [31:0]        regroupV0_hi_lo_lo_hi_lo_hi_3 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_3, regroupV0_hi_lo_lo_hi_lo_hi_lo_3};
  wire [63:0]        regroupV0_hi_lo_lo_hi_lo_3 = {regroupV0_hi_lo_lo_hi_lo_hi_3, regroupV0_hi_lo_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_2 = {regroupV0_hi[795:792], regroupV0_hi[779:776]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_2 = {regroupV0_hi[827:824], regroupV0_hi[811:808]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_lo_lo_3 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_2, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_2 = {regroupV0_hi[859:856], regroupV0_hi[843:840]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_2 = {regroupV0_hi[891:888], regroupV0_hi[875:872]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_lo_hi_3 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_2, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_2};
  wire [31:0]        regroupV0_hi_lo_lo_hi_hi_lo_3 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_3, regroupV0_hi_lo_lo_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_2 = {regroupV0_hi[923:920], regroupV0_hi[907:904]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_2 = {regroupV0_hi[955:952], regroupV0_hi[939:936]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_hi_lo_3 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_2, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_2 = {regroupV0_hi[987:984], regroupV0_hi[971:968]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_2 = {regroupV0_hi[1019:1016], regroupV0_hi[1003:1000]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_hi_hi_3 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_2, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_2};
  wire [31:0]        regroupV0_hi_lo_lo_hi_hi_hi_3 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_3, regroupV0_hi_lo_lo_hi_hi_hi_lo_3};
  wire [63:0]        regroupV0_hi_lo_lo_hi_hi_3 = {regroupV0_hi_lo_lo_hi_hi_hi_3, regroupV0_hi_lo_lo_hi_hi_lo_3};
  wire [127:0]       regroupV0_hi_lo_lo_hi_3 = {regroupV0_hi_lo_lo_hi_hi_3, regroupV0_hi_lo_lo_hi_lo_3};
  wire [255:0]       regroupV0_hi_lo_lo_3 = {regroupV0_hi_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_2 = {regroupV0_hi[1051:1048], regroupV0_hi[1035:1032]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_2 = {regroupV0_hi[1083:1080], regroupV0_hi[1067:1064]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_lo_lo_3 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_2, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_2 = {regroupV0_hi[1115:1112], regroupV0_hi[1099:1096]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_2 = {regroupV0_hi[1147:1144], regroupV0_hi[1131:1128]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_lo_hi_3 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_2, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_2};
  wire [31:0]        regroupV0_hi_lo_hi_lo_lo_lo_3 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_3, regroupV0_hi_lo_hi_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_2 = {regroupV0_hi[1179:1176], regroupV0_hi[1163:1160]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_2 = {regroupV0_hi[1211:1208], regroupV0_hi[1195:1192]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_hi_lo_3 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_2, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_2 = {regroupV0_hi[1243:1240], regroupV0_hi[1227:1224]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_2 = {regroupV0_hi[1275:1272], regroupV0_hi[1259:1256]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_hi_hi_3 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_2, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_2};
  wire [31:0]        regroupV0_hi_lo_hi_lo_lo_hi_3 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_3, regroupV0_hi_lo_hi_lo_lo_hi_lo_3};
  wire [63:0]        regroupV0_hi_lo_hi_lo_lo_3 = {regroupV0_hi_lo_hi_lo_lo_hi_3, regroupV0_hi_lo_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_2 = {regroupV0_hi[1307:1304], regroupV0_hi[1291:1288]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_2 = {regroupV0_hi[1339:1336], regroupV0_hi[1323:1320]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_lo_lo_3 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_2, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_2 = {regroupV0_hi[1371:1368], regroupV0_hi[1355:1352]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_2 = {regroupV0_hi[1403:1400], regroupV0_hi[1387:1384]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_lo_hi_3 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_2, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_2};
  wire [31:0]        regroupV0_hi_lo_hi_lo_hi_lo_3 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_3, regroupV0_hi_lo_hi_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_2 = {regroupV0_hi[1435:1432], regroupV0_hi[1419:1416]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_2 = {regroupV0_hi[1467:1464], regroupV0_hi[1451:1448]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_hi_lo_3 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_2, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_2 = {regroupV0_hi[1499:1496], regroupV0_hi[1483:1480]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_2 = {regroupV0_hi[1531:1528], regroupV0_hi[1515:1512]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_hi_hi_3 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_2, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_2};
  wire [31:0]        regroupV0_hi_lo_hi_lo_hi_hi_3 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_3, regroupV0_hi_lo_hi_lo_hi_hi_lo_3};
  wire [63:0]        regroupV0_hi_lo_hi_lo_hi_3 = {regroupV0_hi_lo_hi_lo_hi_hi_3, regroupV0_hi_lo_hi_lo_hi_lo_3};
  wire [127:0]       regroupV0_hi_lo_hi_lo_3 = {regroupV0_hi_lo_hi_lo_hi_3, regroupV0_hi_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_2 = {regroupV0_hi[1563:1560], regroupV0_hi[1547:1544]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_2 = {regroupV0_hi[1595:1592], regroupV0_hi[1579:1576]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_lo_lo_3 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_2, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_2 = {regroupV0_hi[1627:1624], regroupV0_hi[1611:1608]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_2 = {regroupV0_hi[1659:1656], regroupV0_hi[1643:1640]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_lo_hi_3 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_2, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_2};
  wire [31:0]        regroupV0_hi_lo_hi_hi_lo_lo_3 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_3, regroupV0_hi_lo_hi_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_2 = {regroupV0_hi[1691:1688], regroupV0_hi[1675:1672]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_2 = {regroupV0_hi[1723:1720], regroupV0_hi[1707:1704]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_hi_lo_3 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_2, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_2 = {regroupV0_hi[1755:1752], regroupV0_hi[1739:1736]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_2 = {regroupV0_hi[1787:1784], regroupV0_hi[1771:1768]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_hi_hi_3 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_2, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_2};
  wire [31:0]        regroupV0_hi_lo_hi_hi_lo_hi_3 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_3, regroupV0_hi_lo_hi_hi_lo_hi_lo_3};
  wire [63:0]        regroupV0_hi_lo_hi_hi_lo_3 = {regroupV0_hi_lo_hi_hi_lo_hi_3, regroupV0_hi_lo_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_2 = {regroupV0_hi[1819:1816], regroupV0_hi[1803:1800]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_2 = {regroupV0_hi[1851:1848], regroupV0_hi[1835:1832]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_lo_lo_3 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_2, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_2 = {regroupV0_hi[1883:1880], regroupV0_hi[1867:1864]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_2 = {regroupV0_hi[1915:1912], regroupV0_hi[1899:1896]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_lo_hi_3 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_2, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_2};
  wire [31:0]        regroupV0_hi_lo_hi_hi_hi_lo_3 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_3, regroupV0_hi_lo_hi_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_2 = {regroupV0_hi[1947:1944], regroupV0_hi[1931:1928]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_2 = {regroupV0_hi[1979:1976], regroupV0_hi[1963:1960]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_hi_lo_3 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_2, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_2 = {regroupV0_hi[2011:2008], regroupV0_hi[1995:1992]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_2 = {regroupV0_hi[2043:2040], regroupV0_hi[2027:2024]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_hi_hi_3 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_2, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_2};
  wire [31:0]        regroupV0_hi_lo_hi_hi_hi_hi_3 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_3, regroupV0_hi_lo_hi_hi_hi_hi_lo_3};
  wire [63:0]        regroupV0_hi_lo_hi_hi_hi_3 = {regroupV0_hi_lo_hi_hi_hi_hi_3, regroupV0_hi_lo_hi_hi_hi_lo_3};
  wire [127:0]       regroupV0_hi_lo_hi_hi_3 = {regroupV0_hi_lo_hi_hi_hi_3, regroupV0_hi_lo_hi_hi_lo_3};
  wire [255:0]       regroupV0_hi_lo_hi_3 = {regroupV0_hi_lo_hi_hi_3, regroupV0_hi_lo_hi_lo_3};
  wire [511:0]       regroupV0_hi_lo_3 = {regroupV0_hi_lo_hi_3, regroupV0_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_2 = {regroupV0_hi[2075:2072], regroupV0_hi[2059:2056]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_2 = {regroupV0_hi[2107:2104], regroupV0_hi[2091:2088]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_lo_lo_3 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_2, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_2 = {regroupV0_hi[2139:2136], regroupV0_hi[2123:2120]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_2 = {regroupV0_hi[2171:2168], regroupV0_hi[2155:2152]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_lo_hi_3 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_2, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_2};
  wire [31:0]        regroupV0_hi_hi_lo_lo_lo_lo_3 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_3, regroupV0_hi_hi_lo_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_2 = {regroupV0_hi[2203:2200], regroupV0_hi[2187:2184]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_2 = {regroupV0_hi[2235:2232], regroupV0_hi[2219:2216]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_hi_lo_3 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_2, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_2 = {regroupV0_hi[2267:2264], regroupV0_hi[2251:2248]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_2 = {regroupV0_hi[2299:2296], regroupV0_hi[2283:2280]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_hi_hi_3 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_2, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_2};
  wire [31:0]        regroupV0_hi_hi_lo_lo_lo_hi_3 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_3, regroupV0_hi_hi_lo_lo_lo_hi_lo_3};
  wire [63:0]        regroupV0_hi_hi_lo_lo_lo_3 = {regroupV0_hi_hi_lo_lo_lo_hi_3, regroupV0_hi_hi_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_2 = {regroupV0_hi[2331:2328], regroupV0_hi[2315:2312]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_2 = {regroupV0_hi[2363:2360], regroupV0_hi[2347:2344]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_lo_lo_3 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_2, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_2 = {regroupV0_hi[2395:2392], regroupV0_hi[2379:2376]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_2 = {regroupV0_hi[2427:2424], regroupV0_hi[2411:2408]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_lo_hi_3 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_2, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_2};
  wire [31:0]        regroupV0_hi_hi_lo_lo_hi_lo_3 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_3, regroupV0_hi_hi_lo_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_2 = {regroupV0_hi[2459:2456], regroupV0_hi[2443:2440]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_2 = {regroupV0_hi[2491:2488], regroupV0_hi[2475:2472]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_hi_lo_3 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_2, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_2 = {regroupV0_hi[2523:2520], regroupV0_hi[2507:2504]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_2 = {regroupV0_hi[2555:2552], regroupV0_hi[2539:2536]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_hi_hi_3 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_2, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_2};
  wire [31:0]        regroupV0_hi_hi_lo_lo_hi_hi_3 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_3, regroupV0_hi_hi_lo_lo_hi_hi_lo_3};
  wire [63:0]        regroupV0_hi_hi_lo_lo_hi_3 = {regroupV0_hi_hi_lo_lo_hi_hi_3, regroupV0_hi_hi_lo_lo_hi_lo_3};
  wire [127:0]       regroupV0_hi_hi_lo_lo_3 = {regroupV0_hi_hi_lo_lo_hi_3, regroupV0_hi_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_2 = {regroupV0_hi[2587:2584], regroupV0_hi[2571:2568]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_2 = {regroupV0_hi[2619:2616], regroupV0_hi[2603:2600]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_lo_lo_3 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_2, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_2 = {regroupV0_hi[2651:2648], regroupV0_hi[2635:2632]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_2 = {regroupV0_hi[2683:2680], regroupV0_hi[2667:2664]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_lo_hi_3 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_2, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_2};
  wire [31:0]        regroupV0_hi_hi_lo_hi_lo_lo_3 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_3, regroupV0_hi_hi_lo_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_2 = {regroupV0_hi[2715:2712], regroupV0_hi[2699:2696]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_2 = {regroupV0_hi[2747:2744], regroupV0_hi[2731:2728]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_hi_lo_3 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_2, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_2 = {regroupV0_hi[2779:2776], regroupV0_hi[2763:2760]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_2 = {regroupV0_hi[2811:2808], regroupV0_hi[2795:2792]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_hi_hi_3 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_2, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_2};
  wire [31:0]        regroupV0_hi_hi_lo_hi_lo_hi_3 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_3, regroupV0_hi_hi_lo_hi_lo_hi_lo_3};
  wire [63:0]        regroupV0_hi_hi_lo_hi_lo_3 = {regroupV0_hi_hi_lo_hi_lo_hi_3, regroupV0_hi_hi_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_2 = {regroupV0_hi[2843:2840], regroupV0_hi[2827:2824]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_2 = {regroupV0_hi[2875:2872], regroupV0_hi[2859:2856]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_lo_lo_3 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_2, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_2 = {regroupV0_hi[2907:2904], regroupV0_hi[2891:2888]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_2 = {regroupV0_hi[2939:2936], regroupV0_hi[2923:2920]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_lo_hi_3 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_2, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_2};
  wire [31:0]        regroupV0_hi_hi_lo_hi_hi_lo_3 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_3, regroupV0_hi_hi_lo_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_2 = {regroupV0_hi[2971:2968], regroupV0_hi[2955:2952]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_2 = {regroupV0_hi[3003:3000], regroupV0_hi[2987:2984]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_hi_lo_3 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_2, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_2 = {regroupV0_hi[3035:3032], regroupV0_hi[3019:3016]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_2 = {regroupV0_hi[3067:3064], regroupV0_hi[3051:3048]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_hi_hi_3 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_2, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_2};
  wire [31:0]        regroupV0_hi_hi_lo_hi_hi_hi_3 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_3, regroupV0_hi_hi_lo_hi_hi_hi_lo_3};
  wire [63:0]        regroupV0_hi_hi_lo_hi_hi_3 = {regroupV0_hi_hi_lo_hi_hi_hi_3, regroupV0_hi_hi_lo_hi_hi_lo_3};
  wire [127:0]       regroupV0_hi_hi_lo_hi_3 = {regroupV0_hi_hi_lo_hi_hi_3, regroupV0_hi_hi_lo_hi_lo_3};
  wire [255:0]       regroupV0_hi_hi_lo_3 = {regroupV0_hi_hi_lo_hi_3, regroupV0_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_2 = {regroupV0_hi[3099:3096], regroupV0_hi[3083:3080]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_2 = {regroupV0_hi[3131:3128], regroupV0_hi[3115:3112]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_lo_lo_3 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_2, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_2 = {regroupV0_hi[3163:3160], regroupV0_hi[3147:3144]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_2 = {regroupV0_hi[3195:3192], regroupV0_hi[3179:3176]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_lo_hi_3 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_2, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_2};
  wire [31:0]        regroupV0_hi_hi_hi_lo_lo_lo_3 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_3, regroupV0_hi_hi_hi_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_2 = {regroupV0_hi[3227:3224], regroupV0_hi[3211:3208]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_2 = {regroupV0_hi[3259:3256], regroupV0_hi[3243:3240]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_hi_lo_3 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_2, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_2 = {regroupV0_hi[3291:3288], regroupV0_hi[3275:3272]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_2 = {regroupV0_hi[3323:3320], regroupV0_hi[3307:3304]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_hi_hi_3 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_2, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_2};
  wire [31:0]        regroupV0_hi_hi_hi_lo_lo_hi_3 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_3, regroupV0_hi_hi_hi_lo_lo_hi_lo_3};
  wire [63:0]        regroupV0_hi_hi_hi_lo_lo_3 = {regroupV0_hi_hi_hi_lo_lo_hi_3, regroupV0_hi_hi_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_2 = {regroupV0_hi[3355:3352], regroupV0_hi[3339:3336]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_2 = {regroupV0_hi[3387:3384], regroupV0_hi[3371:3368]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_lo_lo_3 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_2, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_2 = {regroupV0_hi[3419:3416], regroupV0_hi[3403:3400]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_2 = {regroupV0_hi[3451:3448], regroupV0_hi[3435:3432]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_lo_hi_3 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_2, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_2};
  wire [31:0]        regroupV0_hi_hi_hi_lo_hi_lo_3 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_3, regroupV0_hi_hi_hi_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_2 = {regroupV0_hi[3483:3480], regroupV0_hi[3467:3464]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_2 = {regroupV0_hi[3515:3512], regroupV0_hi[3499:3496]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_hi_lo_3 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_2, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_2 = {regroupV0_hi[3547:3544], regroupV0_hi[3531:3528]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_2 = {regroupV0_hi[3579:3576], regroupV0_hi[3563:3560]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_hi_hi_3 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_2};
  wire [31:0]        regroupV0_hi_hi_hi_lo_hi_hi_3 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_3, regroupV0_hi_hi_hi_lo_hi_hi_lo_3};
  wire [63:0]        regroupV0_hi_hi_hi_lo_hi_3 = {regroupV0_hi_hi_hi_lo_hi_hi_3, regroupV0_hi_hi_hi_lo_hi_lo_3};
  wire [127:0]       regroupV0_hi_hi_hi_lo_3 = {regroupV0_hi_hi_hi_lo_hi_3, regroupV0_hi_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_2 = {regroupV0_hi[3611:3608], regroupV0_hi[3595:3592]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_2 = {regroupV0_hi[3643:3640], regroupV0_hi[3627:3624]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_lo_lo_3 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_2, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_2 = {regroupV0_hi[3675:3672], regroupV0_hi[3659:3656]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_2 = {regroupV0_hi[3707:3704], regroupV0_hi[3691:3688]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_lo_hi_3 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_2, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_2};
  wire [31:0]        regroupV0_hi_hi_hi_hi_lo_lo_3 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_3, regroupV0_hi_hi_hi_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_2 = {regroupV0_hi[3739:3736], regroupV0_hi[3723:3720]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_2 = {regroupV0_hi[3771:3768], regroupV0_hi[3755:3752]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_hi_lo_3 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_2, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_2 = {regroupV0_hi[3803:3800], regroupV0_hi[3787:3784]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_2 = {regroupV0_hi[3835:3832], regroupV0_hi[3819:3816]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_hi_hi_3 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_2, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_2};
  wire [31:0]        regroupV0_hi_hi_hi_hi_lo_hi_3 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_3, regroupV0_hi_hi_hi_hi_lo_hi_lo_3};
  wire [63:0]        regroupV0_hi_hi_hi_hi_lo_3 = {regroupV0_hi_hi_hi_hi_lo_hi_3, regroupV0_hi_hi_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_2 = {regroupV0_hi[3867:3864], regroupV0_hi[3851:3848]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_2 = {regroupV0_hi[3899:3896], regroupV0_hi[3883:3880]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_lo_lo_3 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_2, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_2 = {regroupV0_hi[3931:3928], regroupV0_hi[3915:3912]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_2 = {regroupV0_hi[3963:3960], regroupV0_hi[3947:3944]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_lo_hi_3 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_2, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_2};
  wire [31:0]        regroupV0_hi_hi_hi_hi_hi_lo_3 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_3, regroupV0_hi_hi_hi_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_2 = {regroupV0_hi[3995:3992], regroupV0_hi[3979:3976]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_2 = {regroupV0_hi[4027:4024], regroupV0_hi[4011:4008]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_hi_lo_3 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_2, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_2 = {regroupV0_hi[4059:4056], regroupV0_hi[4043:4040]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_2 = {regroupV0_hi[4091:4088], regroupV0_hi[4075:4072]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_hi_hi_3 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_2};
  wire [31:0]        regroupV0_hi_hi_hi_hi_hi_hi_3 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_hi_hi_hi_lo_3};
  wire [63:0]        regroupV0_hi_hi_hi_hi_hi_3 = {regroupV0_hi_hi_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_hi_hi_lo_3};
  wire [127:0]       regroupV0_hi_hi_hi_hi_3 = {regroupV0_hi_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_hi_lo_3};
  wire [255:0]       regroupV0_hi_hi_hi_3 = {regroupV0_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_lo_3};
  wire [511:0]       regroupV0_hi_hi_3 = {regroupV0_hi_hi_hi_3, regroupV0_hi_hi_lo_3};
  wire [1023:0]      regroupV0_hi_3 = {regroupV0_hi_hi_3, regroupV0_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_3 = {regroupV0_lo[31:28], regroupV0_lo[15:12]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_3 = {regroupV0_lo[63:60], regroupV0_lo[47:44]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_lo_lo_4 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_3 = {regroupV0_lo[95:92], regroupV0_lo[79:76]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_3 = {regroupV0_lo[127:124], regroupV0_lo[111:108]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_lo_hi_4 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_3, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_3};
  wire [31:0]        regroupV0_lo_lo_lo_lo_lo_lo_4 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_4, regroupV0_lo_lo_lo_lo_lo_lo_lo_4};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_3 = {regroupV0_lo[159:156], regroupV0_lo[143:140]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_3 = {regroupV0_lo[191:188], regroupV0_lo[175:172]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_hi_lo_4 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_3, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_3 = {regroupV0_lo[223:220], regroupV0_lo[207:204]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_3 = {regroupV0_lo[255:252], regroupV0_lo[239:236]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_hi_hi_4 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_3, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_3};
  wire [31:0]        regroupV0_lo_lo_lo_lo_lo_hi_4 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_4, regroupV0_lo_lo_lo_lo_lo_hi_lo_4};
  wire [63:0]        regroupV0_lo_lo_lo_lo_lo_4 = {regroupV0_lo_lo_lo_lo_lo_hi_4, regroupV0_lo_lo_lo_lo_lo_lo_4};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_3 = {regroupV0_lo[287:284], regroupV0_lo[271:268]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_3 = {regroupV0_lo[319:316], regroupV0_lo[303:300]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_lo_lo_4 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_3 = {regroupV0_lo[351:348], regroupV0_lo[335:332]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_3 = {regroupV0_lo[383:380], regroupV0_lo[367:364]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_lo_hi_4 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_3, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_3};
  wire [31:0]        regroupV0_lo_lo_lo_lo_hi_lo_4 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_4, regroupV0_lo_lo_lo_lo_hi_lo_lo_4};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_3 = {regroupV0_lo[415:412], regroupV0_lo[399:396]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_3 = {regroupV0_lo[447:444], regroupV0_lo[431:428]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_hi_lo_4 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_3, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_3 = {regroupV0_lo[479:476], regroupV0_lo[463:460]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_3 = {regroupV0_lo[511:508], regroupV0_lo[495:492]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_hi_hi_4 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_3, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_3};
  wire [31:0]        regroupV0_lo_lo_lo_lo_hi_hi_4 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_4, regroupV0_lo_lo_lo_lo_hi_hi_lo_4};
  wire [63:0]        regroupV0_lo_lo_lo_lo_hi_4 = {regroupV0_lo_lo_lo_lo_hi_hi_4, regroupV0_lo_lo_lo_lo_hi_lo_4};
  wire [127:0]       regroupV0_lo_lo_lo_lo_4 = {regroupV0_lo_lo_lo_lo_hi_4, regroupV0_lo_lo_lo_lo_lo_4};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_3 = {regroupV0_lo[543:540], regroupV0_lo[527:524]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_3 = {regroupV0_lo[575:572], regroupV0_lo[559:556]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_lo_lo_4 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_3 = {regroupV0_lo[607:604], regroupV0_lo[591:588]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_3 = {regroupV0_lo[639:636], regroupV0_lo[623:620]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_lo_hi_4 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_3, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_3};
  wire [31:0]        regroupV0_lo_lo_lo_hi_lo_lo_4 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_4, regroupV0_lo_lo_lo_hi_lo_lo_lo_4};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_3 = {regroupV0_lo[671:668], regroupV0_lo[655:652]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_3 = {regroupV0_lo[703:700], regroupV0_lo[687:684]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_hi_lo_4 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_3, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_3 = {regroupV0_lo[735:732], regroupV0_lo[719:716]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_3 = {regroupV0_lo[767:764], regroupV0_lo[751:748]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_hi_hi_4 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_3, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_3};
  wire [31:0]        regroupV0_lo_lo_lo_hi_lo_hi_4 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_4, regroupV0_lo_lo_lo_hi_lo_hi_lo_4};
  wire [63:0]        regroupV0_lo_lo_lo_hi_lo_4 = {regroupV0_lo_lo_lo_hi_lo_hi_4, regroupV0_lo_lo_lo_hi_lo_lo_4};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_3 = {regroupV0_lo[799:796], regroupV0_lo[783:780]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_3 = {regroupV0_lo[831:828], regroupV0_lo[815:812]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_lo_lo_4 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_3, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_3 = {regroupV0_lo[863:860], regroupV0_lo[847:844]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_3 = {regroupV0_lo[895:892], regroupV0_lo[879:876]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_lo_hi_4 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_3, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_3};
  wire [31:0]        regroupV0_lo_lo_lo_hi_hi_lo_4 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_4, regroupV0_lo_lo_lo_hi_hi_lo_lo_4};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_3 = {regroupV0_lo[927:924], regroupV0_lo[911:908]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_3 = {regroupV0_lo[959:956], regroupV0_lo[943:940]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_hi_lo_4 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_3, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_3 = {regroupV0_lo[991:988], regroupV0_lo[975:972]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_3 = {regroupV0_lo[1023:1020], regroupV0_lo[1007:1004]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_hi_hi_4 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_3, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_3};
  wire [31:0]        regroupV0_lo_lo_lo_hi_hi_hi_4 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_4, regroupV0_lo_lo_lo_hi_hi_hi_lo_4};
  wire [63:0]        regroupV0_lo_lo_lo_hi_hi_4 = {regroupV0_lo_lo_lo_hi_hi_hi_4, regroupV0_lo_lo_lo_hi_hi_lo_4};
  wire [127:0]       regroupV0_lo_lo_lo_hi_4 = {regroupV0_lo_lo_lo_hi_hi_4, regroupV0_lo_lo_lo_hi_lo_4};
  wire [255:0]       regroupV0_lo_lo_lo_4 = {regroupV0_lo_lo_lo_hi_4, regroupV0_lo_lo_lo_lo_4};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_3 = {regroupV0_lo[1055:1052], regroupV0_lo[1039:1036]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_3 = {regroupV0_lo[1087:1084], regroupV0_lo[1071:1068]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_lo_lo_4 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_3, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_3 = {regroupV0_lo[1119:1116], regroupV0_lo[1103:1100]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_3 = {regroupV0_lo[1151:1148], regroupV0_lo[1135:1132]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_lo_hi_4 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_3, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_3};
  wire [31:0]        regroupV0_lo_lo_hi_lo_lo_lo_4 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_4, regroupV0_lo_lo_hi_lo_lo_lo_lo_4};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_3 = {regroupV0_lo[1183:1180], regroupV0_lo[1167:1164]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_3 = {regroupV0_lo[1215:1212], regroupV0_lo[1199:1196]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_hi_lo_4 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_3, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_3 = {regroupV0_lo[1247:1244], regroupV0_lo[1231:1228]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_3 = {regroupV0_lo[1279:1276], regroupV0_lo[1263:1260]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_hi_hi_4 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_3, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_3};
  wire [31:0]        regroupV0_lo_lo_hi_lo_lo_hi_4 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_4, regroupV0_lo_lo_hi_lo_lo_hi_lo_4};
  wire [63:0]        regroupV0_lo_lo_hi_lo_lo_4 = {regroupV0_lo_lo_hi_lo_lo_hi_4, regroupV0_lo_lo_hi_lo_lo_lo_4};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_3 = {regroupV0_lo[1311:1308], regroupV0_lo[1295:1292]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_3 = {regroupV0_lo[1343:1340], regroupV0_lo[1327:1324]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_lo_lo_4 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_3, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_3 = {regroupV0_lo[1375:1372], regroupV0_lo[1359:1356]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_3 = {regroupV0_lo[1407:1404], regroupV0_lo[1391:1388]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_lo_hi_4 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_3, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_3};
  wire [31:0]        regroupV0_lo_lo_hi_lo_hi_lo_4 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_4, regroupV0_lo_lo_hi_lo_hi_lo_lo_4};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_3 = {regroupV0_lo[1439:1436], regroupV0_lo[1423:1420]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_3 = {regroupV0_lo[1471:1468], regroupV0_lo[1455:1452]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_hi_lo_4 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_3, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_3 = {regroupV0_lo[1503:1500], regroupV0_lo[1487:1484]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_3 = {regroupV0_lo[1535:1532], regroupV0_lo[1519:1516]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_hi_hi_4 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_3, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_3};
  wire [31:0]        regroupV0_lo_lo_hi_lo_hi_hi_4 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_4, regroupV0_lo_lo_hi_lo_hi_hi_lo_4};
  wire [63:0]        regroupV0_lo_lo_hi_lo_hi_4 = {regroupV0_lo_lo_hi_lo_hi_hi_4, regroupV0_lo_lo_hi_lo_hi_lo_4};
  wire [127:0]       regroupV0_lo_lo_hi_lo_4 = {regroupV0_lo_lo_hi_lo_hi_4, regroupV0_lo_lo_hi_lo_lo_4};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_3 = {regroupV0_lo[1567:1564], regroupV0_lo[1551:1548]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_3 = {regroupV0_lo[1599:1596], regroupV0_lo[1583:1580]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_lo_lo_4 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_3, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_3 = {regroupV0_lo[1631:1628], regroupV0_lo[1615:1612]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_3 = {regroupV0_lo[1663:1660], regroupV0_lo[1647:1644]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_lo_hi_4 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_3, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_3};
  wire [31:0]        regroupV0_lo_lo_hi_hi_lo_lo_4 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_4, regroupV0_lo_lo_hi_hi_lo_lo_lo_4};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_3 = {regroupV0_lo[1695:1692], regroupV0_lo[1679:1676]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_3 = {regroupV0_lo[1727:1724], regroupV0_lo[1711:1708]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_hi_lo_4 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_3, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_3 = {regroupV0_lo[1759:1756], regroupV0_lo[1743:1740]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_3 = {regroupV0_lo[1791:1788], regroupV0_lo[1775:1772]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_hi_hi_4 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_3, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_3};
  wire [31:0]        regroupV0_lo_lo_hi_hi_lo_hi_4 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_4, regroupV0_lo_lo_hi_hi_lo_hi_lo_4};
  wire [63:0]        regroupV0_lo_lo_hi_hi_lo_4 = {regroupV0_lo_lo_hi_hi_lo_hi_4, regroupV0_lo_lo_hi_hi_lo_lo_4};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_3 = {regroupV0_lo[1823:1820], regroupV0_lo[1807:1804]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_3 = {regroupV0_lo[1855:1852], regroupV0_lo[1839:1836]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_lo_lo_4 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_3, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_3 = {regroupV0_lo[1887:1884], regroupV0_lo[1871:1868]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_3 = {regroupV0_lo[1919:1916], regroupV0_lo[1903:1900]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_lo_hi_4 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_3, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_3};
  wire [31:0]        regroupV0_lo_lo_hi_hi_hi_lo_4 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_4, regroupV0_lo_lo_hi_hi_hi_lo_lo_4};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_3 = {regroupV0_lo[1951:1948], regroupV0_lo[1935:1932]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_3 = {regroupV0_lo[1983:1980], regroupV0_lo[1967:1964]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_hi_lo_4 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_3, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_3 = {regroupV0_lo[2015:2012], regroupV0_lo[1999:1996]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_3 = {regroupV0_lo[2047:2044], regroupV0_lo[2031:2028]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_hi_hi_4 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_3, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_3};
  wire [31:0]        regroupV0_lo_lo_hi_hi_hi_hi_4 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_4, regroupV0_lo_lo_hi_hi_hi_hi_lo_4};
  wire [63:0]        regroupV0_lo_lo_hi_hi_hi_4 = {regroupV0_lo_lo_hi_hi_hi_hi_4, regroupV0_lo_lo_hi_hi_hi_lo_4};
  wire [127:0]       regroupV0_lo_lo_hi_hi_4 = {regroupV0_lo_lo_hi_hi_hi_4, regroupV0_lo_lo_hi_hi_lo_4};
  wire [255:0]       regroupV0_lo_lo_hi_4 = {regroupV0_lo_lo_hi_hi_4, regroupV0_lo_lo_hi_lo_4};
  wire [511:0]       regroupV0_lo_lo_4 = {regroupV0_lo_lo_hi_4, regroupV0_lo_lo_lo_4};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_3 = {regroupV0_lo[2079:2076], regroupV0_lo[2063:2060]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_3 = {regroupV0_lo[2111:2108], regroupV0_lo[2095:2092]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_lo_lo_4 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_3, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_3 = {regroupV0_lo[2143:2140], regroupV0_lo[2127:2124]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_3 = {regroupV0_lo[2175:2172], regroupV0_lo[2159:2156]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_lo_hi_4 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_3, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_3};
  wire [31:0]        regroupV0_lo_hi_lo_lo_lo_lo_4 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_4, regroupV0_lo_hi_lo_lo_lo_lo_lo_4};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_3 = {regroupV0_lo[2207:2204], regroupV0_lo[2191:2188]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_3 = {regroupV0_lo[2239:2236], regroupV0_lo[2223:2220]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_hi_lo_4 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_3, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_3 = {regroupV0_lo[2271:2268], regroupV0_lo[2255:2252]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_3 = {regroupV0_lo[2303:2300], regroupV0_lo[2287:2284]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_hi_hi_4 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_3, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_3};
  wire [31:0]        regroupV0_lo_hi_lo_lo_lo_hi_4 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_4, regroupV0_lo_hi_lo_lo_lo_hi_lo_4};
  wire [63:0]        regroupV0_lo_hi_lo_lo_lo_4 = {regroupV0_lo_hi_lo_lo_lo_hi_4, regroupV0_lo_hi_lo_lo_lo_lo_4};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_3 = {regroupV0_lo[2335:2332], regroupV0_lo[2319:2316]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_3 = {regroupV0_lo[2367:2364], regroupV0_lo[2351:2348]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_lo_lo_4 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_3, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_3 = {regroupV0_lo[2399:2396], regroupV0_lo[2383:2380]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_3 = {regroupV0_lo[2431:2428], regroupV0_lo[2415:2412]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_lo_hi_4 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_3, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_3};
  wire [31:0]        regroupV0_lo_hi_lo_lo_hi_lo_4 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_4, regroupV0_lo_hi_lo_lo_hi_lo_lo_4};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_3 = {regroupV0_lo[2463:2460], regroupV0_lo[2447:2444]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_3 = {regroupV0_lo[2495:2492], regroupV0_lo[2479:2476]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_hi_lo_4 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_3, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_3 = {regroupV0_lo[2527:2524], regroupV0_lo[2511:2508]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_3 = {regroupV0_lo[2559:2556], regroupV0_lo[2543:2540]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_hi_hi_4 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_3, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_3};
  wire [31:0]        regroupV0_lo_hi_lo_lo_hi_hi_4 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_4, regroupV0_lo_hi_lo_lo_hi_hi_lo_4};
  wire [63:0]        regroupV0_lo_hi_lo_lo_hi_4 = {regroupV0_lo_hi_lo_lo_hi_hi_4, regroupV0_lo_hi_lo_lo_hi_lo_4};
  wire [127:0]       regroupV0_lo_hi_lo_lo_4 = {regroupV0_lo_hi_lo_lo_hi_4, regroupV0_lo_hi_lo_lo_lo_4};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_3 = {regroupV0_lo[2591:2588], regroupV0_lo[2575:2572]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_3 = {regroupV0_lo[2623:2620], regroupV0_lo[2607:2604]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_lo_lo_4 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_3, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_3 = {regroupV0_lo[2655:2652], regroupV0_lo[2639:2636]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_3 = {regroupV0_lo[2687:2684], regroupV0_lo[2671:2668]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_lo_hi_4 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_3, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_3};
  wire [31:0]        regroupV0_lo_hi_lo_hi_lo_lo_4 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_4, regroupV0_lo_hi_lo_hi_lo_lo_lo_4};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_3 = {regroupV0_lo[2719:2716], regroupV0_lo[2703:2700]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_3 = {regroupV0_lo[2751:2748], regroupV0_lo[2735:2732]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_hi_lo_4 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_3, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_3 = {regroupV0_lo[2783:2780], regroupV0_lo[2767:2764]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_3 = {regroupV0_lo[2815:2812], regroupV0_lo[2799:2796]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_hi_hi_4 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_3, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_3};
  wire [31:0]        regroupV0_lo_hi_lo_hi_lo_hi_4 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_4, regroupV0_lo_hi_lo_hi_lo_hi_lo_4};
  wire [63:0]        regroupV0_lo_hi_lo_hi_lo_4 = {regroupV0_lo_hi_lo_hi_lo_hi_4, regroupV0_lo_hi_lo_hi_lo_lo_4};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_3 = {regroupV0_lo[2847:2844], regroupV0_lo[2831:2828]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_3 = {regroupV0_lo[2879:2876], regroupV0_lo[2863:2860]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_lo_lo_4 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_3, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_3 = {regroupV0_lo[2911:2908], regroupV0_lo[2895:2892]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_3 = {regroupV0_lo[2943:2940], regroupV0_lo[2927:2924]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_lo_hi_4 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_3, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_3};
  wire [31:0]        regroupV0_lo_hi_lo_hi_hi_lo_4 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_4, regroupV0_lo_hi_lo_hi_hi_lo_lo_4};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_3 = {regroupV0_lo[2975:2972], regroupV0_lo[2959:2956]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_3 = {regroupV0_lo[3007:3004], regroupV0_lo[2991:2988]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_hi_lo_4 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_3, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_3 = {regroupV0_lo[3039:3036], regroupV0_lo[3023:3020]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_3 = {regroupV0_lo[3071:3068], regroupV0_lo[3055:3052]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_hi_hi_4 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_3, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_3};
  wire [31:0]        regroupV0_lo_hi_lo_hi_hi_hi_4 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_4, regroupV0_lo_hi_lo_hi_hi_hi_lo_4};
  wire [63:0]        regroupV0_lo_hi_lo_hi_hi_4 = {regroupV0_lo_hi_lo_hi_hi_hi_4, regroupV0_lo_hi_lo_hi_hi_lo_4};
  wire [127:0]       regroupV0_lo_hi_lo_hi_4 = {regroupV0_lo_hi_lo_hi_hi_4, regroupV0_lo_hi_lo_hi_lo_4};
  wire [255:0]       regroupV0_lo_hi_lo_4 = {regroupV0_lo_hi_lo_hi_4, regroupV0_lo_hi_lo_lo_4};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_3 = {regroupV0_lo[3103:3100], regroupV0_lo[3087:3084]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_3 = {regroupV0_lo[3135:3132], regroupV0_lo[3119:3116]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_lo_lo_4 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_3, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_3 = {regroupV0_lo[3167:3164], regroupV0_lo[3151:3148]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_3 = {regroupV0_lo[3199:3196], regroupV0_lo[3183:3180]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_lo_hi_4 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_3, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_3};
  wire [31:0]        regroupV0_lo_hi_hi_lo_lo_lo_4 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_4, regroupV0_lo_hi_hi_lo_lo_lo_lo_4};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_3 = {regroupV0_lo[3231:3228], regroupV0_lo[3215:3212]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_3 = {regroupV0_lo[3263:3260], regroupV0_lo[3247:3244]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_hi_lo_4 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_3, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_3 = {regroupV0_lo[3295:3292], regroupV0_lo[3279:3276]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_3 = {regroupV0_lo[3327:3324], regroupV0_lo[3311:3308]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_hi_hi_4 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_3, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_3};
  wire [31:0]        regroupV0_lo_hi_hi_lo_lo_hi_4 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_4, regroupV0_lo_hi_hi_lo_lo_hi_lo_4};
  wire [63:0]        regroupV0_lo_hi_hi_lo_lo_4 = {regroupV0_lo_hi_hi_lo_lo_hi_4, regroupV0_lo_hi_hi_lo_lo_lo_4};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_3 = {regroupV0_lo[3359:3356], regroupV0_lo[3343:3340]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_3 = {regroupV0_lo[3391:3388], regroupV0_lo[3375:3372]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_lo_lo_4 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_3, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_3 = {regroupV0_lo[3423:3420], regroupV0_lo[3407:3404]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_3 = {regroupV0_lo[3455:3452], regroupV0_lo[3439:3436]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_lo_hi_4 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_3, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_3};
  wire [31:0]        regroupV0_lo_hi_hi_lo_hi_lo_4 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_4, regroupV0_lo_hi_hi_lo_hi_lo_lo_4};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_3 = {regroupV0_lo[3487:3484], regroupV0_lo[3471:3468]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_3 = {regroupV0_lo[3519:3516], regroupV0_lo[3503:3500]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_hi_lo_4 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_3, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_3 = {regroupV0_lo[3551:3548], regroupV0_lo[3535:3532]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_3 = {regroupV0_lo[3583:3580], regroupV0_lo[3567:3564]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_hi_hi_4 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_3, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_3};
  wire [31:0]        regroupV0_lo_hi_hi_lo_hi_hi_4 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_4, regroupV0_lo_hi_hi_lo_hi_hi_lo_4};
  wire [63:0]        regroupV0_lo_hi_hi_lo_hi_4 = {regroupV0_lo_hi_hi_lo_hi_hi_4, regroupV0_lo_hi_hi_lo_hi_lo_4};
  wire [127:0]       regroupV0_lo_hi_hi_lo_4 = {regroupV0_lo_hi_hi_lo_hi_4, regroupV0_lo_hi_hi_lo_lo_4};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_3 = {regroupV0_lo[3615:3612], regroupV0_lo[3599:3596]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_3 = {regroupV0_lo[3647:3644], regroupV0_lo[3631:3628]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_lo_lo_4 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_3, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_3 = {regroupV0_lo[3679:3676], regroupV0_lo[3663:3660]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_3 = {regroupV0_lo[3711:3708], regroupV0_lo[3695:3692]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_lo_hi_4 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_3, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_3};
  wire [31:0]        regroupV0_lo_hi_hi_hi_lo_lo_4 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_4, regroupV0_lo_hi_hi_hi_lo_lo_lo_4};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_3 = {regroupV0_lo[3743:3740], regroupV0_lo[3727:3724]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_3 = {regroupV0_lo[3775:3772], regroupV0_lo[3759:3756]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_hi_lo_4 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_3, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_3 = {regroupV0_lo[3807:3804], regroupV0_lo[3791:3788]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_3 = {regroupV0_lo[3839:3836], regroupV0_lo[3823:3820]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_hi_hi_4 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_3, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_3};
  wire [31:0]        regroupV0_lo_hi_hi_hi_lo_hi_4 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_4, regroupV0_lo_hi_hi_hi_lo_hi_lo_4};
  wire [63:0]        regroupV0_lo_hi_hi_hi_lo_4 = {regroupV0_lo_hi_hi_hi_lo_hi_4, regroupV0_lo_hi_hi_hi_lo_lo_4};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_3 = {regroupV0_lo[3871:3868], regroupV0_lo[3855:3852]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_3 = {regroupV0_lo[3903:3900], regroupV0_lo[3887:3884]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_lo_lo_4 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_3, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_3 = {regroupV0_lo[3935:3932], regroupV0_lo[3919:3916]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_3 = {regroupV0_lo[3967:3964], regroupV0_lo[3951:3948]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_lo_hi_4 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_3, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_3};
  wire [31:0]        regroupV0_lo_hi_hi_hi_hi_lo_4 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_4, regroupV0_lo_hi_hi_hi_hi_lo_lo_4};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_3 = {regroupV0_lo[3999:3996], regroupV0_lo[3983:3980]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_3 = {regroupV0_lo[4031:4028], regroupV0_lo[4015:4012]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_hi_lo_4 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_3, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_3 = {regroupV0_lo[4063:4060], regroupV0_lo[4047:4044]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_3 = {regroupV0_lo[4095:4092], regroupV0_lo[4079:4076]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_hi_hi_4 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_3, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_3};
  wire [31:0]        regroupV0_lo_hi_hi_hi_hi_hi_4 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_4, regroupV0_lo_hi_hi_hi_hi_hi_lo_4};
  wire [63:0]        regroupV0_lo_hi_hi_hi_hi_4 = {regroupV0_lo_hi_hi_hi_hi_hi_4, regroupV0_lo_hi_hi_hi_hi_lo_4};
  wire [127:0]       regroupV0_lo_hi_hi_hi_4 = {regroupV0_lo_hi_hi_hi_hi_4, regroupV0_lo_hi_hi_hi_lo_4};
  wire [255:0]       regroupV0_lo_hi_hi_4 = {regroupV0_lo_hi_hi_hi_4, regroupV0_lo_hi_hi_lo_4};
  wire [511:0]       regroupV0_lo_hi_4 = {regroupV0_lo_hi_hi_4, regroupV0_lo_hi_lo_4};
  wire [1023:0]      regroupV0_lo_4 = {regroupV0_lo_hi_4, regroupV0_lo_lo_4};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_3 = {regroupV0_hi[31:28], regroupV0_hi[15:12]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_3 = {regroupV0_hi[63:60], regroupV0_hi[47:44]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_lo_lo_4 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_3 = {regroupV0_hi[95:92], regroupV0_hi[79:76]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_3 = {regroupV0_hi[127:124], regroupV0_hi[111:108]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_lo_hi_4 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_3, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_3};
  wire [31:0]        regroupV0_hi_lo_lo_lo_lo_lo_4 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_4, regroupV0_hi_lo_lo_lo_lo_lo_lo_4};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_3 = {regroupV0_hi[159:156], regroupV0_hi[143:140]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_3 = {regroupV0_hi[191:188], regroupV0_hi[175:172]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_hi_lo_4 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_3, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_3 = {regroupV0_hi[223:220], regroupV0_hi[207:204]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_3 = {regroupV0_hi[255:252], regroupV0_hi[239:236]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_hi_hi_4 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_3, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_3};
  wire [31:0]        regroupV0_hi_lo_lo_lo_lo_hi_4 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_4, regroupV0_hi_lo_lo_lo_lo_hi_lo_4};
  wire [63:0]        regroupV0_hi_lo_lo_lo_lo_4 = {regroupV0_hi_lo_lo_lo_lo_hi_4, regroupV0_hi_lo_lo_lo_lo_lo_4};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_3 = {regroupV0_hi[287:284], regroupV0_hi[271:268]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_3 = {regroupV0_hi[319:316], regroupV0_hi[303:300]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_lo_lo_4 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_3 = {regroupV0_hi[351:348], regroupV0_hi[335:332]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_3 = {regroupV0_hi[383:380], regroupV0_hi[367:364]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_lo_hi_4 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_3, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_3};
  wire [31:0]        regroupV0_hi_lo_lo_lo_hi_lo_4 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_4, regroupV0_hi_lo_lo_lo_hi_lo_lo_4};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_3 = {regroupV0_hi[415:412], regroupV0_hi[399:396]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_3 = {regroupV0_hi[447:444], regroupV0_hi[431:428]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_hi_lo_4 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_3, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_3 = {regroupV0_hi[479:476], regroupV0_hi[463:460]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_3 = {regroupV0_hi[511:508], regroupV0_hi[495:492]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_hi_hi_4 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_3, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_3};
  wire [31:0]        regroupV0_hi_lo_lo_lo_hi_hi_4 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_4, regroupV0_hi_lo_lo_lo_hi_hi_lo_4};
  wire [63:0]        regroupV0_hi_lo_lo_lo_hi_4 = {regroupV0_hi_lo_lo_lo_hi_hi_4, regroupV0_hi_lo_lo_lo_hi_lo_4};
  wire [127:0]       regroupV0_hi_lo_lo_lo_4 = {regroupV0_hi_lo_lo_lo_hi_4, regroupV0_hi_lo_lo_lo_lo_4};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_3 = {regroupV0_hi[543:540], regroupV0_hi[527:524]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_3 = {regroupV0_hi[575:572], regroupV0_hi[559:556]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_lo_lo_4 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_3, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_3 = {regroupV0_hi[607:604], regroupV0_hi[591:588]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_3 = {regroupV0_hi[639:636], regroupV0_hi[623:620]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_lo_hi_4 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_3, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_3};
  wire [31:0]        regroupV0_hi_lo_lo_hi_lo_lo_4 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_4, regroupV0_hi_lo_lo_hi_lo_lo_lo_4};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_3 = {regroupV0_hi[671:668], regroupV0_hi[655:652]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_3 = {regroupV0_hi[703:700], regroupV0_hi[687:684]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_hi_lo_4 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_3, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_3 = {regroupV0_hi[735:732], regroupV0_hi[719:716]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_3 = {regroupV0_hi[767:764], regroupV0_hi[751:748]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_hi_hi_4 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_3, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_3};
  wire [31:0]        regroupV0_hi_lo_lo_hi_lo_hi_4 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_4, regroupV0_hi_lo_lo_hi_lo_hi_lo_4};
  wire [63:0]        regroupV0_hi_lo_lo_hi_lo_4 = {regroupV0_hi_lo_lo_hi_lo_hi_4, regroupV0_hi_lo_lo_hi_lo_lo_4};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_3 = {regroupV0_hi[799:796], regroupV0_hi[783:780]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_3 = {regroupV0_hi[831:828], regroupV0_hi[815:812]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_lo_lo_4 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_3, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_3 = {regroupV0_hi[863:860], regroupV0_hi[847:844]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_3 = {regroupV0_hi[895:892], regroupV0_hi[879:876]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_lo_hi_4 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_3, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_3};
  wire [31:0]        regroupV0_hi_lo_lo_hi_hi_lo_4 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_4, regroupV0_hi_lo_lo_hi_hi_lo_lo_4};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_3 = {regroupV0_hi[927:924], regroupV0_hi[911:908]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_3 = {regroupV0_hi[959:956], regroupV0_hi[943:940]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_hi_lo_4 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_3, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_3 = {regroupV0_hi[991:988], regroupV0_hi[975:972]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_3 = {regroupV0_hi[1023:1020], regroupV0_hi[1007:1004]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_hi_hi_4 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_3, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_3};
  wire [31:0]        regroupV0_hi_lo_lo_hi_hi_hi_4 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_4, regroupV0_hi_lo_lo_hi_hi_hi_lo_4};
  wire [63:0]        regroupV0_hi_lo_lo_hi_hi_4 = {regroupV0_hi_lo_lo_hi_hi_hi_4, regroupV0_hi_lo_lo_hi_hi_lo_4};
  wire [127:0]       regroupV0_hi_lo_lo_hi_4 = {regroupV0_hi_lo_lo_hi_hi_4, regroupV0_hi_lo_lo_hi_lo_4};
  wire [255:0]       regroupV0_hi_lo_lo_4 = {regroupV0_hi_lo_lo_hi_4, regroupV0_hi_lo_lo_lo_4};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_3 = {regroupV0_hi[1055:1052], regroupV0_hi[1039:1036]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_3 = {regroupV0_hi[1087:1084], regroupV0_hi[1071:1068]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_lo_lo_4 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_3, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_3 = {regroupV0_hi[1119:1116], regroupV0_hi[1103:1100]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_3 = {regroupV0_hi[1151:1148], regroupV0_hi[1135:1132]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_lo_hi_4 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_3, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_3};
  wire [31:0]        regroupV0_hi_lo_hi_lo_lo_lo_4 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_4, regroupV0_hi_lo_hi_lo_lo_lo_lo_4};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_3 = {regroupV0_hi[1183:1180], regroupV0_hi[1167:1164]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_3 = {regroupV0_hi[1215:1212], regroupV0_hi[1199:1196]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_hi_lo_4 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_3, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_3 = {regroupV0_hi[1247:1244], regroupV0_hi[1231:1228]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_3 = {regroupV0_hi[1279:1276], regroupV0_hi[1263:1260]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_hi_hi_4 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_3, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_3};
  wire [31:0]        regroupV0_hi_lo_hi_lo_lo_hi_4 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_4, regroupV0_hi_lo_hi_lo_lo_hi_lo_4};
  wire [63:0]        regroupV0_hi_lo_hi_lo_lo_4 = {regroupV0_hi_lo_hi_lo_lo_hi_4, regroupV0_hi_lo_hi_lo_lo_lo_4};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_3 = {regroupV0_hi[1311:1308], regroupV0_hi[1295:1292]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_3 = {regroupV0_hi[1343:1340], regroupV0_hi[1327:1324]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_lo_lo_4 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_3, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_3 = {regroupV0_hi[1375:1372], regroupV0_hi[1359:1356]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_3 = {regroupV0_hi[1407:1404], regroupV0_hi[1391:1388]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_lo_hi_4 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_3, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_3};
  wire [31:0]        regroupV0_hi_lo_hi_lo_hi_lo_4 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_4, regroupV0_hi_lo_hi_lo_hi_lo_lo_4};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_3 = {regroupV0_hi[1439:1436], regroupV0_hi[1423:1420]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_3 = {regroupV0_hi[1471:1468], regroupV0_hi[1455:1452]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_hi_lo_4 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_3, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_3 = {regroupV0_hi[1503:1500], regroupV0_hi[1487:1484]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_3 = {regroupV0_hi[1535:1532], regroupV0_hi[1519:1516]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_hi_hi_4 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_3, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_3};
  wire [31:0]        regroupV0_hi_lo_hi_lo_hi_hi_4 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_4, regroupV0_hi_lo_hi_lo_hi_hi_lo_4};
  wire [63:0]        regroupV0_hi_lo_hi_lo_hi_4 = {regroupV0_hi_lo_hi_lo_hi_hi_4, regroupV0_hi_lo_hi_lo_hi_lo_4};
  wire [127:0]       regroupV0_hi_lo_hi_lo_4 = {regroupV0_hi_lo_hi_lo_hi_4, regroupV0_hi_lo_hi_lo_lo_4};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_3 = {regroupV0_hi[1567:1564], regroupV0_hi[1551:1548]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_3 = {regroupV0_hi[1599:1596], regroupV0_hi[1583:1580]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_lo_lo_4 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_3, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_3 = {regroupV0_hi[1631:1628], regroupV0_hi[1615:1612]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_3 = {regroupV0_hi[1663:1660], regroupV0_hi[1647:1644]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_lo_hi_4 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_3, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_3};
  wire [31:0]        regroupV0_hi_lo_hi_hi_lo_lo_4 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_4, regroupV0_hi_lo_hi_hi_lo_lo_lo_4};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_3 = {regroupV0_hi[1695:1692], regroupV0_hi[1679:1676]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_3 = {regroupV0_hi[1727:1724], regroupV0_hi[1711:1708]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_hi_lo_4 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_3, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_3 = {regroupV0_hi[1759:1756], regroupV0_hi[1743:1740]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_3 = {regroupV0_hi[1791:1788], regroupV0_hi[1775:1772]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_hi_hi_4 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_3, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_3};
  wire [31:0]        regroupV0_hi_lo_hi_hi_lo_hi_4 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_4, regroupV0_hi_lo_hi_hi_lo_hi_lo_4};
  wire [63:0]        regroupV0_hi_lo_hi_hi_lo_4 = {regroupV0_hi_lo_hi_hi_lo_hi_4, regroupV0_hi_lo_hi_hi_lo_lo_4};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_3 = {regroupV0_hi[1823:1820], regroupV0_hi[1807:1804]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_3 = {regroupV0_hi[1855:1852], regroupV0_hi[1839:1836]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_lo_lo_4 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_3, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_3 = {regroupV0_hi[1887:1884], regroupV0_hi[1871:1868]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_3 = {regroupV0_hi[1919:1916], regroupV0_hi[1903:1900]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_lo_hi_4 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_3, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_3};
  wire [31:0]        regroupV0_hi_lo_hi_hi_hi_lo_4 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_4, regroupV0_hi_lo_hi_hi_hi_lo_lo_4};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_3 = {regroupV0_hi[1951:1948], regroupV0_hi[1935:1932]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_3 = {regroupV0_hi[1983:1980], regroupV0_hi[1967:1964]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_hi_lo_4 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_3, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_3 = {regroupV0_hi[2015:2012], regroupV0_hi[1999:1996]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_3 = {regroupV0_hi[2047:2044], regroupV0_hi[2031:2028]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_hi_hi_4 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_3, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_3};
  wire [31:0]        regroupV0_hi_lo_hi_hi_hi_hi_4 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_4, regroupV0_hi_lo_hi_hi_hi_hi_lo_4};
  wire [63:0]        regroupV0_hi_lo_hi_hi_hi_4 = {regroupV0_hi_lo_hi_hi_hi_hi_4, regroupV0_hi_lo_hi_hi_hi_lo_4};
  wire [127:0]       regroupV0_hi_lo_hi_hi_4 = {regroupV0_hi_lo_hi_hi_hi_4, regroupV0_hi_lo_hi_hi_lo_4};
  wire [255:0]       regroupV0_hi_lo_hi_4 = {regroupV0_hi_lo_hi_hi_4, regroupV0_hi_lo_hi_lo_4};
  wire [511:0]       regroupV0_hi_lo_4 = {regroupV0_hi_lo_hi_4, regroupV0_hi_lo_lo_4};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_3 = {regroupV0_hi[2079:2076], regroupV0_hi[2063:2060]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_3 = {regroupV0_hi[2111:2108], regroupV0_hi[2095:2092]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_lo_lo_4 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_3, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_3 = {regroupV0_hi[2143:2140], regroupV0_hi[2127:2124]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_3 = {regroupV0_hi[2175:2172], regroupV0_hi[2159:2156]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_lo_hi_4 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_3, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_3};
  wire [31:0]        regroupV0_hi_hi_lo_lo_lo_lo_4 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_4, regroupV0_hi_hi_lo_lo_lo_lo_lo_4};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_3 = {regroupV0_hi[2207:2204], regroupV0_hi[2191:2188]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_3 = {regroupV0_hi[2239:2236], regroupV0_hi[2223:2220]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_hi_lo_4 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_3, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_3 = {regroupV0_hi[2271:2268], regroupV0_hi[2255:2252]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_3 = {regroupV0_hi[2303:2300], regroupV0_hi[2287:2284]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_hi_hi_4 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_3, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_3};
  wire [31:0]        regroupV0_hi_hi_lo_lo_lo_hi_4 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_4, regroupV0_hi_hi_lo_lo_lo_hi_lo_4};
  wire [63:0]        regroupV0_hi_hi_lo_lo_lo_4 = {regroupV0_hi_hi_lo_lo_lo_hi_4, regroupV0_hi_hi_lo_lo_lo_lo_4};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_3 = {regroupV0_hi[2335:2332], regroupV0_hi[2319:2316]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_3 = {regroupV0_hi[2367:2364], regroupV0_hi[2351:2348]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_lo_lo_4 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_3, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_3 = {regroupV0_hi[2399:2396], regroupV0_hi[2383:2380]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_3 = {regroupV0_hi[2431:2428], regroupV0_hi[2415:2412]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_lo_hi_4 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_3, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_3};
  wire [31:0]        regroupV0_hi_hi_lo_lo_hi_lo_4 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_4, regroupV0_hi_hi_lo_lo_hi_lo_lo_4};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_3 = {regroupV0_hi[2463:2460], regroupV0_hi[2447:2444]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_3 = {regroupV0_hi[2495:2492], regroupV0_hi[2479:2476]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_hi_lo_4 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_3, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_3 = {regroupV0_hi[2527:2524], regroupV0_hi[2511:2508]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_3 = {regroupV0_hi[2559:2556], regroupV0_hi[2543:2540]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_hi_hi_4 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_3, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_3};
  wire [31:0]        regroupV0_hi_hi_lo_lo_hi_hi_4 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_4, regroupV0_hi_hi_lo_lo_hi_hi_lo_4};
  wire [63:0]        regroupV0_hi_hi_lo_lo_hi_4 = {regroupV0_hi_hi_lo_lo_hi_hi_4, regroupV0_hi_hi_lo_lo_hi_lo_4};
  wire [127:0]       regroupV0_hi_hi_lo_lo_4 = {regroupV0_hi_hi_lo_lo_hi_4, regroupV0_hi_hi_lo_lo_lo_4};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_3 = {regroupV0_hi[2591:2588], regroupV0_hi[2575:2572]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_3 = {regroupV0_hi[2623:2620], regroupV0_hi[2607:2604]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_lo_lo_4 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_3, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_3 = {regroupV0_hi[2655:2652], regroupV0_hi[2639:2636]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_3 = {regroupV0_hi[2687:2684], regroupV0_hi[2671:2668]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_lo_hi_4 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_3, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_3};
  wire [31:0]        regroupV0_hi_hi_lo_hi_lo_lo_4 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_4, regroupV0_hi_hi_lo_hi_lo_lo_lo_4};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_3 = {regroupV0_hi[2719:2716], regroupV0_hi[2703:2700]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_3 = {regroupV0_hi[2751:2748], regroupV0_hi[2735:2732]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_hi_lo_4 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_3, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_3 = {regroupV0_hi[2783:2780], regroupV0_hi[2767:2764]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_3 = {regroupV0_hi[2815:2812], regroupV0_hi[2799:2796]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_hi_hi_4 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_3, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_3};
  wire [31:0]        regroupV0_hi_hi_lo_hi_lo_hi_4 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_4, regroupV0_hi_hi_lo_hi_lo_hi_lo_4};
  wire [63:0]        regroupV0_hi_hi_lo_hi_lo_4 = {regroupV0_hi_hi_lo_hi_lo_hi_4, regroupV0_hi_hi_lo_hi_lo_lo_4};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_3 = {regroupV0_hi[2847:2844], regroupV0_hi[2831:2828]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_3 = {regroupV0_hi[2879:2876], regroupV0_hi[2863:2860]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_lo_lo_4 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_3, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_3 = {regroupV0_hi[2911:2908], regroupV0_hi[2895:2892]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_3 = {regroupV0_hi[2943:2940], regroupV0_hi[2927:2924]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_lo_hi_4 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_3, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_3};
  wire [31:0]        regroupV0_hi_hi_lo_hi_hi_lo_4 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_4, regroupV0_hi_hi_lo_hi_hi_lo_lo_4};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_3 = {regroupV0_hi[2975:2972], regroupV0_hi[2959:2956]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_3 = {regroupV0_hi[3007:3004], regroupV0_hi[2991:2988]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_hi_lo_4 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_3, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_3 = {regroupV0_hi[3039:3036], regroupV0_hi[3023:3020]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_3 = {regroupV0_hi[3071:3068], regroupV0_hi[3055:3052]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_hi_hi_4 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_3, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_3};
  wire [31:0]        regroupV0_hi_hi_lo_hi_hi_hi_4 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_4, regroupV0_hi_hi_lo_hi_hi_hi_lo_4};
  wire [63:0]        regroupV0_hi_hi_lo_hi_hi_4 = {regroupV0_hi_hi_lo_hi_hi_hi_4, regroupV0_hi_hi_lo_hi_hi_lo_4};
  wire [127:0]       regroupV0_hi_hi_lo_hi_4 = {regroupV0_hi_hi_lo_hi_hi_4, regroupV0_hi_hi_lo_hi_lo_4};
  wire [255:0]       regroupV0_hi_hi_lo_4 = {regroupV0_hi_hi_lo_hi_4, regroupV0_hi_hi_lo_lo_4};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_3 = {regroupV0_hi[3103:3100], regroupV0_hi[3087:3084]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_3 = {regroupV0_hi[3135:3132], regroupV0_hi[3119:3116]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_lo_lo_4 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_3, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_3 = {regroupV0_hi[3167:3164], regroupV0_hi[3151:3148]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_3 = {regroupV0_hi[3199:3196], regroupV0_hi[3183:3180]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_lo_hi_4 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_3, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_3};
  wire [31:0]        regroupV0_hi_hi_hi_lo_lo_lo_4 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_4, regroupV0_hi_hi_hi_lo_lo_lo_lo_4};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_3 = {regroupV0_hi[3231:3228], regroupV0_hi[3215:3212]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_3 = {regroupV0_hi[3263:3260], regroupV0_hi[3247:3244]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_hi_lo_4 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_3, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_3 = {regroupV0_hi[3295:3292], regroupV0_hi[3279:3276]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_3 = {regroupV0_hi[3327:3324], regroupV0_hi[3311:3308]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_hi_hi_4 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_3, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_3};
  wire [31:0]        regroupV0_hi_hi_hi_lo_lo_hi_4 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_4, regroupV0_hi_hi_hi_lo_lo_hi_lo_4};
  wire [63:0]        regroupV0_hi_hi_hi_lo_lo_4 = {regroupV0_hi_hi_hi_lo_lo_hi_4, regroupV0_hi_hi_hi_lo_lo_lo_4};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_3 = {regroupV0_hi[3359:3356], regroupV0_hi[3343:3340]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_3 = {regroupV0_hi[3391:3388], regroupV0_hi[3375:3372]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_lo_lo_4 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_3, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_3 = {regroupV0_hi[3423:3420], regroupV0_hi[3407:3404]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_3 = {regroupV0_hi[3455:3452], regroupV0_hi[3439:3436]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_lo_hi_4 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_3, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_3};
  wire [31:0]        regroupV0_hi_hi_hi_lo_hi_lo_4 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_4, regroupV0_hi_hi_hi_lo_hi_lo_lo_4};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_3 = {regroupV0_hi[3487:3484], regroupV0_hi[3471:3468]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_3 = {regroupV0_hi[3519:3516], regroupV0_hi[3503:3500]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_hi_lo_4 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_3, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_3 = {regroupV0_hi[3551:3548], regroupV0_hi[3535:3532]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_3 = {regroupV0_hi[3583:3580], regroupV0_hi[3567:3564]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_hi_hi_4 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_3};
  wire [31:0]        regroupV0_hi_hi_hi_lo_hi_hi_4 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_4, regroupV0_hi_hi_hi_lo_hi_hi_lo_4};
  wire [63:0]        regroupV0_hi_hi_hi_lo_hi_4 = {regroupV0_hi_hi_hi_lo_hi_hi_4, regroupV0_hi_hi_hi_lo_hi_lo_4};
  wire [127:0]       regroupV0_hi_hi_hi_lo_4 = {regroupV0_hi_hi_hi_lo_hi_4, regroupV0_hi_hi_hi_lo_lo_4};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_3 = {regroupV0_hi[3615:3612], regroupV0_hi[3599:3596]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_3 = {regroupV0_hi[3647:3644], regroupV0_hi[3631:3628]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_lo_lo_4 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_3, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_3 = {regroupV0_hi[3679:3676], regroupV0_hi[3663:3660]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_3 = {regroupV0_hi[3711:3708], regroupV0_hi[3695:3692]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_lo_hi_4 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_3, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_3};
  wire [31:0]        regroupV0_hi_hi_hi_hi_lo_lo_4 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_4, regroupV0_hi_hi_hi_hi_lo_lo_lo_4};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_3 = {regroupV0_hi[3743:3740], regroupV0_hi[3727:3724]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_3 = {regroupV0_hi[3775:3772], regroupV0_hi[3759:3756]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_hi_lo_4 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_3, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_3 = {regroupV0_hi[3807:3804], regroupV0_hi[3791:3788]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_3 = {regroupV0_hi[3839:3836], regroupV0_hi[3823:3820]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_hi_hi_4 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_3, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_3};
  wire [31:0]        regroupV0_hi_hi_hi_hi_lo_hi_4 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_4, regroupV0_hi_hi_hi_hi_lo_hi_lo_4};
  wire [63:0]        regroupV0_hi_hi_hi_hi_lo_4 = {regroupV0_hi_hi_hi_hi_lo_hi_4, regroupV0_hi_hi_hi_hi_lo_lo_4};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_3 = {regroupV0_hi[3871:3868], regroupV0_hi[3855:3852]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_3 = {regroupV0_hi[3903:3900], regroupV0_hi[3887:3884]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_lo_lo_4 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_3, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_3 = {regroupV0_hi[3935:3932], regroupV0_hi[3919:3916]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_3 = {regroupV0_hi[3967:3964], regroupV0_hi[3951:3948]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_lo_hi_4 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_3, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_3};
  wire [31:0]        regroupV0_hi_hi_hi_hi_hi_lo_4 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_4, regroupV0_hi_hi_hi_hi_hi_lo_lo_4};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_3 = {regroupV0_hi[3999:3996], regroupV0_hi[3983:3980]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_3 = {regroupV0_hi[4031:4028], regroupV0_hi[4015:4012]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_hi_lo_4 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_3, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_3 = {regroupV0_hi[4063:4060], regroupV0_hi[4047:4044]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_3 = {regroupV0_hi[4095:4092], regroupV0_hi[4079:4076]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_hi_hi_4 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_3};
  wire [31:0]        regroupV0_hi_hi_hi_hi_hi_hi_4 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_4, regroupV0_hi_hi_hi_hi_hi_hi_lo_4};
  wire [63:0]        regroupV0_hi_hi_hi_hi_hi_4 = {regroupV0_hi_hi_hi_hi_hi_hi_4, regroupV0_hi_hi_hi_hi_hi_lo_4};
  wire [127:0]       regroupV0_hi_hi_hi_hi_4 = {regroupV0_hi_hi_hi_hi_hi_4, regroupV0_hi_hi_hi_hi_lo_4};
  wire [255:0]       regroupV0_hi_hi_hi_4 = {regroupV0_hi_hi_hi_hi_4, regroupV0_hi_hi_hi_lo_4};
  wire [511:0]       regroupV0_hi_hi_4 = {regroupV0_hi_hi_hi_4, regroupV0_hi_hi_lo_4};
  wire [1023:0]      regroupV0_hi_4 = {regroupV0_hi_hi_4, regroupV0_hi_lo_4};
  wire [4095:0]      regroupV0_lo_5 = {regroupV0_hi_2, regroupV0_lo_2, regroupV0_hi_1, regroupV0_lo_1};
  wire [4095:0]      regroupV0_hi_5 = {regroupV0_hi_4, regroupV0_lo_4, regroupV0_hi_3, regroupV0_lo_3};
  wire [8191:0]      regroupV0_0 = {regroupV0_hi_5, regroupV0_lo_5};
  wire [127:0]       regroupV0_lo_lo_lo_lo_lo_lo_5 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_5, regroupV0_lo_lo_lo_lo_lo_lo_lo_5};
  wire [127:0]       regroupV0_lo_lo_lo_lo_lo_hi_5 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_5, regroupV0_lo_lo_lo_lo_lo_hi_lo_5};
  wire [255:0]       regroupV0_lo_lo_lo_lo_lo_5 = {regroupV0_lo_lo_lo_lo_lo_hi_5, regroupV0_lo_lo_lo_lo_lo_lo_5};
  wire [127:0]       regroupV0_lo_lo_lo_lo_hi_lo_5 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_5, regroupV0_lo_lo_lo_lo_hi_lo_lo_5};
  wire [127:0]       regroupV0_lo_lo_lo_lo_hi_hi_5 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_5, regroupV0_lo_lo_lo_lo_hi_hi_lo_5};
  wire [255:0]       regroupV0_lo_lo_lo_lo_hi_5 = {regroupV0_lo_lo_lo_lo_hi_hi_5, regroupV0_lo_lo_lo_lo_hi_lo_5};
  wire [511:0]       regroupV0_lo_lo_lo_lo_5 = {regroupV0_lo_lo_lo_lo_hi_5, regroupV0_lo_lo_lo_lo_lo_5};
  wire [127:0]       regroupV0_lo_lo_lo_hi_lo_lo_5 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_5, regroupV0_lo_lo_lo_hi_lo_lo_lo_5};
  wire [127:0]       regroupV0_lo_lo_lo_hi_lo_hi_5 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_5, regroupV0_lo_lo_lo_hi_lo_hi_lo_5};
  wire [255:0]       regroupV0_lo_lo_lo_hi_lo_5 = {regroupV0_lo_lo_lo_hi_lo_hi_5, regroupV0_lo_lo_lo_hi_lo_lo_5};
  wire [127:0]       regroupV0_lo_lo_lo_hi_hi_lo_5 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_5, regroupV0_lo_lo_lo_hi_hi_lo_lo_5};
  wire [127:0]       regroupV0_lo_lo_lo_hi_hi_hi_5 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_5, regroupV0_lo_lo_lo_hi_hi_hi_lo_5};
  wire [255:0]       regroupV0_lo_lo_lo_hi_hi_5 = {regroupV0_lo_lo_lo_hi_hi_hi_5, regroupV0_lo_lo_lo_hi_hi_lo_5};
  wire [511:0]       regroupV0_lo_lo_lo_hi_5 = {regroupV0_lo_lo_lo_hi_hi_5, regroupV0_lo_lo_lo_hi_lo_5};
  wire [1023:0]      regroupV0_lo_lo_lo_5 = {regroupV0_lo_lo_lo_hi_5, regroupV0_lo_lo_lo_lo_5};
  wire [127:0]       regroupV0_lo_lo_hi_lo_lo_lo_5 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_5, regroupV0_lo_lo_hi_lo_lo_lo_lo_5};
  wire [127:0]       regroupV0_lo_lo_hi_lo_lo_hi_5 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_5, regroupV0_lo_lo_hi_lo_lo_hi_lo_5};
  wire [255:0]       regroupV0_lo_lo_hi_lo_lo_5 = {regroupV0_lo_lo_hi_lo_lo_hi_5, regroupV0_lo_lo_hi_lo_lo_lo_5};
  wire [127:0]       regroupV0_lo_lo_hi_lo_hi_lo_5 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_5, regroupV0_lo_lo_hi_lo_hi_lo_lo_5};
  wire [127:0]       regroupV0_lo_lo_hi_lo_hi_hi_5 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_5, regroupV0_lo_lo_hi_lo_hi_hi_lo_5};
  wire [255:0]       regroupV0_lo_lo_hi_lo_hi_5 = {regroupV0_lo_lo_hi_lo_hi_hi_5, regroupV0_lo_lo_hi_lo_hi_lo_5};
  wire [511:0]       regroupV0_lo_lo_hi_lo_5 = {regroupV0_lo_lo_hi_lo_hi_5, regroupV0_lo_lo_hi_lo_lo_5};
  wire [127:0]       regroupV0_lo_lo_hi_hi_lo_lo_5 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_5, regroupV0_lo_lo_hi_hi_lo_lo_lo_5};
  wire [127:0]       regroupV0_lo_lo_hi_hi_lo_hi_5 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_5, regroupV0_lo_lo_hi_hi_lo_hi_lo_5};
  wire [255:0]       regroupV0_lo_lo_hi_hi_lo_5 = {regroupV0_lo_lo_hi_hi_lo_hi_5, regroupV0_lo_lo_hi_hi_lo_lo_5};
  wire [127:0]       regroupV0_lo_lo_hi_hi_hi_lo_5 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_5, regroupV0_lo_lo_hi_hi_hi_lo_lo_5};
  wire [127:0]       regroupV0_lo_lo_hi_hi_hi_hi_5 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_5, regroupV0_lo_lo_hi_hi_hi_hi_lo_5};
  wire [255:0]       regroupV0_lo_lo_hi_hi_hi_5 = {regroupV0_lo_lo_hi_hi_hi_hi_5, regroupV0_lo_lo_hi_hi_hi_lo_5};
  wire [511:0]       regroupV0_lo_lo_hi_hi_5 = {regroupV0_lo_lo_hi_hi_hi_5, regroupV0_lo_lo_hi_hi_lo_5};
  wire [1023:0]      regroupV0_lo_lo_hi_5 = {regroupV0_lo_lo_hi_hi_5, regroupV0_lo_lo_hi_lo_5};
  wire [2047:0]      regroupV0_lo_lo_5 = {regroupV0_lo_lo_hi_5, regroupV0_lo_lo_lo_5};
  wire [127:0]       regroupV0_lo_hi_lo_lo_lo_lo_5 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_5, regroupV0_lo_hi_lo_lo_lo_lo_lo_5};
  wire [127:0]       regroupV0_lo_hi_lo_lo_lo_hi_5 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_5, regroupV0_lo_hi_lo_lo_lo_hi_lo_5};
  wire [255:0]       regroupV0_lo_hi_lo_lo_lo_5 = {regroupV0_lo_hi_lo_lo_lo_hi_5, regroupV0_lo_hi_lo_lo_lo_lo_5};
  wire [127:0]       regroupV0_lo_hi_lo_lo_hi_lo_5 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_5, regroupV0_lo_hi_lo_lo_hi_lo_lo_5};
  wire [127:0]       regroupV0_lo_hi_lo_lo_hi_hi_5 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_5, regroupV0_lo_hi_lo_lo_hi_hi_lo_5};
  wire [255:0]       regroupV0_lo_hi_lo_lo_hi_5 = {regroupV0_lo_hi_lo_lo_hi_hi_5, regroupV0_lo_hi_lo_lo_hi_lo_5};
  wire [511:0]       regroupV0_lo_hi_lo_lo_5 = {regroupV0_lo_hi_lo_lo_hi_5, regroupV0_lo_hi_lo_lo_lo_5};
  wire [127:0]       regroupV0_lo_hi_lo_hi_lo_lo_5 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_5, regroupV0_lo_hi_lo_hi_lo_lo_lo_5};
  wire [127:0]       regroupV0_lo_hi_lo_hi_lo_hi_5 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_5, regroupV0_lo_hi_lo_hi_lo_hi_lo_5};
  wire [255:0]       regroupV0_lo_hi_lo_hi_lo_5 = {regroupV0_lo_hi_lo_hi_lo_hi_5, regroupV0_lo_hi_lo_hi_lo_lo_5};
  wire [127:0]       regroupV0_lo_hi_lo_hi_hi_lo_5 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_5, regroupV0_lo_hi_lo_hi_hi_lo_lo_5};
  wire [127:0]       regroupV0_lo_hi_lo_hi_hi_hi_5 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_5, regroupV0_lo_hi_lo_hi_hi_hi_lo_5};
  wire [255:0]       regroupV0_lo_hi_lo_hi_hi_5 = {regroupV0_lo_hi_lo_hi_hi_hi_5, regroupV0_lo_hi_lo_hi_hi_lo_5};
  wire [511:0]       regroupV0_lo_hi_lo_hi_5 = {regroupV0_lo_hi_lo_hi_hi_5, regroupV0_lo_hi_lo_hi_lo_5};
  wire [1023:0]      regroupV0_lo_hi_lo_5 = {regroupV0_lo_hi_lo_hi_5, regroupV0_lo_hi_lo_lo_5};
  wire [127:0]       regroupV0_lo_hi_hi_lo_lo_lo_5 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_5, regroupV0_lo_hi_hi_lo_lo_lo_lo_5};
  wire [127:0]       regroupV0_lo_hi_hi_lo_lo_hi_5 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_5, regroupV0_lo_hi_hi_lo_lo_hi_lo_5};
  wire [255:0]       regroupV0_lo_hi_hi_lo_lo_5 = {regroupV0_lo_hi_hi_lo_lo_hi_5, regroupV0_lo_hi_hi_lo_lo_lo_5};
  wire [127:0]       regroupV0_lo_hi_hi_lo_hi_lo_5 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_5, regroupV0_lo_hi_hi_lo_hi_lo_lo_5};
  wire [127:0]       regroupV0_lo_hi_hi_lo_hi_hi_5 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_5, regroupV0_lo_hi_hi_lo_hi_hi_lo_5};
  wire [255:0]       regroupV0_lo_hi_hi_lo_hi_5 = {regroupV0_lo_hi_hi_lo_hi_hi_5, regroupV0_lo_hi_hi_lo_hi_lo_5};
  wire [511:0]       regroupV0_lo_hi_hi_lo_5 = {regroupV0_lo_hi_hi_lo_hi_5, regroupV0_lo_hi_hi_lo_lo_5};
  wire [127:0]       regroupV0_lo_hi_hi_hi_lo_lo_5 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_5, regroupV0_lo_hi_hi_hi_lo_lo_lo_5};
  wire [127:0]       regroupV0_lo_hi_hi_hi_lo_hi_5 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_5, regroupV0_lo_hi_hi_hi_lo_hi_lo_5};
  wire [255:0]       regroupV0_lo_hi_hi_hi_lo_5 = {regroupV0_lo_hi_hi_hi_lo_hi_5, regroupV0_lo_hi_hi_hi_lo_lo_5};
  wire [127:0]       regroupV0_lo_hi_hi_hi_hi_lo_5 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_5, regroupV0_lo_hi_hi_hi_hi_lo_lo_5};
  wire [127:0]       regroupV0_lo_hi_hi_hi_hi_hi_5 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_5, regroupV0_lo_hi_hi_hi_hi_hi_lo_5};
  wire [255:0]       regroupV0_lo_hi_hi_hi_hi_5 = {regroupV0_lo_hi_hi_hi_hi_hi_5, regroupV0_lo_hi_hi_hi_hi_lo_5};
  wire [511:0]       regroupV0_lo_hi_hi_hi_5 = {regroupV0_lo_hi_hi_hi_hi_5, regroupV0_lo_hi_hi_hi_lo_5};
  wire [1023:0]      regroupV0_lo_hi_hi_5 = {regroupV0_lo_hi_hi_hi_5, regroupV0_lo_hi_hi_lo_5};
  wire [2047:0]      regroupV0_lo_hi_5 = {regroupV0_lo_hi_hi_5, regroupV0_lo_hi_lo_5};
  wire [4095:0]      regroupV0_lo_6 = {regroupV0_lo_hi_5, regroupV0_lo_lo_5};
  wire [127:0]       regroupV0_hi_lo_lo_lo_lo_lo_5 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_5, regroupV0_hi_lo_lo_lo_lo_lo_lo_5};
  wire [127:0]       regroupV0_hi_lo_lo_lo_lo_hi_5 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_5, regroupV0_hi_lo_lo_lo_lo_hi_lo_5};
  wire [255:0]       regroupV0_hi_lo_lo_lo_lo_5 = {regroupV0_hi_lo_lo_lo_lo_hi_5, regroupV0_hi_lo_lo_lo_lo_lo_5};
  wire [127:0]       regroupV0_hi_lo_lo_lo_hi_lo_5 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_5, regroupV0_hi_lo_lo_lo_hi_lo_lo_5};
  wire [127:0]       regroupV0_hi_lo_lo_lo_hi_hi_5 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_5, regroupV0_hi_lo_lo_lo_hi_hi_lo_5};
  wire [255:0]       regroupV0_hi_lo_lo_lo_hi_5 = {regroupV0_hi_lo_lo_lo_hi_hi_5, regroupV0_hi_lo_lo_lo_hi_lo_5};
  wire [511:0]       regroupV0_hi_lo_lo_lo_5 = {regroupV0_hi_lo_lo_lo_hi_5, regroupV0_hi_lo_lo_lo_lo_5};
  wire [127:0]       regroupV0_hi_lo_lo_hi_lo_lo_5 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_5, regroupV0_hi_lo_lo_hi_lo_lo_lo_5};
  wire [127:0]       regroupV0_hi_lo_lo_hi_lo_hi_5 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_5, regroupV0_hi_lo_lo_hi_lo_hi_lo_5};
  wire [255:0]       regroupV0_hi_lo_lo_hi_lo_5 = {regroupV0_hi_lo_lo_hi_lo_hi_5, regroupV0_hi_lo_lo_hi_lo_lo_5};
  wire [127:0]       regroupV0_hi_lo_lo_hi_hi_lo_5 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_5, regroupV0_hi_lo_lo_hi_hi_lo_lo_5};
  wire [127:0]       regroupV0_hi_lo_lo_hi_hi_hi_5 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_5, regroupV0_hi_lo_lo_hi_hi_hi_lo_5};
  wire [255:0]       regroupV0_hi_lo_lo_hi_hi_5 = {regroupV0_hi_lo_lo_hi_hi_hi_5, regroupV0_hi_lo_lo_hi_hi_lo_5};
  wire [511:0]       regroupV0_hi_lo_lo_hi_5 = {regroupV0_hi_lo_lo_hi_hi_5, regroupV0_hi_lo_lo_hi_lo_5};
  wire [1023:0]      regroupV0_hi_lo_lo_5 = {regroupV0_hi_lo_lo_hi_5, regroupV0_hi_lo_lo_lo_5};
  wire [127:0]       regroupV0_hi_lo_hi_lo_lo_lo_5 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_5, regroupV0_hi_lo_hi_lo_lo_lo_lo_5};
  wire [127:0]       regroupV0_hi_lo_hi_lo_lo_hi_5 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_5, regroupV0_hi_lo_hi_lo_lo_hi_lo_5};
  wire [255:0]       regroupV0_hi_lo_hi_lo_lo_5 = {regroupV0_hi_lo_hi_lo_lo_hi_5, regroupV0_hi_lo_hi_lo_lo_lo_5};
  wire [127:0]       regroupV0_hi_lo_hi_lo_hi_lo_5 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_5, regroupV0_hi_lo_hi_lo_hi_lo_lo_5};
  wire [127:0]       regroupV0_hi_lo_hi_lo_hi_hi_5 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_5, regroupV0_hi_lo_hi_lo_hi_hi_lo_5};
  wire [255:0]       regroupV0_hi_lo_hi_lo_hi_5 = {regroupV0_hi_lo_hi_lo_hi_hi_5, regroupV0_hi_lo_hi_lo_hi_lo_5};
  wire [511:0]       regroupV0_hi_lo_hi_lo_5 = {regroupV0_hi_lo_hi_lo_hi_5, regroupV0_hi_lo_hi_lo_lo_5};
  wire [127:0]       regroupV0_hi_lo_hi_hi_lo_lo_5 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_5, regroupV0_hi_lo_hi_hi_lo_lo_lo_5};
  wire [127:0]       regroupV0_hi_lo_hi_hi_lo_hi_5 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_5, regroupV0_hi_lo_hi_hi_lo_hi_lo_5};
  wire [255:0]       regroupV0_hi_lo_hi_hi_lo_5 = {regroupV0_hi_lo_hi_hi_lo_hi_5, regroupV0_hi_lo_hi_hi_lo_lo_5};
  wire [127:0]       regroupV0_hi_lo_hi_hi_hi_lo_5 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_5, regroupV0_hi_lo_hi_hi_hi_lo_lo_5};
  wire [127:0]       regroupV0_hi_lo_hi_hi_hi_hi_5 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_5, regroupV0_hi_lo_hi_hi_hi_hi_lo_5};
  wire [255:0]       regroupV0_hi_lo_hi_hi_hi_5 = {regroupV0_hi_lo_hi_hi_hi_hi_5, regroupV0_hi_lo_hi_hi_hi_lo_5};
  wire [511:0]       regroupV0_hi_lo_hi_hi_5 = {regroupV0_hi_lo_hi_hi_hi_5, regroupV0_hi_lo_hi_hi_lo_5};
  wire [1023:0]      regroupV0_hi_lo_hi_5 = {regroupV0_hi_lo_hi_hi_5, regroupV0_hi_lo_hi_lo_5};
  wire [2047:0]      regroupV0_hi_lo_5 = {regroupV0_hi_lo_hi_5, regroupV0_hi_lo_lo_5};
  wire [127:0]       regroupV0_hi_hi_lo_lo_lo_lo_5 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_5, regroupV0_hi_hi_lo_lo_lo_lo_lo_5};
  wire [127:0]       regroupV0_hi_hi_lo_lo_lo_hi_5 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_5, regroupV0_hi_hi_lo_lo_lo_hi_lo_5};
  wire [255:0]       regroupV0_hi_hi_lo_lo_lo_5 = {regroupV0_hi_hi_lo_lo_lo_hi_5, regroupV0_hi_hi_lo_lo_lo_lo_5};
  wire [127:0]       regroupV0_hi_hi_lo_lo_hi_lo_5 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_5, regroupV0_hi_hi_lo_lo_hi_lo_lo_5};
  wire [127:0]       regroupV0_hi_hi_lo_lo_hi_hi_5 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_5, regroupV0_hi_hi_lo_lo_hi_hi_lo_5};
  wire [255:0]       regroupV0_hi_hi_lo_lo_hi_5 = {regroupV0_hi_hi_lo_lo_hi_hi_5, regroupV0_hi_hi_lo_lo_hi_lo_5};
  wire [511:0]       regroupV0_hi_hi_lo_lo_5 = {regroupV0_hi_hi_lo_lo_hi_5, regroupV0_hi_hi_lo_lo_lo_5};
  wire [127:0]       regroupV0_hi_hi_lo_hi_lo_lo_5 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_5, regroupV0_hi_hi_lo_hi_lo_lo_lo_5};
  wire [127:0]       regroupV0_hi_hi_lo_hi_lo_hi_5 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_5, regroupV0_hi_hi_lo_hi_lo_hi_lo_5};
  wire [255:0]       regroupV0_hi_hi_lo_hi_lo_5 = {regroupV0_hi_hi_lo_hi_lo_hi_5, regroupV0_hi_hi_lo_hi_lo_lo_5};
  wire [127:0]       regroupV0_hi_hi_lo_hi_hi_lo_5 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_5, regroupV0_hi_hi_lo_hi_hi_lo_lo_5};
  wire [127:0]       regroupV0_hi_hi_lo_hi_hi_hi_5 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_5, regroupV0_hi_hi_lo_hi_hi_hi_lo_5};
  wire [255:0]       regroupV0_hi_hi_lo_hi_hi_5 = {regroupV0_hi_hi_lo_hi_hi_hi_5, regroupV0_hi_hi_lo_hi_hi_lo_5};
  wire [511:0]       regroupV0_hi_hi_lo_hi_5 = {regroupV0_hi_hi_lo_hi_hi_5, regroupV0_hi_hi_lo_hi_lo_5};
  wire [1023:0]      regroupV0_hi_hi_lo_5 = {regroupV0_hi_hi_lo_hi_5, regroupV0_hi_hi_lo_lo_5};
  wire [127:0]       regroupV0_hi_hi_hi_lo_lo_lo_5 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_5, regroupV0_hi_hi_hi_lo_lo_lo_lo_5};
  wire [127:0]       regroupV0_hi_hi_hi_lo_lo_hi_5 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_5, regroupV0_hi_hi_hi_lo_lo_hi_lo_5};
  wire [255:0]       regroupV0_hi_hi_hi_lo_lo_5 = {regroupV0_hi_hi_hi_lo_lo_hi_5, regroupV0_hi_hi_hi_lo_lo_lo_5};
  wire [127:0]       regroupV0_hi_hi_hi_lo_hi_lo_5 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_5, regroupV0_hi_hi_hi_lo_hi_lo_lo_5};
  wire [127:0]       regroupV0_hi_hi_hi_lo_hi_hi_5 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_5, regroupV0_hi_hi_hi_lo_hi_hi_lo_5};
  wire [255:0]       regroupV0_hi_hi_hi_lo_hi_5 = {regroupV0_hi_hi_hi_lo_hi_hi_5, regroupV0_hi_hi_hi_lo_hi_lo_5};
  wire [511:0]       regroupV0_hi_hi_hi_lo_5 = {regroupV0_hi_hi_hi_lo_hi_5, regroupV0_hi_hi_hi_lo_lo_5};
  wire [127:0]       regroupV0_hi_hi_hi_hi_lo_lo_5 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_5, regroupV0_hi_hi_hi_hi_lo_lo_lo_5};
  wire [127:0]       regroupV0_hi_hi_hi_hi_lo_hi_5 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_5, regroupV0_hi_hi_hi_hi_lo_hi_lo_5};
  wire [255:0]       regroupV0_hi_hi_hi_hi_lo_5 = {regroupV0_hi_hi_hi_hi_lo_hi_5, regroupV0_hi_hi_hi_hi_lo_lo_5};
  wire [127:0]       regroupV0_hi_hi_hi_hi_hi_lo_5 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_5, regroupV0_hi_hi_hi_hi_hi_lo_lo_5};
  wire [127:0]       regroupV0_hi_hi_hi_hi_hi_hi_5 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_5, regroupV0_hi_hi_hi_hi_hi_hi_lo_5};
  wire [255:0]       regroupV0_hi_hi_hi_hi_hi_5 = {regroupV0_hi_hi_hi_hi_hi_hi_5, regroupV0_hi_hi_hi_hi_hi_lo_5};
  wire [511:0]       regroupV0_hi_hi_hi_hi_5 = {regroupV0_hi_hi_hi_hi_hi_5, regroupV0_hi_hi_hi_hi_lo_5};
  wire [1023:0]      regroupV0_hi_hi_hi_5 = {regroupV0_hi_hi_hi_hi_5, regroupV0_hi_hi_hi_lo_5};
  wire [2047:0]      regroupV0_hi_hi_5 = {regroupV0_hi_hi_hi_5, regroupV0_hi_hi_lo_5};
  wire [4095:0]      regroupV0_hi_6 = {regroupV0_hi_hi_5, regroupV0_hi_lo_5};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo = {regroupV0_lo_6[9:8], regroupV0_lo_6[1:0]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi = {regroupV0_lo_6[25:24], regroupV0_lo_6[17:16]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_4 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo = {regroupV0_lo_6[41:40], regroupV0_lo_6[33:32]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi = {regroupV0_lo_6[57:56], regroupV0_lo_6[49:48]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_4 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi, regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_lo_lo_6 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_4, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_4};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo = {regroupV0_lo_6[73:72], regroupV0_lo_6[65:64]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi = {regroupV0_lo_6[89:88], regroupV0_lo_6[81:80]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_4 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo = {regroupV0_lo_6[105:104], regroupV0_lo_6[97:96]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi = {regroupV0_lo_6[121:120], regroupV0_lo_6[113:112]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_4 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi, regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_lo_hi_6 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_4, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_4};
  wire [31:0]        regroupV0_lo_lo_lo_lo_lo_lo_6 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_6, regroupV0_lo_lo_lo_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo = {regroupV0_lo_6[137:136], regroupV0_lo_6[129:128]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi = {regroupV0_lo_6[153:152], regroupV0_lo_6[145:144]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_4 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo = {regroupV0_lo_6[169:168], regroupV0_lo_6[161:160]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi = {regroupV0_lo_6[185:184], regroupV0_lo_6[177:176]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_4 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi, regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_hi_lo_6 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_4, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_4};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo = {regroupV0_lo_6[201:200], regroupV0_lo_6[193:192]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi = {regroupV0_lo_6[217:216], regroupV0_lo_6[209:208]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_4 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo = {regroupV0_lo_6[233:232], regroupV0_lo_6[225:224]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi = {regroupV0_lo_6[249:248], regroupV0_lo_6[241:240]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_4 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi, regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_hi_hi_6 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_4, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_4};
  wire [31:0]        regroupV0_lo_lo_lo_lo_lo_hi_6 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_6, regroupV0_lo_lo_lo_lo_lo_hi_lo_6};
  wire [63:0]        regroupV0_lo_lo_lo_lo_lo_6 = {regroupV0_lo_lo_lo_lo_lo_hi_6, regroupV0_lo_lo_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo = {regroupV0_lo_6[265:264], regroupV0_lo_6[257:256]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi = {regroupV0_lo_6[281:280], regroupV0_lo_6[273:272]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_4 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo = {regroupV0_lo_6[297:296], regroupV0_lo_6[289:288]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi = {regroupV0_lo_6[313:312], regroupV0_lo_6[305:304]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_4 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi, regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_lo_lo_6 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_4, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_4};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo = {regroupV0_lo_6[329:328], regroupV0_lo_6[321:320]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi = {regroupV0_lo_6[345:344], regroupV0_lo_6[337:336]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_4 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo = {regroupV0_lo_6[361:360], regroupV0_lo_6[353:352]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi = {regroupV0_lo_6[377:376], regroupV0_lo_6[369:368]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_4 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi, regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_lo_hi_6 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_4, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_4};
  wire [31:0]        regroupV0_lo_lo_lo_lo_hi_lo_6 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_6, regroupV0_lo_lo_lo_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo = {regroupV0_lo_6[393:392], regroupV0_lo_6[385:384]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi = {regroupV0_lo_6[409:408], regroupV0_lo_6[401:400]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_4 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo = {regroupV0_lo_6[425:424], regroupV0_lo_6[417:416]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi = {regroupV0_lo_6[441:440], regroupV0_lo_6[433:432]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_4 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi, regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_hi_lo_6 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_4, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_4};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo = {regroupV0_lo_6[457:456], regroupV0_lo_6[449:448]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi = {regroupV0_lo_6[473:472], regroupV0_lo_6[465:464]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_4 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo = {regroupV0_lo_6[489:488], regroupV0_lo_6[481:480]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi = {regroupV0_lo_6[505:504], regroupV0_lo_6[497:496]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_4 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi, regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_hi_hi_6 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_4, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_4};
  wire [31:0]        regroupV0_lo_lo_lo_lo_hi_hi_6 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_6, regroupV0_lo_lo_lo_lo_hi_hi_lo_6};
  wire [63:0]        regroupV0_lo_lo_lo_lo_hi_6 = {regroupV0_lo_lo_lo_lo_hi_hi_6, regroupV0_lo_lo_lo_lo_hi_lo_6};
  wire [127:0]       regroupV0_lo_lo_lo_lo_6 = {regroupV0_lo_lo_lo_lo_hi_6, regroupV0_lo_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo = {regroupV0_lo_6[521:520], regroupV0_lo_6[513:512]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi = {regroupV0_lo_6[537:536], regroupV0_lo_6[529:528]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_4 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo = {regroupV0_lo_6[553:552], regroupV0_lo_6[545:544]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi = {regroupV0_lo_6[569:568], regroupV0_lo_6[561:560]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_4 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi, regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_lo_lo_6 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_4, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_4};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo = {regroupV0_lo_6[585:584], regroupV0_lo_6[577:576]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi = {regroupV0_lo_6[601:600], regroupV0_lo_6[593:592]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_4 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo = {regroupV0_lo_6[617:616], regroupV0_lo_6[609:608]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi = {regroupV0_lo_6[633:632], regroupV0_lo_6[625:624]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_4 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi, regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_lo_hi_6 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_4, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_4};
  wire [31:0]        regroupV0_lo_lo_lo_hi_lo_lo_6 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_6, regroupV0_lo_lo_lo_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo = {regroupV0_lo_6[649:648], regroupV0_lo_6[641:640]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi = {regroupV0_lo_6[665:664], regroupV0_lo_6[657:656]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_4 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo = {regroupV0_lo_6[681:680], regroupV0_lo_6[673:672]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi = {regroupV0_lo_6[697:696], regroupV0_lo_6[689:688]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_4 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi, regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_hi_lo_6 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_4, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_4};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo = {regroupV0_lo_6[713:712], regroupV0_lo_6[705:704]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi = {regroupV0_lo_6[729:728], regroupV0_lo_6[721:720]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_4 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo = {regroupV0_lo_6[745:744], regroupV0_lo_6[737:736]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi = {regroupV0_lo_6[761:760], regroupV0_lo_6[753:752]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_4 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi, regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_hi_hi_6 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_4, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_4};
  wire [31:0]        regroupV0_lo_lo_lo_hi_lo_hi_6 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_6, regroupV0_lo_lo_lo_hi_lo_hi_lo_6};
  wire [63:0]        regroupV0_lo_lo_lo_hi_lo_6 = {regroupV0_lo_lo_lo_hi_lo_hi_6, regroupV0_lo_lo_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo = {regroupV0_lo_6[777:776], regroupV0_lo_6[769:768]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi = {regroupV0_lo_6[793:792], regroupV0_lo_6[785:784]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_4 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo = {regroupV0_lo_6[809:808], regroupV0_lo_6[801:800]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi = {regroupV0_lo_6[825:824], regroupV0_lo_6[817:816]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_4 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi, regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_lo_lo_6 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_4, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_4};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo = {regroupV0_lo_6[841:840], regroupV0_lo_6[833:832]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi = {regroupV0_lo_6[857:856], regroupV0_lo_6[849:848]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_4 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo = {regroupV0_lo_6[873:872], regroupV0_lo_6[865:864]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi = {regroupV0_lo_6[889:888], regroupV0_lo_6[881:880]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_4 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi, regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_lo_hi_6 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_4, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_4};
  wire [31:0]        regroupV0_lo_lo_lo_hi_hi_lo_6 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_6, regroupV0_lo_lo_lo_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo = {regroupV0_lo_6[905:904], regroupV0_lo_6[897:896]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi = {regroupV0_lo_6[921:920], regroupV0_lo_6[913:912]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_4 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo = {regroupV0_lo_6[937:936], regroupV0_lo_6[929:928]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi = {regroupV0_lo_6[953:952], regroupV0_lo_6[945:944]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_4 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi, regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_hi_lo_6 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_4, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_4};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo = {regroupV0_lo_6[969:968], regroupV0_lo_6[961:960]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi = {regroupV0_lo_6[985:984], regroupV0_lo_6[977:976]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_4 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo = {regroupV0_lo_6[1001:1000], regroupV0_lo_6[993:992]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi = {regroupV0_lo_6[1017:1016], regroupV0_lo_6[1009:1008]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_4 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi, regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_hi_hi_6 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_4, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_4};
  wire [31:0]        regroupV0_lo_lo_lo_hi_hi_hi_6 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_6, regroupV0_lo_lo_lo_hi_hi_hi_lo_6};
  wire [63:0]        regroupV0_lo_lo_lo_hi_hi_6 = {regroupV0_lo_lo_lo_hi_hi_hi_6, regroupV0_lo_lo_lo_hi_hi_lo_6};
  wire [127:0]       regroupV0_lo_lo_lo_hi_6 = {regroupV0_lo_lo_lo_hi_hi_6, regroupV0_lo_lo_lo_hi_lo_6};
  wire [255:0]       regroupV0_lo_lo_lo_6 = {regroupV0_lo_lo_lo_hi_6, regroupV0_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo = {regroupV0_lo_6[1033:1032], regroupV0_lo_6[1025:1024]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi = {regroupV0_lo_6[1049:1048], regroupV0_lo_6[1041:1040]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_4 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo = {regroupV0_lo_6[1065:1064], regroupV0_lo_6[1057:1056]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi = {regroupV0_lo_6[1081:1080], regroupV0_lo_6[1073:1072]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_4 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi, regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_lo_lo_6 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_4, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_4};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo = {regroupV0_lo_6[1097:1096], regroupV0_lo_6[1089:1088]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi = {regroupV0_lo_6[1113:1112], regroupV0_lo_6[1105:1104]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_4 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo = {regroupV0_lo_6[1129:1128], regroupV0_lo_6[1121:1120]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi = {regroupV0_lo_6[1145:1144], regroupV0_lo_6[1137:1136]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_4 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi, regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_lo_hi_6 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_4, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_4};
  wire [31:0]        regroupV0_lo_lo_hi_lo_lo_lo_6 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_6, regroupV0_lo_lo_hi_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo = {regroupV0_lo_6[1161:1160], regroupV0_lo_6[1153:1152]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi = {regroupV0_lo_6[1177:1176], regroupV0_lo_6[1169:1168]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_4 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo = {regroupV0_lo_6[1193:1192], regroupV0_lo_6[1185:1184]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi = {regroupV0_lo_6[1209:1208], regroupV0_lo_6[1201:1200]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_4 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi, regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_hi_lo_6 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_4, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_4};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo = {regroupV0_lo_6[1225:1224], regroupV0_lo_6[1217:1216]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi = {regroupV0_lo_6[1241:1240], regroupV0_lo_6[1233:1232]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_4 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo = {regroupV0_lo_6[1257:1256], regroupV0_lo_6[1249:1248]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi = {regroupV0_lo_6[1273:1272], regroupV0_lo_6[1265:1264]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_4 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi, regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_hi_hi_6 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_4, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_4};
  wire [31:0]        regroupV0_lo_lo_hi_lo_lo_hi_6 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_6, regroupV0_lo_lo_hi_lo_lo_hi_lo_6};
  wire [63:0]        regroupV0_lo_lo_hi_lo_lo_6 = {regroupV0_lo_lo_hi_lo_lo_hi_6, regroupV0_lo_lo_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo = {regroupV0_lo_6[1289:1288], regroupV0_lo_6[1281:1280]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi = {regroupV0_lo_6[1305:1304], regroupV0_lo_6[1297:1296]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_4 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo = {regroupV0_lo_6[1321:1320], regroupV0_lo_6[1313:1312]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi = {regroupV0_lo_6[1337:1336], regroupV0_lo_6[1329:1328]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_4 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi, regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_lo_lo_6 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_4, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_4};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo = {regroupV0_lo_6[1353:1352], regroupV0_lo_6[1345:1344]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi = {regroupV0_lo_6[1369:1368], regroupV0_lo_6[1361:1360]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_4 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo = {regroupV0_lo_6[1385:1384], regroupV0_lo_6[1377:1376]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi = {regroupV0_lo_6[1401:1400], regroupV0_lo_6[1393:1392]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_4 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi, regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_lo_hi_6 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_4, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_4};
  wire [31:0]        regroupV0_lo_lo_hi_lo_hi_lo_6 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_6, regroupV0_lo_lo_hi_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo = {regroupV0_lo_6[1417:1416], regroupV0_lo_6[1409:1408]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi = {regroupV0_lo_6[1433:1432], regroupV0_lo_6[1425:1424]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_4 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo = {regroupV0_lo_6[1449:1448], regroupV0_lo_6[1441:1440]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi = {regroupV0_lo_6[1465:1464], regroupV0_lo_6[1457:1456]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_4 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi, regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_hi_lo_6 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_4, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_4};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo = {regroupV0_lo_6[1481:1480], regroupV0_lo_6[1473:1472]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi = {regroupV0_lo_6[1497:1496], regroupV0_lo_6[1489:1488]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_4 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo = {regroupV0_lo_6[1513:1512], regroupV0_lo_6[1505:1504]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi = {regroupV0_lo_6[1529:1528], regroupV0_lo_6[1521:1520]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_4 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi, regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_hi_hi_6 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_4, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_4};
  wire [31:0]        regroupV0_lo_lo_hi_lo_hi_hi_6 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_6, regroupV0_lo_lo_hi_lo_hi_hi_lo_6};
  wire [63:0]        regroupV0_lo_lo_hi_lo_hi_6 = {regroupV0_lo_lo_hi_lo_hi_hi_6, regroupV0_lo_lo_hi_lo_hi_lo_6};
  wire [127:0]       regroupV0_lo_lo_hi_lo_6 = {regroupV0_lo_lo_hi_lo_hi_6, regroupV0_lo_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo = {regroupV0_lo_6[1545:1544], regroupV0_lo_6[1537:1536]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi = {regroupV0_lo_6[1561:1560], regroupV0_lo_6[1553:1552]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_4 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo = {regroupV0_lo_6[1577:1576], regroupV0_lo_6[1569:1568]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi = {regroupV0_lo_6[1593:1592], regroupV0_lo_6[1585:1584]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_4 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi, regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_lo_lo_6 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_4, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_4};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo = {regroupV0_lo_6[1609:1608], regroupV0_lo_6[1601:1600]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi = {regroupV0_lo_6[1625:1624], regroupV0_lo_6[1617:1616]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_4 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo = {regroupV0_lo_6[1641:1640], regroupV0_lo_6[1633:1632]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi = {regroupV0_lo_6[1657:1656], regroupV0_lo_6[1649:1648]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_4 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi, regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_lo_hi_6 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_4, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_4};
  wire [31:0]        regroupV0_lo_lo_hi_hi_lo_lo_6 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_6, regroupV0_lo_lo_hi_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo = {regroupV0_lo_6[1673:1672], regroupV0_lo_6[1665:1664]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi = {regroupV0_lo_6[1689:1688], regroupV0_lo_6[1681:1680]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_4 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo = {regroupV0_lo_6[1705:1704], regroupV0_lo_6[1697:1696]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi = {regroupV0_lo_6[1721:1720], regroupV0_lo_6[1713:1712]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_4 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi, regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_hi_lo_6 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_4, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_4};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo = {regroupV0_lo_6[1737:1736], regroupV0_lo_6[1729:1728]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi = {regroupV0_lo_6[1753:1752], regroupV0_lo_6[1745:1744]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_4 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo = {regroupV0_lo_6[1769:1768], regroupV0_lo_6[1761:1760]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi = {regroupV0_lo_6[1785:1784], regroupV0_lo_6[1777:1776]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_4 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi, regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_hi_hi_6 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_4, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_4};
  wire [31:0]        regroupV0_lo_lo_hi_hi_lo_hi_6 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_6, regroupV0_lo_lo_hi_hi_lo_hi_lo_6};
  wire [63:0]        regroupV0_lo_lo_hi_hi_lo_6 = {regroupV0_lo_lo_hi_hi_lo_hi_6, regroupV0_lo_lo_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo = {regroupV0_lo_6[1801:1800], regroupV0_lo_6[1793:1792]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi = {regroupV0_lo_6[1817:1816], regroupV0_lo_6[1809:1808]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_4 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo = {regroupV0_lo_6[1833:1832], regroupV0_lo_6[1825:1824]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi = {regroupV0_lo_6[1849:1848], regroupV0_lo_6[1841:1840]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_4 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi, regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_lo_lo_6 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_4, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_4};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo = {regroupV0_lo_6[1865:1864], regroupV0_lo_6[1857:1856]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi = {regroupV0_lo_6[1881:1880], regroupV0_lo_6[1873:1872]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_4 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo = {regroupV0_lo_6[1897:1896], regroupV0_lo_6[1889:1888]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi = {regroupV0_lo_6[1913:1912], regroupV0_lo_6[1905:1904]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_4 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi, regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_lo_hi_6 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_4, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_4};
  wire [31:0]        regroupV0_lo_lo_hi_hi_hi_lo_6 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_6, regroupV0_lo_lo_hi_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo = {regroupV0_lo_6[1929:1928], regroupV0_lo_6[1921:1920]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi = {regroupV0_lo_6[1945:1944], regroupV0_lo_6[1937:1936]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_4 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo = {regroupV0_lo_6[1961:1960], regroupV0_lo_6[1953:1952]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi = {regroupV0_lo_6[1977:1976], regroupV0_lo_6[1969:1968]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_4 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi, regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_hi_lo_6 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_4, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_4};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo = {regroupV0_lo_6[1993:1992], regroupV0_lo_6[1985:1984]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi = {regroupV0_lo_6[2009:2008], regroupV0_lo_6[2001:2000]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_4 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo = {regroupV0_lo_6[2025:2024], regroupV0_lo_6[2017:2016]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi = {regroupV0_lo_6[2041:2040], regroupV0_lo_6[2033:2032]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_4 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi, regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_hi_hi_6 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_4, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_4};
  wire [31:0]        regroupV0_lo_lo_hi_hi_hi_hi_6 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_6, regroupV0_lo_lo_hi_hi_hi_hi_lo_6};
  wire [63:0]        regroupV0_lo_lo_hi_hi_hi_6 = {regroupV0_lo_lo_hi_hi_hi_hi_6, regroupV0_lo_lo_hi_hi_hi_lo_6};
  wire [127:0]       regroupV0_lo_lo_hi_hi_6 = {regroupV0_lo_lo_hi_hi_hi_6, regroupV0_lo_lo_hi_hi_lo_6};
  wire [255:0]       regroupV0_lo_lo_hi_6 = {regroupV0_lo_lo_hi_hi_6, regroupV0_lo_lo_hi_lo_6};
  wire [511:0]       regroupV0_lo_lo_6 = {regroupV0_lo_lo_hi_6, regroupV0_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo = {regroupV0_lo_6[2057:2056], regroupV0_lo_6[2049:2048]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi = {regroupV0_lo_6[2073:2072], regroupV0_lo_6[2065:2064]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_4 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo = {regroupV0_lo_6[2089:2088], regroupV0_lo_6[2081:2080]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi = {regroupV0_lo_6[2105:2104], regroupV0_lo_6[2097:2096]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_4 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi, regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_lo_lo_6 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_4, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_4};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo = {regroupV0_lo_6[2121:2120], regroupV0_lo_6[2113:2112]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi = {regroupV0_lo_6[2137:2136], regroupV0_lo_6[2129:2128]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_4 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo = {regroupV0_lo_6[2153:2152], regroupV0_lo_6[2145:2144]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi = {regroupV0_lo_6[2169:2168], regroupV0_lo_6[2161:2160]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_4 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi, regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_lo_hi_6 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_4, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_4};
  wire [31:0]        regroupV0_lo_hi_lo_lo_lo_lo_6 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_6, regroupV0_lo_hi_lo_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo = {regroupV0_lo_6[2185:2184], regroupV0_lo_6[2177:2176]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi = {regroupV0_lo_6[2201:2200], regroupV0_lo_6[2193:2192]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_4 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo = {regroupV0_lo_6[2217:2216], regroupV0_lo_6[2209:2208]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi = {regroupV0_lo_6[2233:2232], regroupV0_lo_6[2225:2224]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_4 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi, regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_hi_lo_6 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_4, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_4};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo = {regroupV0_lo_6[2249:2248], regroupV0_lo_6[2241:2240]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi = {regroupV0_lo_6[2265:2264], regroupV0_lo_6[2257:2256]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_4 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo = {regroupV0_lo_6[2281:2280], regroupV0_lo_6[2273:2272]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi = {regroupV0_lo_6[2297:2296], regroupV0_lo_6[2289:2288]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_4 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi, regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_hi_hi_6 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_4, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_4};
  wire [31:0]        regroupV0_lo_hi_lo_lo_lo_hi_6 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_6, regroupV0_lo_hi_lo_lo_lo_hi_lo_6};
  wire [63:0]        regroupV0_lo_hi_lo_lo_lo_6 = {regroupV0_lo_hi_lo_lo_lo_hi_6, regroupV0_lo_hi_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo = {regroupV0_lo_6[2313:2312], regroupV0_lo_6[2305:2304]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi = {regroupV0_lo_6[2329:2328], regroupV0_lo_6[2321:2320]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_4 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo = {regroupV0_lo_6[2345:2344], regroupV0_lo_6[2337:2336]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi = {regroupV0_lo_6[2361:2360], regroupV0_lo_6[2353:2352]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_4 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi, regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_lo_lo_6 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_4, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_4};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo = {regroupV0_lo_6[2377:2376], regroupV0_lo_6[2369:2368]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi = {regroupV0_lo_6[2393:2392], regroupV0_lo_6[2385:2384]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_4 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo = {regroupV0_lo_6[2409:2408], regroupV0_lo_6[2401:2400]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi = {regroupV0_lo_6[2425:2424], regroupV0_lo_6[2417:2416]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_4 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi, regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_lo_hi_6 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_4, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_4};
  wire [31:0]        regroupV0_lo_hi_lo_lo_hi_lo_6 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_6, regroupV0_lo_hi_lo_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo = {regroupV0_lo_6[2441:2440], regroupV0_lo_6[2433:2432]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi = {regroupV0_lo_6[2457:2456], regroupV0_lo_6[2449:2448]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_4 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo = {regroupV0_lo_6[2473:2472], regroupV0_lo_6[2465:2464]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi = {regroupV0_lo_6[2489:2488], regroupV0_lo_6[2481:2480]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_4 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi, regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_hi_lo_6 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_4, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_4};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo = {regroupV0_lo_6[2505:2504], regroupV0_lo_6[2497:2496]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi = {regroupV0_lo_6[2521:2520], regroupV0_lo_6[2513:2512]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_4 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo = {regroupV0_lo_6[2537:2536], regroupV0_lo_6[2529:2528]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi = {regroupV0_lo_6[2553:2552], regroupV0_lo_6[2545:2544]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_4 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi, regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_hi_hi_6 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_4, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_4};
  wire [31:0]        regroupV0_lo_hi_lo_lo_hi_hi_6 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_6, regroupV0_lo_hi_lo_lo_hi_hi_lo_6};
  wire [63:0]        regroupV0_lo_hi_lo_lo_hi_6 = {regroupV0_lo_hi_lo_lo_hi_hi_6, regroupV0_lo_hi_lo_lo_hi_lo_6};
  wire [127:0]       regroupV0_lo_hi_lo_lo_6 = {regroupV0_lo_hi_lo_lo_hi_6, regroupV0_lo_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo = {regroupV0_lo_6[2569:2568], regroupV0_lo_6[2561:2560]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi = {regroupV0_lo_6[2585:2584], regroupV0_lo_6[2577:2576]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_4 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo = {regroupV0_lo_6[2601:2600], regroupV0_lo_6[2593:2592]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi = {regroupV0_lo_6[2617:2616], regroupV0_lo_6[2609:2608]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_4 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi, regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_lo_lo_6 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_4, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_4};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo = {regroupV0_lo_6[2633:2632], regroupV0_lo_6[2625:2624]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi = {regroupV0_lo_6[2649:2648], regroupV0_lo_6[2641:2640]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_4 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo = {regroupV0_lo_6[2665:2664], regroupV0_lo_6[2657:2656]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi = {regroupV0_lo_6[2681:2680], regroupV0_lo_6[2673:2672]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_4 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi, regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_lo_hi_6 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_4, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_4};
  wire [31:0]        regroupV0_lo_hi_lo_hi_lo_lo_6 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_6, regroupV0_lo_hi_lo_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo = {regroupV0_lo_6[2697:2696], regroupV0_lo_6[2689:2688]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi = {regroupV0_lo_6[2713:2712], regroupV0_lo_6[2705:2704]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_4 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo = {regroupV0_lo_6[2729:2728], regroupV0_lo_6[2721:2720]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi = {regroupV0_lo_6[2745:2744], regroupV0_lo_6[2737:2736]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_4 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi, regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_hi_lo_6 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_4, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_4};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo = {regroupV0_lo_6[2761:2760], regroupV0_lo_6[2753:2752]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi = {regroupV0_lo_6[2777:2776], regroupV0_lo_6[2769:2768]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_4 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo = {regroupV0_lo_6[2793:2792], regroupV0_lo_6[2785:2784]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi = {regroupV0_lo_6[2809:2808], regroupV0_lo_6[2801:2800]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_4 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi, regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_hi_hi_6 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_4, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_4};
  wire [31:0]        regroupV0_lo_hi_lo_hi_lo_hi_6 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_6, regroupV0_lo_hi_lo_hi_lo_hi_lo_6};
  wire [63:0]        regroupV0_lo_hi_lo_hi_lo_6 = {regroupV0_lo_hi_lo_hi_lo_hi_6, regroupV0_lo_hi_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo = {regroupV0_lo_6[2825:2824], regroupV0_lo_6[2817:2816]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi = {regroupV0_lo_6[2841:2840], regroupV0_lo_6[2833:2832]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_4 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo = {regroupV0_lo_6[2857:2856], regroupV0_lo_6[2849:2848]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi = {regroupV0_lo_6[2873:2872], regroupV0_lo_6[2865:2864]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_4 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi, regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_lo_lo_6 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_4, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_4};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo = {regroupV0_lo_6[2889:2888], regroupV0_lo_6[2881:2880]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi = {regroupV0_lo_6[2905:2904], regroupV0_lo_6[2897:2896]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_4 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo = {regroupV0_lo_6[2921:2920], regroupV0_lo_6[2913:2912]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi = {regroupV0_lo_6[2937:2936], regroupV0_lo_6[2929:2928]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_4 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi, regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_lo_hi_6 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_4, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_4};
  wire [31:0]        regroupV0_lo_hi_lo_hi_hi_lo_6 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_6, regroupV0_lo_hi_lo_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo = {regroupV0_lo_6[2953:2952], regroupV0_lo_6[2945:2944]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi = {regroupV0_lo_6[2969:2968], regroupV0_lo_6[2961:2960]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_4 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo = {regroupV0_lo_6[2985:2984], regroupV0_lo_6[2977:2976]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi = {regroupV0_lo_6[3001:3000], regroupV0_lo_6[2993:2992]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_4 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi, regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_hi_lo_6 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_4, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_4};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo = {regroupV0_lo_6[3017:3016], regroupV0_lo_6[3009:3008]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi = {regroupV0_lo_6[3033:3032], regroupV0_lo_6[3025:3024]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_4 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo = {regroupV0_lo_6[3049:3048], regroupV0_lo_6[3041:3040]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi = {regroupV0_lo_6[3065:3064], regroupV0_lo_6[3057:3056]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_4 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi, regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_hi_hi_6 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_4, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_4};
  wire [31:0]        regroupV0_lo_hi_lo_hi_hi_hi_6 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_6, regroupV0_lo_hi_lo_hi_hi_hi_lo_6};
  wire [63:0]        regroupV0_lo_hi_lo_hi_hi_6 = {regroupV0_lo_hi_lo_hi_hi_hi_6, regroupV0_lo_hi_lo_hi_hi_lo_6};
  wire [127:0]       regroupV0_lo_hi_lo_hi_6 = {regroupV0_lo_hi_lo_hi_hi_6, regroupV0_lo_hi_lo_hi_lo_6};
  wire [255:0]       regroupV0_lo_hi_lo_6 = {regroupV0_lo_hi_lo_hi_6, regroupV0_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo = {regroupV0_lo_6[3081:3080], regroupV0_lo_6[3073:3072]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi = {regroupV0_lo_6[3097:3096], regroupV0_lo_6[3089:3088]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_4 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo = {regroupV0_lo_6[3113:3112], regroupV0_lo_6[3105:3104]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi = {regroupV0_lo_6[3129:3128], regroupV0_lo_6[3121:3120]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_4 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi, regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_lo_lo_6 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_4, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_4};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo = {regroupV0_lo_6[3145:3144], regroupV0_lo_6[3137:3136]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi = {regroupV0_lo_6[3161:3160], regroupV0_lo_6[3153:3152]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_4 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo = {regroupV0_lo_6[3177:3176], regroupV0_lo_6[3169:3168]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi = {regroupV0_lo_6[3193:3192], regroupV0_lo_6[3185:3184]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_4 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi, regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_lo_hi_6 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_4, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_4};
  wire [31:0]        regroupV0_lo_hi_hi_lo_lo_lo_6 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_6, regroupV0_lo_hi_hi_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo = {regroupV0_lo_6[3209:3208], regroupV0_lo_6[3201:3200]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi = {regroupV0_lo_6[3225:3224], regroupV0_lo_6[3217:3216]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_4 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo = {regroupV0_lo_6[3241:3240], regroupV0_lo_6[3233:3232]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi = {regroupV0_lo_6[3257:3256], regroupV0_lo_6[3249:3248]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_4 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi, regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_hi_lo_6 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_4, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_4};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo = {regroupV0_lo_6[3273:3272], regroupV0_lo_6[3265:3264]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi = {regroupV0_lo_6[3289:3288], regroupV0_lo_6[3281:3280]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_4 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo = {regroupV0_lo_6[3305:3304], regroupV0_lo_6[3297:3296]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi = {regroupV0_lo_6[3321:3320], regroupV0_lo_6[3313:3312]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_4 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi, regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_hi_hi_6 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_4, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_4};
  wire [31:0]        regroupV0_lo_hi_hi_lo_lo_hi_6 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_6, regroupV0_lo_hi_hi_lo_lo_hi_lo_6};
  wire [63:0]        regroupV0_lo_hi_hi_lo_lo_6 = {regroupV0_lo_hi_hi_lo_lo_hi_6, regroupV0_lo_hi_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo = {regroupV0_lo_6[3337:3336], regroupV0_lo_6[3329:3328]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi = {regroupV0_lo_6[3353:3352], regroupV0_lo_6[3345:3344]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_4 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo = {regroupV0_lo_6[3369:3368], regroupV0_lo_6[3361:3360]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi = {regroupV0_lo_6[3385:3384], regroupV0_lo_6[3377:3376]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_4 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi, regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_lo_lo_6 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_4, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_4};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo = {regroupV0_lo_6[3401:3400], regroupV0_lo_6[3393:3392]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi = {regroupV0_lo_6[3417:3416], regroupV0_lo_6[3409:3408]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_4 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo = {regroupV0_lo_6[3433:3432], regroupV0_lo_6[3425:3424]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi = {regroupV0_lo_6[3449:3448], regroupV0_lo_6[3441:3440]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_4 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi, regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_lo_hi_6 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_4, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_4};
  wire [31:0]        regroupV0_lo_hi_hi_lo_hi_lo_6 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_6, regroupV0_lo_hi_hi_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo = {regroupV0_lo_6[3465:3464], regroupV0_lo_6[3457:3456]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi = {regroupV0_lo_6[3481:3480], regroupV0_lo_6[3473:3472]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_4 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo = {regroupV0_lo_6[3497:3496], regroupV0_lo_6[3489:3488]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi = {regroupV0_lo_6[3513:3512], regroupV0_lo_6[3505:3504]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_4 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi, regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_hi_lo_6 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_4, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_4};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo = {regroupV0_lo_6[3529:3528], regroupV0_lo_6[3521:3520]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi = {regroupV0_lo_6[3545:3544], regroupV0_lo_6[3537:3536]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_4 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo = {regroupV0_lo_6[3561:3560], regroupV0_lo_6[3553:3552]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi = {regroupV0_lo_6[3577:3576], regroupV0_lo_6[3569:3568]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_4 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi, regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_hi_hi_6 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_4, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_4};
  wire [31:0]        regroupV0_lo_hi_hi_lo_hi_hi_6 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_6, regroupV0_lo_hi_hi_lo_hi_hi_lo_6};
  wire [63:0]        regroupV0_lo_hi_hi_lo_hi_6 = {regroupV0_lo_hi_hi_lo_hi_hi_6, regroupV0_lo_hi_hi_lo_hi_lo_6};
  wire [127:0]       regroupV0_lo_hi_hi_lo_6 = {regroupV0_lo_hi_hi_lo_hi_6, regroupV0_lo_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo = {regroupV0_lo_6[3593:3592], regroupV0_lo_6[3585:3584]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi = {regroupV0_lo_6[3609:3608], regroupV0_lo_6[3601:3600]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_4 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo = {regroupV0_lo_6[3625:3624], regroupV0_lo_6[3617:3616]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi = {regroupV0_lo_6[3641:3640], regroupV0_lo_6[3633:3632]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_4 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi, regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_lo_lo_6 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_4, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_4};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo = {regroupV0_lo_6[3657:3656], regroupV0_lo_6[3649:3648]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi = {regroupV0_lo_6[3673:3672], regroupV0_lo_6[3665:3664]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_4 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo = {regroupV0_lo_6[3689:3688], regroupV0_lo_6[3681:3680]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi = {regroupV0_lo_6[3705:3704], regroupV0_lo_6[3697:3696]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_4 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi, regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_lo_hi_6 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_4, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_4};
  wire [31:0]        regroupV0_lo_hi_hi_hi_lo_lo_6 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_6, regroupV0_lo_hi_hi_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo = {regroupV0_lo_6[3721:3720], regroupV0_lo_6[3713:3712]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi = {regroupV0_lo_6[3737:3736], regroupV0_lo_6[3729:3728]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_4 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo = {regroupV0_lo_6[3753:3752], regroupV0_lo_6[3745:3744]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi = {regroupV0_lo_6[3769:3768], regroupV0_lo_6[3761:3760]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_4 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi, regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_hi_lo_6 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_4, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_4};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo = {regroupV0_lo_6[3785:3784], regroupV0_lo_6[3777:3776]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi = {regroupV0_lo_6[3801:3800], regroupV0_lo_6[3793:3792]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_4 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo = {regroupV0_lo_6[3817:3816], regroupV0_lo_6[3809:3808]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi = {regroupV0_lo_6[3833:3832], regroupV0_lo_6[3825:3824]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_4 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi, regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_hi_hi_6 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_4, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_4};
  wire [31:0]        regroupV0_lo_hi_hi_hi_lo_hi_6 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_6, regroupV0_lo_hi_hi_hi_lo_hi_lo_6};
  wire [63:0]        regroupV0_lo_hi_hi_hi_lo_6 = {regroupV0_lo_hi_hi_hi_lo_hi_6, regroupV0_lo_hi_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo = {regroupV0_lo_6[3849:3848], regroupV0_lo_6[3841:3840]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi = {regroupV0_lo_6[3865:3864], regroupV0_lo_6[3857:3856]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_4 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo = {regroupV0_lo_6[3881:3880], regroupV0_lo_6[3873:3872]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi = {regroupV0_lo_6[3897:3896], regroupV0_lo_6[3889:3888]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_4 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi, regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_lo_lo_6 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_4, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_4};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo = {regroupV0_lo_6[3913:3912], regroupV0_lo_6[3905:3904]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi = {regroupV0_lo_6[3929:3928], regroupV0_lo_6[3921:3920]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_4 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo = {regroupV0_lo_6[3945:3944], regroupV0_lo_6[3937:3936]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi = {regroupV0_lo_6[3961:3960], regroupV0_lo_6[3953:3952]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_4 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi, regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_lo_hi_6 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_4, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_4};
  wire [31:0]        regroupV0_lo_hi_hi_hi_hi_lo_6 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_6, regroupV0_lo_hi_hi_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo = {regroupV0_lo_6[3977:3976], regroupV0_lo_6[3969:3968]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi = {regroupV0_lo_6[3993:3992], regroupV0_lo_6[3985:3984]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_4 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo = {regroupV0_lo_6[4009:4008], regroupV0_lo_6[4001:4000]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi = {regroupV0_lo_6[4025:4024], regroupV0_lo_6[4017:4016]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_4 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi, regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_hi_lo_6 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_4, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_4};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo = {regroupV0_lo_6[4041:4040], regroupV0_lo_6[4033:4032]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi = {regroupV0_lo_6[4057:4056], regroupV0_lo_6[4049:4048]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_4 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo = {regroupV0_lo_6[4073:4072], regroupV0_lo_6[4065:4064]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi = {regroupV0_lo_6[4089:4088], regroupV0_lo_6[4081:4080]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_4 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi, regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_hi_hi_6 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_4, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_4};
  wire [31:0]        regroupV0_lo_hi_hi_hi_hi_hi_6 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_6, regroupV0_lo_hi_hi_hi_hi_hi_lo_6};
  wire [63:0]        regroupV0_lo_hi_hi_hi_hi_6 = {regroupV0_lo_hi_hi_hi_hi_hi_6, regroupV0_lo_hi_hi_hi_hi_lo_6};
  wire [127:0]       regroupV0_lo_hi_hi_hi_6 = {regroupV0_lo_hi_hi_hi_hi_6, regroupV0_lo_hi_hi_hi_lo_6};
  wire [255:0]       regroupV0_lo_hi_hi_6 = {regroupV0_lo_hi_hi_hi_6, regroupV0_lo_hi_hi_lo_6};
  wire [511:0]       regroupV0_lo_hi_6 = {regroupV0_lo_hi_hi_6, regroupV0_lo_hi_lo_6};
  wire [1023:0]      regroupV0_lo_7 = {regroupV0_lo_hi_6, regroupV0_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo = {regroupV0_hi_6[9:8], regroupV0_hi_6[1:0]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi = {regroupV0_hi_6[25:24], regroupV0_hi_6[17:16]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_4 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo = {regroupV0_hi_6[41:40], regroupV0_hi_6[33:32]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi = {regroupV0_hi_6[57:56], regroupV0_hi_6[49:48]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_4 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi, regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_lo_lo_6 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_4, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_4};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo = {regroupV0_hi_6[73:72], regroupV0_hi_6[65:64]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi = {regroupV0_hi_6[89:88], regroupV0_hi_6[81:80]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_4 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo = {regroupV0_hi_6[105:104], regroupV0_hi_6[97:96]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi = {regroupV0_hi_6[121:120], regroupV0_hi_6[113:112]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_4 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi, regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_lo_hi_6 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_4, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_4};
  wire [31:0]        regroupV0_hi_lo_lo_lo_lo_lo_6 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_6, regroupV0_hi_lo_lo_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo = {regroupV0_hi_6[137:136], regroupV0_hi_6[129:128]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi = {regroupV0_hi_6[153:152], regroupV0_hi_6[145:144]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_4 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo = {regroupV0_hi_6[169:168], regroupV0_hi_6[161:160]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi = {regroupV0_hi_6[185:184], regroupV0_hi_6[177:176]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_4 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi, regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_hi_lo_6 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_4, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_4};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo = {regroupV0_hi_6[201:200], regroupV0_hi_6[193:192]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi = {regroupV0_hi_6[217:216], regroupV0_hi_6[209:208]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_4 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo = {regroupV0_hi_6[233:232], regroupV0_hi_6[225:224]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi = {regroupV0_hi_6[249:248], regroupV0_hi_6[241:240]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_4 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi, regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_hi_hi_6 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_4, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_4};
  wire [31:0]        regroupV0_hi_lo_lo_lo_lo_hi_6 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_6, regroupV0_hi_lo_lo_lo_lo_hi_lo_6};
  wire [63:0]        regroupV0_hi_lo_lo_lo_lo_6 = {regroupV0_hi_lo_lo_lo_lo_hi_6, regroupV0_hi_lo_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo = {regroupV0_hi_6[265:264], regroupV0_hi_6[257:256]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi = {regroupV0_hi_6[281:280], regroupV0_hi_6[273:272]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_4 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo = {regroupV0_hi_6[297:296], regroupV0_hi_6[289:288]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi = {regroupV0_hi_6[313:312], regroupV0_hi_6[305:304]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_4 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi, regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_lo_lo_6 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_4, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_4};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo = {regroupV0_hi_6[329:328], regroupV0_hi_6[321:320]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi = {regroupV0_hi_6[345:344], regroupV0_hi_6[337:336]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_4 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo = {regroupV0_hi_6[361:360], regroupV0_hi_6[353:352]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi = {regroupV0_hi_6[377:376], regroupV0_hi_6[369:368]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_4 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi, regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_lo_hi_6 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_4, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_4};
  wire [31:0]        regroupV0_hi_lo_lo_lo_hi_lo_6 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_6, regroupV0_hi_lo_lo_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo = {regroupV0_hi_6[393:392], regroupV0_hi_6[385:384]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi = {regroupV0_hi_6[409:408], regroupV0_hi_6[401:400]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_4 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo = {regroupV0_hi_6[425:424], regroupV0_hi_6[417:416]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi = {regroupV0_hi_6[441:440], regroupV0_hi_6[433:432]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_4 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi, regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_hi_lo_6 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_4, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_4};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo = {regroupV0_hi_6[457:456], regroupV0_hi_6[449:448]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi = {regroupV0_hi_6[473:472], regroupV0_hi_6[465:464]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_4 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo = {regroupV0_hi_6[489:488], regroupV0_hi_6[481:480]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi = {regroupV0_hi_6[505:504], regroupV0_hi_6[497:496]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_4 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi, regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_hi_hi_6 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_4, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_4};
  wire [31:0]        regroupV0_hi_lo_lo_lo_hi_hi_6 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_6, regroupV0_hi_lo_lo_lo_hi_hi_lo_6};
  wire [63:0]        regroupV0_hi_lo_lo_lo_hi_6 = {regroupV0_hi_lo_lo_lo_hi_hi_6, regroupV0_hi_lo_lo_lo_hi_lo_6};
  wire [127:0]       regroupV0_hi_lo_lo_lo_6 = {regroupV0_hi_lo_lo_lo_hi_6, regroupV0_hi_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo = {regroupV0_hi_6[521:520], regroupV0_hi_6[513:512]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi = {regroupV0_hi_6[537:536], regroupV0_hi_6[529:528]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_4 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo = {regroupV0_hi_6[553:552], regroupV0_hi_6[545:544]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi = {regroupV0_hi_6[569:568], regroupV0_hi_6[561:560]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_4 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi, regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_lo_lo_6 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_4, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_4};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo = {regroupV0_hi_6[585:584], regroupV0_hi_6[577:576]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi = {regroupV0_hi_6[601:600], regroupV0_hi_6[593:592]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_4 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo = {regroupV0_hi_6[617:616], regroupV0_hi_6[609:608]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi = {regroupV0_hi_6[633:632], regroupV0_hi_6[625:624]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_4 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi, regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_lo_hi_6 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_4, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_4};
  wire [31:0]        regroupV0_hi_lo_lo_hi_lo_lo_6 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_6, regroupV0_hi_lo_lo_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo = {regroupV0_hi_6[649:648], regroupV0_hi_6[641:640]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi = {regroupV0_hi_6[665:664], regroupV0_hi_6[657:656]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_4 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo = {regroupV0_hi_6[681:680], regroupV0_hi_6[673:672]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi = {regroupV0_hi_6[697:696], regroupV0_hi_6[689:688]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_4 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi, regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_hi_lo_6 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_4, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_4};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo = {regroupV0_hi_6[713:712], regroupV0_hi_6[705:704]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi = {regroupV0_hi_6[729:728], regroupV0_hi_6[721:720]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_4 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo = {regroupV0_hi_6[745:744], regroupV0_hi_6[737:736]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi = {regroupV0_hi_6[761:760], regroupV0_hi_6[753:752]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_4 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi, regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_hi_hi_6 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_4, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_4};
  wire [31:0]        regroupV0_hi_lo_lo_hi_lo_hi_6 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_6, regroupV0_hi_lo_lo_hi_lo_hi_lo_6};
  wire [63:0]        regroupV0_hi_lo_lo_hi_lo_6 = {regroupV0_hi_lo_lo_hi_lo_hi_6, regroupV0_hi_lo_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo = {regroupV0_hi_6[777:776], regroupV0_hi_6[769:768]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi = {regroupV0_hi_6[793:792], regroupV0_hi_6[785:784]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_4 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo = {regroupV0_hi_6[809:808], regroupV0_hi_6[801:800]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi = {regroupV0_hi_6[825:824], regroupV0_hi_6[817:816]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_4 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi, regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_lo_lo_6 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_4, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_4};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo = {regroupV0_hi_6[841:840], regroupV0_hi_6[833:832]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi = {regroupV0_hi_6[857:856], regroupV0_hi_6[849:848]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_4 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo = {regroupV0_hi_6[873:872], regroupV0_hi_6[865:864]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi = {regroupV0_hi_6[889:888], regroupV0_hi_6[881:880]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_4 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi, regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_lo_hi_6 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_4, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_4};
  wire [31:0]        regroupV0_hi_lo_lo_hi_hi_lo_6 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_6, regroupV0_hi_lo_lo_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo = {regroupV0_hi_6[905:904], regroupV0_hi_6[897:896]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi = {regroupV0_hi_6[921:920], regroupV0_hi_6[913:912]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_4 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo = {regroupV0_hi_6[937:936], regroupV0_hi_6[929:928]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi = {regroupV0_hi_6[953:952], regroupV0_hi_6[945:944]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_4 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi, regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_hi_lo_6 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_4, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_4};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo = {regroupV0_hi_6[969:968], regroupV0_hi_6[961:960]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi = {regroupV0_hi_6[985:984], regroupV0_hi_6[977:976]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_4 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo = {regroupV0_hi_6[1001:1000], regroupV0_hi_6[993:992]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi = {regroupV0_hi_6[1017:1016], regroupV0_hi_6[1009:1008]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_4 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi, regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_hi_hi_6 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_4, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_4};
  wire [31:0]        regroupV0_hi_lo_lo_hi_hi_hi_6 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_6, regroupV0_hi_lo_lo_hi_hi_hi_lo_6};
  wire [63:0]        regroupV0_hi_lo_lo_hi_hi_6 = {regroupV0_hi_lo_lo_hi_hi_hi_6, regroupV0_hi_lo_lo_hi_hi_lo_6};
  wire [127:0]       regroupV0_hi_lo_lo_hi_6 = {regroupV0_hi_lo_lo_hi_hi_6, regroupV0_hi_lo_lo_hi_lo_6};
  wire [255:0]       regroupV0_hi_lo_lo_6 = {regroupV0_hi_lo_lo_hi_6, regroupV0_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo = {regroupV0_hi_6[1033:1032], regroupV0_hi_6[1025:1024]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi = {regroupV0_hi_6[1049:1048], regroupV0_hi_6[1041:1040]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_4 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo = {regroupV0_hi_6[1065:1064], regroupV0_hi_6[1057:1056]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi = {regroupV0_hi_6[1081:1080], regroupV0_hi_6[1073:1072]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_4 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi, regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_lo_lo_6 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_4, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_4};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo = {regroupV0_hi_6[1097:1096], regroupV0_hi_6[1089:1088]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi = {regroupV0_hi_6[1113:1112], regroupV0_hi_6[1105:1104]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_4 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo = {regroupV0_hi_6[1129:1128], regroupV0_hi_6[1121:1120]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi = {regroupV0_hi_6[1145:1144], regroupV0_hi_6[1137:1136]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_4 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi, regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_lo_hi_6 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_4, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_4};
  wire [31:0]        regroupV0_hi_lo_hi_lo_lo_lo_6 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_6, regroupV0_hi_lo_hi_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo = {regroupV0_hi_6[1161:1160], regroupV0_hi_6[1153:1152]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi = {regroupV0_hi_6[1177:1176], regroupV0_hi_6[1169:1168]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_4 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo = {regroupV0_hi_6[1193:1192], regroupV0_hi_6[1185:1184]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi = {regroupV0_hi_6[1209:1208], regroupV0_hi_6[1201:1200]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_4 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi, regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_hi_lo_6 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_4, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_4};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo = {regroupV0_hi_6[1225:1224], regroupV0_hi_6[1217:1216]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi = {regroupV0_hi_6[1241:1240], regroupV0_hi_6[1233:1232]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_4 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo = {regroupV0_hi_6[1257:1256], regroupV0_hi_6[1249:1248]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi = {regroupV0_hi_6[1273:1272], regroupV0_hi_6[1265:1264]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_4 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi, regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_hi_hi_6 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_4, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_4};
  wire [31:0]        regroupV0_hi_lo_hi_lo_lo_hi_6 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_6, regroupV0_hi_lo_hi_lo_lo_hi_lo_6};
  wire [63:0]        regroupV0_hi_lo_hi_lo_lo_6 = {regroupV0_hi_lo_hi_lo_lo_hi_6, regroupV0_hi_lo_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo = {regroupV0_hi_6[1289:1288], regroupV0_hi_6[1281:1280]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi = {regroupV0_hi_6[1305:1304], regroupV0_hi_6[1297:1296]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_4 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo = {regroupV0_hi_6[1321:1320], regroupV0_hi_6[1313:1312]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi = {regroupV0_hi_6[1337:1336], regroupV0_hi_6[1329:1328]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_4 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi, regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_lo_lo_6 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_4, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_4};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo = {regroupV0_hi_6[1353:1352], regroupV0_hi_6[1345:1344]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi = {regroupV0_hi_6[1369:1368], regroupV0_hi_6[1361:1360]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_4 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo = {regroupV0_hi_6[1385:1384], regroupV0_hi_6[1377:1376]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi = {regroupV0_hi_6[1401:1400], regroupV0_hi_6[1393:1392]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_4 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi, regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_lo_hi_6 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_4, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_4};
  wire [31:0]        regroupV0_hi_lo_hi_lo_hi_lo_6 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_6, regroupV0_hi_lo_hi_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo = {regroupV0_hi_6[1417:1416], regroupV0_hi_6[1409:1408]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi = {regroupV0_hi_6[1433:1432], regroupV0_hi_6[1425:1424]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_4 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo = {regroupV0_hi_6[1449:1448], regroupV0_hi_6[1441:1440]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi = {regroupV0_hi_6[1465:1464], regroupV0_hi_6[1457:1456]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_4 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi, regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_hi_lo_6 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_4, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_4};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo = {regroupV0_hi_6[1481:1480], regroupV0_hi_6[1473:1472]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi = {regroupV0_hi_6[1497:1496], regroupV0_hi_6[1489:1488]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_4 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo = {regroupV0_hi_6[1513:1512], regroupV0_hi_6[1505:1504]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi = {regroupV0_hi_6[1529:1528], regroupV0_hi_6[1521:1520]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_4 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi, regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_hi_hi_6 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_4, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_4};
  wire [31:0]        regroupV0_hi_lo_hi_lo_hi_hi_6 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_6, regroupV0_hi_lo_hi_lo_hi_hi_lo_6};
  wire [63:0]        regroupV0_hi_lo_hi_lo_hi_6 = {regroupV0_hi_lo_hi_lo_hi_hi_6, regroupV0_hi_lo_hi_lo_hi_lo_6};
  wire [127:0]       regroupV0_hi_lo_hi_lo_6 = {regroupV0_hi_lo_hi_lo_hi_6, regroupV0_hi_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo = {regroupV0_hi_6[1545:1544], regroupV0_hi_6[1537:1536]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi = {regroupV0_hi_6[1561:1560], regroupV0_hi_6[1553:1552]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_4 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo = {regroupV0_hi_6[1577:1576], regroupV0_hi_6[1569:1568]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi = {regroupV0_hi_6[1593:1592], regroupV0_hi_6[1585:1584]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_4 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi, regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_lo_lo_6 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_4, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_4};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo = {regroupV0_hi_6[1609:1608], regroupV0_hi_6[1601:1600]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi = {regroupV0_hi_6[1625:1624], regroupV0_hi_6[1617:1616]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_4 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo = {regroupV0_hi_6[1641:1640], regroupV0_hi_6[1633:1632]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi = {regroupV0_hi_6[1657:1656], regroupV0_hi_6[1649:1648]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_4 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi, regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_lo_hi_6 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_4, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_4};
  wire [31:0]        regroupV0_hi_lo_hi_hi_lo_lo_6 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_6, regroupV0_hi_lo_hi_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo = {regroupV0_hi_6[1673:1672], regroupV0_hi_6[1665:1664]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi = {regroupV0_hi_6[1689:1688], regroupV0_hi_6[1681:1680]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_4 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo = {regroupV0_hi_6[1705:1704], regroupV0_hi_6[1697:1696]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi = {regroupV0_hi_6[1721:1720], regroupV0_hi_6[1713:1712]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_4 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi, regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_hi_lo_6 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_4, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_4};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo = {regroupV0_hi_6[1737:1736], regroupV0_hi_6[1729:1728]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi = {regroupV0_hi_6[1753:1752], regroupV0_hi_6[1745:1744]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_4 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo = {regroupV0_hi_6[1769:1768], regroupV0_hi_6[1761:1760]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi = {regroupV0_hi_6[1785:1784], regroupV0_hi_6[1777:1776]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_4 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi, regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_hi_hi_6 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_4, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_4};
  wire [31:0]        regroupV0_hi_lo_hi_hi_lo_hi_6 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_6, regroupV0_hi_lo_hi_hi_lo_hi_lo_6};
  wire [63:0]        regroupV0_hi_lo_hi_hi_lo_6 = {regroupV0_hi_lo_hi_hi_lo_hi_6, regroupV0_hi_lo_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo = {regroupV0_hi_6[1801:1800], regroupV0_hi_6[1793:1792]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi = {regroupV0_hi_6[1817:1816], regroupV0_hi_6[1809:1808]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_4 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo = {regroupV0_hi_6[1833:1832], regroupV0_hi_6[1825:1824]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi = {regroupV0_hi_6[1849:1848], regroupV0_hi_6[1841:1840]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_4 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi, regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_lo_lo_6 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_4, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_4};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo = {regroupV0_hi_6[1865:1864], regroupV0_hi_6[1857:1856]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi = {regroupV0_hi_6[1881:1880], regroupV0_hi_6[1873:1872]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_4 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo = {regroupV0_hi_6[1897:1896], regroupV0_hi_6[1889:1888]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi = {regroupV0_hi_6[1913:1912], regroupV0_hi_6[1905:1904]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_4 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi, regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_lo_hi_6 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_4, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_4};
  wire [31:0]        regroupV0_hi_lo_hi_hi_hi_lo_6 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_6, regroupV0_hi_lo_hi_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo = {regroupV0_hi_6[1929:1928], regroupV0_hi_6[1921:1920]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi = {regroupV0_hi_6[1945:1944], regroupV0_hi_6[1937:1936]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_4 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo = {regroupV0_hi_6[1961:1960], regroupV0_hi_6[1953:1952]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi = {regroupV0_hi_6[1977:1976], regroupV0_hi_6[1969:1968]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_4 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi, regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_hi_lo_6 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_4, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_4};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo = {regroupV0_hi_6[1993:1992], regroupV0_hi_6[1985:1984]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi = {regroupV0_hi_6[2009:2008], regroupV0_hi_6[2001:2000]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_4 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo = {regroupV0_hi_6[2025:2024], regroupV0_hi_6[2017:2016]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi = {regroupV0_hi_6[2041:2040], regroupV0_hi_6[2033:2032]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_4 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi, regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_hi_hi_6 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_4, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_4};
  wire [31:0]        regroupV0_hi_lo_hi_hi_hi_hi_6 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_6, regroupV0_hi_lo_hi_hi_hi_hi_lo_6};
  wire [63:0]        regroupV0_hi_lo_hi_hi_hi_6 = {regroupV0_hi_lo_hi_hi_hi_hi_6, regroupV0_hi_lo_hi_hi_hi_lo_6};
  wire [127:0]       regroupV0_hi_lo_hi_hi_6 = {regroupV0_hi_lo_hi_hi_hi_6, regroupV0_hi_lo_hi_hi_lo_6};
  wire [255:0]       regroupV0_hi_lo_hi_6 = {regroupV0_hi_lo_hi_hi_6, regroupV0_hi_lo_hi_lo_6};
  wire [511:0]       regroupV0_hi_lo_6 = {regroupV0_hi_lo_hi_6, regroupV0_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo = {regroupV0_hi_6[2057:2056], regroupV0_hi_6[2049:2048]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi = {regroupV0_hi_6[2073:2072], regroupV0_hi_6[2065:2064]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_4 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo = {regroupV0_hi_6[2089:2088], regroupV0_hi_6[2081:2080]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi = {regroupV0_hi_6[2105:2104], regroupV0_hi_6[2097:2096]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_4 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi, regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_lo_lo_6 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_4, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_4};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo = {regroupV0_hi_6[2121:2120], regroupV0_hi_6[2113:2112]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi = {regroupV0_hi_6[2137:2136], regroupV0_hi_6[2129:2128]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_4 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo = {regroupV0_hi_6[2153:2152], regroupV0_hi_6[2145:2144]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi = {regroupV0_hi_6[2169:2168], regroupV0_hi_6[2161:2160]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_4 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi, regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_lo_hi_6 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_4, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_4};
  wire [31:0]        regroupV0_hi_hi_lo_lo_lo_lo_6 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_6, regroupV0_hi_hi_lo_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo = {regroupV0_hi_6[2185:2184], regroupV0_hi_6[2177:2176]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi = {regroupV0_hi_6[2201:2200], regroupV0_hi_6[2193:2192]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_4 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo = {regroupV0_hi_6[2217:2216], regroupV0_hi_6[2209:2208]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi = {regroupV0_hi_6[2233:2232], regroupV0_hi_6[2225:2224]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_4 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi, regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_hi_lo_6 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_4, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_4};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo = {regroupV0_hi_6[2249:2248], regroupV0_hi_6[2241:2240]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi = {regroupV0_hi_6[2265:2264], regroupV0_hi_6[2257:2256]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_4 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo = {regroupV0_hi_6[2281:2280], regroupV0_hi_6[2273:2272]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi = {regroupV0_hi_6[2297:2296], regroupV0_hi_6[2289:2288]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_4 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi, regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_hi_hi_6 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_4, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_4};
  wire [31:0]        regroupV0_hi_hi_lo_lo_lo_hi_6 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_6, regroupV0_hi_hi_lo_lo_lo_hi_lo_6};
  wire [63:0]        regroupV0_hi_hi_lo_lo_lo_6 = {regroupV0_hi_hi_lo_lo_lo_hi_6, regroupV0_hi_hi_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo = {regroupV0_hi_6[2313:2312], regroupV0_hi_6[2305:2304]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi = {regroupV0_hi_6[2329:2328], regroupV0_hi_6[2321:2320]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_4 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo = {regroupV0_hi_6[2345:2344], regroupV0_hi_6[2337:2336]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi = {regroupV0_hi_6[2361:2360], regroupV0_hi_6[2353:2352]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_4 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi, regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_lo_lo_6 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_4, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_4};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo = {regroupV0_hi_6[2377:2376], regroupV0_hi_6[2369:2368]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi = {regroupV0_hi_6[2393:2392], regroupV0_hi_6[2385:2384]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_4 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo = {regroupV0_hi_6[2409:2408], regroupV0_hi_6[2401:2400]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi = {regroupV0_hi_6[2425:2424], regroupV0_hi_6[2417:2416]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_4 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi, regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_lo_hi_6 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_4, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_4};
  wire [31:0]        regroupV0_hi_hi_lo_lo_hi_lo_6 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_6, regroupV0_hi_hi_lo_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo = {regroupV0_hi_6[2441:2440], regroupV0_hi_6[2433:2432]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi = {regroupV0_hi_6[2457:2456], regroupV0_hi_6[2449:2448]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_4 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo = {regroupV0_hi_6[2473:2472], regroupV0_hi_6[2465:2464]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi = {regroupV0_hi_6[2489:2488], regroupV0_hi_6[2481:2480]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_4 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi, regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_hi_lo_6 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_4, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_4};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo = {regroupV0_hi_6[2505:2504], regroupV0_hi_6[2497:2496]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi = {regroupV0_hi_6[2521:2520], regroupV0_hi_6[2513:2512]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_4 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo = {regroupV0_hi_6[2537:2536], regroupV0_hi_6[2529:2528]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi = {regroupV0_hi_6[2553:2552], regroupV0_hi_6[2545:2544]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_4 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi, regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_hi_hi_6 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_4, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_4};
  wire [31:0]        regroupV0_hi_hi_lo_lo_hi_hi_6 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_6, regroupV0_hi_hi_lo_lo_hi_hi_lo_6};
  wire [63:0]        regroupV0_hi_hi_lo_lo_hi_6 = {regroupV0_hi_hi_lo_lo_hi_hi_6, regroupV0_hi_hi_lo_lo_hi_lo_6};
  wire [127:0]       regroupV0_hi_hi_lo_lo_6 = {regroupV0_hi_hi_lo_lo_hi_6, regroupV0_hi_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo = {regroupV0_hi_6[2569:2568], regroupV0_hi_6[2561:2560]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi = {regroupV0_hi_6[2585:2584], regroupV0_hi_6[2577:2576]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_4 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo = {regroupV0_hi_6[2601:2600], regroupV0_hi_6[2593:2592]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi = {regroupV0_hi_6[2617:2616], regroupV0_hi_6[2609:2608]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_4 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi, regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_lo_lo_6 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_4, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_4};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo = {regroupV0_hi_6[2633:2632], regroupV0_hi_6[2625:2624]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi = {regroupV0_hi_6[2649:2648], regroupV0_hi_6[2641:2640]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_4 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo = {regroupV0_hi_6[2665:2664], regroupV0_hi_6[2657:2656]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi = {regroupV0_hi_6[2681:2680], regroupV0_hi_6[2673:2672]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_4 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi, regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_lo_hi_6 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_4, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_4};
  wire [31:0]        regroupV0_hi_hi_lo_hi_lo_lo_6 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_6, regroupV0_hi_hi_lo_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo = {regroupV0_hi_6[2697:2696], regroupV0_hi_6[2689:2688]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi = {regroupV0_hi_6[2713:2712], regroupV0_hi_6[2705:2704]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_4 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo = {regroupV0_hi_6[2729:2728], regroupV0_hi_6[2721:2720]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi = {regroupV0_hi_6[2745:2744], regroupV0_hi_6[2737:2736]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_4 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi, regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_hi_lo_6 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_4, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_4};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo = {regroupV0_hi_6[2761:2760], regroupV0_hi_6[2753:2752]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi = {regroupV0_hi_6[2777:2776], regroupV0_hi_6[2769:2768]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_4 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo = {regroupV0_hi_6[2793:2792], regroupV0_hi_6[2785:2784]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi = {regroupV0_hi_6[2809:2808], regroupV0_hi_6[2801:2800]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_4 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi, regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_hi_hi_6 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_4, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_4};
  wire [31:0]        regroupV0_hi_hi_lo_hi_lo_hi_6 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_6, regroupV0_hi_hi_lo_hi_lo_hi_lo_6};
  wire [63:0]        regroupV0_hi_hi_lo_hi_lo_6 = {regroupV0_hi_hi_lo_hi_lo_hi_6, regroupV0_hi_hi_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo = {regroupV0_hi_6[2825:2824], regroupV0_hi_6[2817:2816]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi = {regroupV0_hi_6[2841:2840], regroupV0_hi_6[2833:2832]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_4 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo = {regroupV0_hi_6[2857:2856], regroupV0_hi_6[2849:2848]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi = {regroupV0_hi_6[2873:2872], regroupV0_hi_6[2865:2864]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_4 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi, regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_lo_lo_6 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_4, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_4};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo = {regroupV0_hi_6[2889:2888], regroupV0_hi_6[2881:2880]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi = {regroupV0_hi_6[2905:2904], regroupV0_hi_6[2897:2896]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_4 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo = {regroupV0_hi_6[2921:2920], regroupV0_hi_6[2913:2912]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi = {regroupV0_hi_6[2937:2936], regroupV0_hi_6[2929:2928]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_4 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi, regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_lo_hi_6 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_4, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_4};
  wire [31:0]        regroupV0_hi_hi_lo_hi_hi_lo_6 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_6, regroupV0_hi_hi_lo_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo = {regroupV0_hi_6[2953:2952], regroupV0_hi_6[2945:2944]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi = {regroupV0_hi_6[2969:2968], regroupV0_hi_6[2961:2960]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_4 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo = {regroupV0_hi_6[2985:2984], regroupV0_hi_6[2977:2976]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi = {regroupV0_hi_6[3001:3000], regroupV0_hi_6[2993:2992]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_4 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi, regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_hi_lo_6 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_4, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_4};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo = {regroupV0_hi_6[3017:3016], regroupV0_hi_6[3009:3008]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi = {regroupV0_hi_6[3033:3032], regroupV0_hi_6[3025:3024]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_4 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo = {regroupV0_hi_6[3049:3048], regroupV0_hi_6[3041:3040]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi = {regroupV0_hi_6[3065:3064], regroupV0_hi_6[3057:3056]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_4 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi, regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_hi_hi_6 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_4, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_4};
  wire [31:0]        regroupV0_hi_hi_lo_hi_hi_hi_6 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_6, regroupV0_hi_hi_lo_hi_hi_hi_lo_6};
  wire [63:0]        regroupV0_hi_hi_lo_hi_hi_6 = {regroupV0_hi_hi_lo_hi_hi_hi_6, regroupV0_hi_hi_lo_hi_hi_lo_6};
  wire [127:0]       regroupV0_hi_hi_lo_hi_6 = {regroupV0_hi_hi_lo_hi_hi_6, regroupV0_hi_hi_lo_hi_lo_6};
  wire [255:0]       regroupV0_hi_hi_lo_6 = {regroupV0_hi_hi_lo_hi_6, regroupV0_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo = {regroupV0_hi_6[3081:3080], regroupV0_hi_6[3073:3072]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi = {regroupV0_hi_6[3097:3096], regroupV0_hi_6[3089:3088]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_4 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo = {regroupV0_hi_6[3113:3112], regroupV0_hi_6[3105:3104]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi = {regroupV0_hi_6[3129:3128], regroupV0_hi_6[3121:3120]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_4 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi, regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_lo_lo_6 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_4, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_4};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo = {regroupV0_hi_6[3145:3144], regroupV0_hi_6[3137:3136]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi = {regroupV0_hi_6[3161:3160], regroupV0_hi_6[3153:3152]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_4 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo = {regroupV0_hi_6[3177:3176], regroupV0_hi_6[3169:3168]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi = {regroupV0_hi_6[3193:3192], regroupV0_hi_6[3185:3184]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_4 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi, regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_lo_hi_6 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_4, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_4};
  wire [31:0]        regroupV0_hi_hi_hi_lo_lo_lo_6 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_6, regroupV0_hi_hi_hi_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo = {regroupV0_hi_6[3209:3208], regroupV0_hi_6[3201:3200]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi = {regroupV0_hi_6[3225:3224], regroupV0_hi_6[3217:3216]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_4 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo = {regroupV0_hi_6[3241:3240], regroupV0_hi_6[3233:3232]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi = {regroupV0_hi_6[3257:3256], regroupV0_hi_6[3249:3248]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_4 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi, regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_hi_lo_6 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_4, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_4};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo = {regroupV0_hi_6[3273:3272], regroupV0_hi_6[3265:3264]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi = {regroupV0_hi_6[3289:3288], regroupV0_hi_6[3281:3280]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_4 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo = {regroupV0_hi_6[3305:3304], regroupV0_hi_6[3297:3296]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi = {regroupV0_hi_6[3321:3320], regroupV0_hi_6[3313:3312]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_4 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi, regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_hi_hi_6 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_4, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_4};
  wire [31:0]        regroupV0_hi_hi_hi_lo_lo_hi_6 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_6, regroupV0_hi_hi_hi_lo_lo_hi_lo_6};
  wire [63:0]        regroupV0_hi_hi_hi_lo_lo_6 = {regroupV0_hi_hi_hi_lo_lo_hi_6, regroupV0_hi_hi_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo = {regroupV0_hi_6[3337:3336], regroupV0_hi_6[3329:3328]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi = {regroupV0_hi_6[3353:3352], regroupV0_hi_6[3345:3344]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_4 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo = {regroupV0_hi_6[3369:3368], regroupV0_hi_6[3361:3360]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi = {regroupV0_hi_6[3385:3384], regroupV0_hi_6[3377:3376]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_4 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi, regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_lo_lo_6 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_4, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_4};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo = {regroupV0_hi_6[3401:3400], regroupV0_hi_6[3393:3392]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi = {regroupV0_hi_6[3417:3416], regroupV0_hi_6[3409:3408]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_4 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo = {regroupV0_hi_6[3433:3432], regroupV0_hi_6[3425:3424]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi = {regroupV0_hi_6[3449:3448], regroupV0_hi_6[3441:3440]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_4 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi, regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_lo_hi_6 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_4, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_4};
  wire [31:0]        regroupV0_hi_hi_hi_lo_hi_lo_6 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_6, regroupV0_hi_hi_hi_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo = {regroupV0_hi_6[3465:3464], regroupV0_hi_6[3457:3456]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi = {regroupV0_hi_6[3481:3480], regroupV0_hi_6[3473:3472]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_4 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo = {regroupV0_hi_6[3497:3496], regroupV0_hi_6[3489:3488]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi = {regroupV0_hi_6[3513:3512], regroupV0_hi_6[3505:3504]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_4 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi, regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_hi_lo_6 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_4, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_4};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo = {regroupV0_hi_6[3529:3528], regroupV0_hi_6[3521:3520]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi = {regroupV0_hi_6[3545:3544], regroupV0_hi_6[3537:3536]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_4 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo = {regroupV0_hi_6[3561:3560], regroupV0_hi_6[3553:3552]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi = {regroupV0_hi_6[3577:3576], regroupV0_hi_6[3569:3568]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_4 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi, regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_hi_hi_6 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_4, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_4};
  wire [31:0]        regroupV0_hi_hi_hi_lo_hi_hi_6 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_6, regroupV0_hi_hi_hi_lo_hi_hi_lo_6};
  wire [63:0]        regroupV0_hi_hi_hi_lo_hi_6 = {regroupV0_hi_hi_hi_lo_hi_hi_6, regroupV0_hi_hi_hi_lo_hi_lo_6};
  wire [127:0]       regroupV0_hi_hi_hi_lo_6 = {regroupV0_hi_hi_hi_lo_hi_6, regroupV0_hi_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo = {regroupV0_hi_6[3593:3592], regroupV0_hi_6[3585:3584]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi = {regroupV0_hi_6[3609:3608], regroupV0_hi_6[3601:3600]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_4 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo = {regroupV0_hi_6[3625:3624], regroupV0_hi_6[3617:3616]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi = {regroupV0_hi_6[3641:3640], regroupV0_hi_6[3633:3632]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_4 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi, regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_lo_lo_6 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_4, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_4};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo = {regroupV0_hi_6[3657:3656], regroupV0_hi_6[3649:3648]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi = {regroupV0_hi_6[3673:3672], regroupV0_hi_6[3665:3664]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_4 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo = {regroupV0_hi_6[3689:3688], regroupV0_hi_6[3681:3680]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi = {regroupV0_hi_6[3705:3704], regroupV0_hi_6[3697:3696]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_4 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi, regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_lo_hi_6 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_4, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_4};
  wire [31:0]        regroupV0_hi_hi_hi_hi_lo_lo_6 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_6, regroupV0_hi_hi_hi_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo = {regroupV0_hi_6[3721:3720], regroupV0_hi_6[3713:3712]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi = {regroupV0_hi_6[3737:3736], regroupV0_hi_6[3729:3728]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_4 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo = {regroupV0_hi_6[3753:3752], regroupV0_hi_6[3745:3744]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi = {regroupV0_hi_6[3769:3768], regroupV0_hi_6[3761:3760]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_4 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi, regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_hi_lo_6 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_4, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_4};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo = {regroupV0_hi_6[3785:3784], regroupV0_hi_6[3777:3776]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi = {regroupV0_hi_6[3801:3800], regroupV0_hi_6[3793:3792]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_4 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo = {regroupV0_hi_6[3817:3816], regroupV0_hi_6[3809:3808]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi = {regroupV0_hi_6[3833:3832], regroupV0_hi_6[3825:3824]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_4 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi, regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_hi_hi_6 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_4, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_4};
  wire [31:0]        regroupV0_hi_hi_hi_hi_lo_hi_6 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_6, regroupV0_hi_hi_hi_hi_lo_hi_lo_6};
  wire [63:0]        regroupV0_hi_hi_hi_hi_lo_6 = {regroupV0_hi_hi_hi_hi_lo_hi_6, regroupV0_hi_hi_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo = {regroupV0_hi_6[3849:3848], regroupV0_hi_6[3841:3840]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi = {regroupV0_hi_6[3865:3864], regroupV0_hi_6[3857:3856]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_4 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo = {regroupV0_hi_6[3881:3880], regroupV0_hi_6[3873:3872]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi = {regroupV0_hi_6[3897:3896], regroupV0_hi_6[3889:3888]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_4 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi, regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_lo_lo_6 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_4, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_4};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo = {regroupV0_hi_6[3913:3912], regroupV0_hi_6[3905:3904]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi = {regroupV0_hi_6[3929:3928], regroupV0_hi_6[3921:3920]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_4 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo = {regroupV0_hi_6[3945:3944], regroupV0_hi_6[3937:3936]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi = {regroupV0_hi_6[3961:3960], regroupV0_hi_6[3953:3952]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_4 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi, regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_lo_hi_6 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_4, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_4};
  wire [31:0]        regroupV0_hi_hi_hi_hi_hi_lo_6 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_6, regroupV0_hi_hi_hi_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo = {regroupV0_hi_6[3977:3976], regroupV0_hi_6[3969:3968]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi = {regroupV0_hi_6[3993:3992], regroupV0_hi_6[3985:3984]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_4 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo = {regroupV0_hi_6[4009:4008], regroupV0_hi_6[4001:4000]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi = {regroupV0_hi_6[4025:4024], regroupV0_hi_6[4017:4016]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_4 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi, regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_hi_lo_6 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_4, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_4};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo = {regroupV0_hi_6[4041:4040], regroupV0_hi_6[4033:4032]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi = {regroupV0_hi_6[4057:4056], regroupV0_hi_6[4049:4048]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_4 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo = {regroupV0_hi_6[4073:4072], regroupV0_hi_6[4065:4064]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi = {regroupV0_hi_6[4089:4088], regroupV0_hi_6[4081:4080]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_4 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi, regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_hi_hi_6 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_4, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_4};
  wire [31:0]        regroupV0_hi_hi_hi_hi_hi_hi_6 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_6, regroupV0_hi_hi_hi_hi_hi_hi_lo_6};
  wire [63:0]        regroupV0_hi_hi_hi_hi_hi_6 = {regroupV0_hi_hi_hi_hi_hi_hi_6, regroupV0_hi_hi_hi_hi_hi_lo_6};
  wire [127:0]       regroupV0_hi_hi_hi_hi_6 = {regroupV0_hi_hi_hi_hi_hi_6, regroupV0_hi_hi_hi_hi_lo_6};
  wire [255:0]       regroupV0_hi_hi_hi_6 = {regroupV0_hi_hi_hi_hi_6, regroupV0_hi_hi_hi_lo_6};
  wire [511:0]       regroupV0_hi_hi_6 = {regroupV0_hi_hi_hi_6, regroupV0_hi_hi_lo_6};
  wire [1023:0]      regroupV0_hi_7 = {regroupV0_hi_hi_6, regroupV0_hi_lo_6};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo_1 = {regroupV0_lo_6[11:10], regroupV0_lo_6[3:2]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi_1 = {regroupV0_lo_6[27:26], regroupV0_lo_6[19:18]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_5 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo_1 = {regroupV0_lo_6[43:42], regroupV0_lo_6[35:34]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi_1 = {regroupV0_lo_6[59:58], regroupV0_lo_6[51:50]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_5 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi_1, regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_lo_lo_7 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_5, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_5};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo_1 = {regroupV0_lo_6[75:74], regroupV0_lo_6[67:66]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi_1 = {regroupV0_lo_6[91:90], regroupV0_lo_6[83:82]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_5 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi_1, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo_1 = {regroupV0_lo_6[107:106], regroupV0_lo_6[99:98]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi_1 = {regroupV0_lo_6[123:122], regroupV0_lo_6[115:114]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_5 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi_1, regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_lo_hi_7 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_5, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_5};
  wire [31:0]        regroupV0_lo_lo_lo_lo_lo_lo_7 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_7, regroupV0_lo_lo_lo_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo_1 = {regroupV0_lo_6[139:138], regroupV0_lo_6[131:130]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi_1 = {regroupV0_lo_6[155:154], regroupV0_lo_6[147:146]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_5 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo_1 = {regroupV0_lo_6[171:170], regroupV0_lo_6[163:162]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi_1 = {regroupV0_lo_6[187:186], regroupV0_lo_6[179:178]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_5 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi_1, regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_hi_lo_7 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_5, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_5};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo_1 = {regroupV0_lo_6[203:202], regroupV0_lo_6[195:194]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi_1 = {regroupV0_lo_6[219:218], regroupV0_lo_6[211:210]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_5 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi_1, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo_1 = {regroupV0_lo_6[235:234], regroupV0_lo_6[227:226]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi_1 = {regroupV0_lo_6[251:250], regroupV0_lo_6[243:242]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_5 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi_1, regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_hi_hi_7 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_5, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_5};
  wire [31:0]        regroupV0_lo_lo_lo_lo_lo_hi_7 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_7, regroupV0_lo_lo_lo_lo_lo_hi_lo_7};
  wire [63:0]        regroupV0_lo_lo_lo_lo_lo_7 = {regroupV0_lo_lo_lo_lo_lo_hi_7, regroupV0_lo_lo_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo_1 = {regroupV0_lo_6[267:266], regroupV0_lo_6[259:258]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi_1 = {regroupV0_lo_6[283:282], regroupV0_lo_6[275:274]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_5 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo_1 = {regroupV0_lo_6[299:298], regroupV0_lo_6[291:290]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi_1 = {regroupV0_lo_6[315:314], regroupV0_lo_6[307:306]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_5 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi_1, regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_lo_lo_7 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_5, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_5};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo_1 = {regroupV0_lo_6[331:330], regroupV0_lo_6[323:322]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi_1 = {regroupV0_lo_6[347:346], regroupV0_lo_6[339:338]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_5 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi_1, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo_1 = {regroupV0_lo_6[363:362], regroupV0_lo_6[355:354]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi_1 = {regroupV0_lo_6[379:378], regroupV0_lo_6[371:370]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_5 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi_1, regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_lo_hi_7 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_5, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_5};
  wire [31:0]        regroupV0_lo_lo_lo_lo_hi_lo_7 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_7, regroupV0_lo_lo_lo_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo_1 = {regroupV0_lo_6[395:394], regroupV0_lo_6[387:386]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi_1 = {regroupV0_lo_6[411:410], regroupV0_lo_6[403:402]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_5 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo_1 = {regroupV0_lo_6[427:426], regroupV0_lo_6[419:418]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi_1 = {regroupV0_lo_6[443:442], regroupV0_lo_6[435:434]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_5 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi_1, regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_hi_lo_7 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_5, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_5};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo_1 = {regroupV0_lo_6[459:458], regroupV0_lo_6[451:450]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi_1 = {regroupV0_lo_6[475:474], regroupV0_lo_6[467:466]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_5 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi_1, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo_1 = {regroupV0_lo_6[491:490], regroupV0_lo_6[483:482]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi_1 = {regroupV0_lo_6[507:506], regroupV0_lo_6[499:498]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_5 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi_1, regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_hi_hi_7 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_5, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_5};
  wire [31:0]        regroupV0_lo_lo_lo_lo_hi_hi_7 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_7, regroupV0_lo_lo_lo_lo_hi_hi_lo_7};
  wire [63:0]        regroupV0_lo_lo_lo_lo_hi_7 = {regroupV0_lo_lo_lo_lo_hi_hi_7, regroupV0_lo_lo_lo_lo_hi_lo_7};
  wire [127:0]       regroupV0_lo_lo_lo_lo_7 = {regroupV0_lo_lo_lo_lo_hi_7, regroupV0_lo_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo_1 = {regroupV0_lo_6[523:522], regroupV0_lo_6[515:514]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi_1 = {regroupV0_lo_6[539:538], regroupV0_lo_6[531:530]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_5 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo_1 = {regroupV0_lo_6[555:554], regroupV0_lo_6[547:546]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi_1 = {regroupV0_lo_6[571:570], regroupV0_lo_6[563:562]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_5 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi_1, regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_lo_lo_7 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_5, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_5};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo_1 = {regroupV0_lo_6[587:586], regroupV0_lo_6[579:578]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi_1 = {regroupV0_lo_6[603:602], regroupV0_lo_6[595:594]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_5 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi_1, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo_1 = {regroupV0_lo_6[619:618], regroupV0_lo_6[611:610]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi_1 = {regroupV0_lo_6[635:634], regroupV0_lo_6[627:626]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_5 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi_1, regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_lo_hi_7 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_5, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_5};
  wire [31:0]        regroupV0_lo_lo_lo_hi_lo_lo_7 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_7, regroupV0_lo_lo_lo_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo_1 = {regroupV0_lo_6[651:650], regroupV0_lo_6[643:642]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi_1 = {regroupV0_lo_6[667:666], regroupV0_lo_6[659:658]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_5 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi_1, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo_1 = {regroupV0_lo_6[683:682], regroupV0_lo_6[675:674]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi_1 = {regroupV0_lo_6[699:698], regroupV0_lo_6[691:690]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_5 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi_1, regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_hi_lo_7 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_5, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_5};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo_1 = {regroupV0_lo_6[715:714], regroupV0_lo_6[707:706]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi_1 = {regroupV0_lo_6[731:730], regroupV0_lo_6[723:722]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_5 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi_1, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo_1 = {regroupV0_lo_6[747:746], regroupV0_lo_6[739:738]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi_1 = {regroupV0_lo_6[763:762], regroupV0_lo_6[755:754]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_5 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi_1, regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_hi_hi_7 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_5, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_5};
  wire [31:0]        regroupV0_lo_lo_lo_hi_lo_hi_7 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_7, regroupV0_lo_lo_lo_hi_lo_hi_lo_7};
  wire [63:0]        regroupV0_lo_lo_lo_hi_lo_7 = {regroupV0_lo_lo_lo_hi_lo_hi_7, regroupV0_lo_lo_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo_1 = {regroupV0_lo_6[779:778], regroupV0_lo_6[771:770]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi_1 = {regroupV0_lo_6[795:794], regroupV0_lo_6[787:786]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_5 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo_1 = {regroupV0_lo_6[811:810], regroupV0_lo_6[803:802]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi_1 = {regroupV0_lo_6[827:826], regroupV0_lo_6[819:818]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_5 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi_1, regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_lo_lo_7 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_5, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_5};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo_1 = {regroupV0_lo_6[843:842], regroupV0_lo_6[835:834]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi_1 = {regroupV0_lo_6[859:858], regroupV0_lo_6[851:850]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_5 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi_1, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo_1 = {regroupV0_lo_6[875:874], regroupV0_lo_6[867:866]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi_1 = {regroupV0_lo_6[891:890], regroupV0_lo_6[883:882]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_5 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi_1, regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_lo_hi_7 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_5, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_5};
  wire [31:0]        regroupV0_lo_lo_lo_hi_hi_lo_7 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_7, regroupV0_lo_lo_lo_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo_1 = {regroupV0_lo_6[907:906], regroupV0_lo_6[899:898]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi_1 = {regroupV0_lo_6[923:922], regroupV0_lo_6[915:914]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_5 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi_1, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo_1 = {regroupV0_lo_6[939:938], regroupV0_lo_6[931:930]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi_1 = {regroupV0_lo_6[955:954], regroupV0_lo_6[947:946]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_5 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi_1, regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_hi_lo_7 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_5, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_5};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo_1 = {regroupV0_lo_6[971:970], regroupV0_lo_6[963:962]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi_1 = {regroupV0_lo_6[987:986], regroupV0_lo_6[979:978]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_5 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi_1, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo_1 = {regroupV0_lo_6[1003:1002], regroupV0_lo_6[995:994]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi_1 = {regroupV0_lo_6[1019:1018], regroupV0_lo_6[1011:1010]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_5 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi_1, regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_hi_hi_7 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_5, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_5};
  wire [31:0]        regroupV0_lo_lo_lo_hi_hi_hi_7 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_7, regroupV0_lo_lo_lo_hi_hi_hi_lo_7};
  wire [63:0]        regroupV0_lo_lo_lo_hi_hi_7 = {regroupV0_lo_lo_lo_hi_hi_hi_7, regroupV0_lo_lo_lo_hi_hi_lo_7};
  wire [127:0]       regroupV0_lo_lo_lo_hi_7 = {regroupV0_lo_lo_lo_hi_hi_7, regroupV0_lo_lo_lo_hi_lo_7};
  wire [255:0]       regroupV0_lo_lo_lo_7 = {regroupV0_lo_lo_lo_hi_7, regroupV0_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo_1 = {regroupV0_lo_6[1035:1034], regroupV0_lo_6[1027:1026]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi_1 = {regroupV0_lo_6[1051:1050], regroupV0_lo_6[1043:1042]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_5 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi_1, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo_1 = {regroupV0_lo_6[1067:1066], regroupV0_lo_6[1059:1058]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi_1 = {regroupV0_lo_6[1083:1082], regroupV0_lo_6[1075:1074]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_5 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi_1, regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_lo_lo_7 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_5, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_5};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo_1 = {regroupV0_lo_6[1099:1098], regroupV0_lo_6[1091:1090]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi_1 = {regroupV0_lo_6[1115:1114], regroupV0_lo_6[1107:1106]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_5 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi_1, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo_1 = {regroupV0_lo_6[1131:1130], regroupV0_lo_6[1123:1122]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi_1 = {regroupV0_lo_6[1147:1146], regroupV0_lo_6[1139:1138]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_5 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi_1, regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_lo_hi_7 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_5, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_5};
  wire [31:0]        regroupV0_lo_lo_hi_lo_lo_lo_7 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_7, regroupV0_lo_lo_hi_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo_1 = {regroupV0_lo_6[1163:1162], regroupV0_lo_6[1155:1154]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi_1 = {regroupV0_lo_6[1179:1178], regroupV0_lo_6[1171:1170]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_5 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi_1, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo_1 = {regroupV0_lo_6[1195:1194], regroupV0_lo_6[1187:1186]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi_1 = {regroupV0_lo_6[1211:1210], regroupV0_lo_6[1203:1202]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_5 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi_1, regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_hi_lo_7 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_5, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_5};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo_1 = {regroupV0_lo_6[1227:1226], regroupV0_lo_6[1219:1218]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi_1 = {regroupV0_lo_6[1243:1242], regroupV0_lo_6[1235:1234]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_5 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi_1, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo_1 = {regroupV0_lo_6[1259:1258], regroupV0_lo_6[1251:1250]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi_1 = {regroupV0_lo_6[1275:1274], regroupV0_lo_6[1267:1266]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_5 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi_1, regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_hi_hi_7 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_5, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_5};
  wire [31:0]        regroupV0_lo_lo_hi_lo_lo_hi_7 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_7, regroupV0_lo_lo_hi_lo_lo_hi_lo_7};
  wire [63:0]        regroupV0_lo_lo_hi_lo_lo_7 = {regroupV0_lo_lo_hi_lo_lo_hi_7, regroupV0_lo_lo_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo_1 = {regroupV0_lo_6[1291:1290], regroupV0_lo_6[1283:1282]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi_1 = {regroupV0_lo_6[1307:1306], regroupV0_lo_6[1299:1298]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_5 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi_1, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo_1 = {regroupV0_lo_6[1323:1322], regroupV0_lo_6[1315:1314]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi_1 = {regroupV0_lo_6[1339:1338], regroupV0_lo_6[1331:1330]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_5 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi_1, regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_lo_lo_7 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_5, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_5};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo_1 = {regroupV0_lo_6[1355:1354], regroupV0_lo_6[1347:1346]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi_1 = {regroupV0_lo_6[1371:1370], regroupV0_lo_6[1363:1362]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_5 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi_1, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo_1 = {regroupV0_lo_6[1387:1386], regroupV0_lo_6[1379:1378]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi_1 = {regroupV0_lo_6[1403:1402], regroupV0_lo_6[1395:1394]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_5 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi_1, regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_lo_hi_7 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_5, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_5};
  wire [31:0]        regroupV0_lo_lo_hi_lo_hi_lo_7 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_7, regroupV0_lo_lo_hi_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo_1 = {regroupV0_lo_6[1419:1418], regroupV0_lo_6[1411:1410]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi_1 = {regroupV0_lo_6[1435:1434], regroupV0_lo_6[1427:1426]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_5 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi_1, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo_1 = {regroupV0_lo_6[1451:1450], regroupV0_lo_6[1443:1442]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi_1 = {regroupV0_lo_6[1467:1466], regroupV0_lo_6[1459:1458]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_5 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi_1, regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_hi_lo_7 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_5, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_5};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo_1 = {regroupV0_lo_6[1483:1482], regroupV0_lo_6[1475:1474]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi_1 = {regroupV0_lo_6[1499:1498], regroupV0_lo_6[1491:1490]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_5 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi_1, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo_1 = {regroupV0_lo_6[1515:1514], regroupV0_lo_6[1507:1506]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi_1 = {regroupV0_lo_6[1531:1530], regroupV0_lo_6[1523:1522]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_5 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi_1, regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_hi_hi_7 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_5, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_5};
  wire [31:0]        regroupV0_lo_lo_hi_lo_hi_hi_7 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_7, regroupV0_lo_lo_hi_lo_hi_hi_lo_7};
  wire [63:0]        regroupV0_lo_lo_hi_lo_hi_7 = {regroupV0_lo_lo_hi_lo_hi_hi_7, regroupV0_lo_lo_hi_lo_hi_lo_7};
  wire [127:0]       regroupV0_lo_lo_hi_lo_7 = {regroupV0_lo_lo_hi_lo_hi_7, regroupV0_lo_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo_1 = {regroupV0_lo_6[1547:1546], regroupV0_lo_6[1539:1538]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi_1 = {regroupV0_lo_6[1563:1562], regroupV0_lo_6[1555:1554]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_5 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi_1, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo_1 = {regroupV0_lo_6[1579:1578], regroupV0_lo_6[1571:1570]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi_1 = {regroupV0_lo_6[1595:1594], regroupV0_lo_6[1587:1586]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_5 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi_1, regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_lo_lo_7 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_5, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_5};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo_1 = {regroupV0_lo_6[1611:1610], regroupV0_lo_6[1603:1602]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi_1 = {regroupV0_lo_6[1627:1626], regroupV0_lo_6[1619:1618]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_5 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi_1, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo_1 = {regroupV0_lo_6[1643:1642], regroupV0_lo_6[1635:1634]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi_1 = {regroupV0_lo_6[1659:1658], regroupV0_lo_6[1651:1650]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_5 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi_1, regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_lo_hi_7 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_5, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_5};
  wire [31:0]        regroupV0_lo_lo_hi_hi_lo_lo_7 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_7, regroupV0_lo_lo_hi_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo_1 = {regroupV0_lo_6[1675:1674], regroupV0_lo_6[1667:1666]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi_1 = {regroupV0_lo_6[1691:1690], regroupV0_lo_6[1683:1682]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_5 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi_1, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo_1 = {regroupV0_lo_6[1707:1706], regroupV0_lo_6[1699:1698]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi_1 = {regroupV0_lo_6[1723:1722], regroupV0_lo_6[1715:1714]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_5 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi_1, regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_hi_lo_7 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_5, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_5};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo_1 = {regroupV0_lo_6[1739:1738], regroupV0_lo_6[1731:1730]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi_1 = {regroupV0_lo_6[1755:1754], regroupV0_lo_6[1747:1746]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_5 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi_1, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo_1 = {regroupV0_lo_6[1771:1770], regroupV0_lo_6[1763:1762]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi_1 = {regroupV0_lo_6[1787:1786], regroupV0_lo_6[1779:1778]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_5 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi_1, regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_hi_hi_7 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_5, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_5};
  wire [31:0]        regroupV0_lo_lo_hi_hi_lo_hi_7 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_7, regroupV0_lo_lo_hi_hi_lo_hi_lo_7};
  wire [63:0]        regroupV0_lo_lo_hi_hi_lo_7 = {regroupV0_lo_lo_hi_hi_lo_hi_7, regroupV0_lo_lo_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo_1 = {regroupV0_lo_6[1803:1802], regroupV0_lo_6[1795:1794]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi_1 = {regroupV0_lo_6[1819:1818], regroupV0_lo_6[1811:1810]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_5 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi_1, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo_1 = {regroupV0_lo_6[1835:1834], regroupV0_lo_6[1827:1826]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi_1 = {regroupV0_lo_6[1851:1850], regroupV0_lo_6[1843:1842]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_5 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi_1, regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_lo_lo_7 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_5, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_5};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo_1 = {regroupV0_lo_6[1867:1866], regroupV0_lo_6[1859:1858]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi_1 = {regroupV0_lo_6[1883:1882], regroupV0_lo_6[1875:1874]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_5 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi_1, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo_1 = {regroupV0_lo_6[1899:1898], regroupV0_lo_6[1891:1890]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi_1 = {regroupV0_lo_6[1915:1914], regroupV0_lo_6[1907:1906]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_5 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi_1, regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_lo_hi_7 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_5, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_5};
  wire [31:0]        regroupV0_lo_lo_hi_hi_hi_lo_7 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_7, regroupV0_lo_lo_hi_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo_1 = {regroupV0_lo_6[1931:1930], regroupV0_lo_6[1923:1922]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi_1 = {regroupV0_lo_6[1947:1946], regroupV0_lo_6[1939:1938]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_5 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi_1, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo_1 = {regroupV0_lo_6[1963:1962], regroupV0_lo_6[1955:1954]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi_1 = {regroupV0_lo_6[1979:1978], regroupV0_lo_6[1971:1970]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_5 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi_1, regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_hi_lo_7 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_5, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_5};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo_1 = {regroupV0_lo_6[1995:1994], regroupV0_lo_6[1987:1986]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi_1 = {regroupV0_lo_6[2011:2010], regroupV0_lo_6[2003:2002]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_5 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi_1, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo_1 = {regroupV0_lo_6[2027:2026], regroupV0_lo_6[2019:2018]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi_1 = {regroupV0_lo_6[2043:2042], regroupV0_lo_6[2035:2034]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_5 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi_1, regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_hi_hi_7 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_5, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_5};
  wire [31:0]        regroupV0_lo_lo_hi_hi_hi_hi_7 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_7, regroupV0_lo_lo_hi_hi_hi_hi_lo_7};
  wire [63:0]        regroupV0_lo_lo_hi_hi_hi_7 = {regroupV0_lo_lo_hi_hi_hi_hi_7, regroupV0_lo_lo_hi_hi_hi_lo_7};
  wire [127:0]       regroupV0_lo_lo_hi_hi_7 = {regroupV0_lo_lo_hi_hi_hi_7, regroupV0_lo_lo_hi_hi_lo_7};
  wire [255:0]       regroupV0_lo_lo_hi_7 = {regroupV0_lo_lo_hi_hi_7, regroupV0_lo_lo_hi_lo_7};
  wire [511:0]       regroupV0_lo_lo_7 = {regroupV0_lo_lo_hi_7, regroupV0_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo_1 = {regroupV0_lo_6[2059:2058], regroupV0_lo_6[2051:2050]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi_1 = {regroupV0_lo_6[2075:2074], regroupV0_lo_6[2067:2066]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_5 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi_1, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo_1 = {regroupV0_lo_6[2091:2090], regroupV0_lo_6[2083:2082]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi_1 = {regroupV0_lo_6[2107:2106], regroupV0_lo_6[2099:2098]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_5 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi_1, regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_lo_lo_7 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_5, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_5};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo_1 = {regroupV0_lo_6[2123:2122], regroupV0_lo_6[2115:2114]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi_1 = {regroupV0_lo_6[2139:2138], regroupV0_lo_6[2131:2130]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_5 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi_1, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo_1 = {regroupV0_lo_6[2155:2154], regroupV0_lo_6[2147:2146]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi_1 = {regroupV0_lo_6[2171:2170], regroupV0_lo_6[2163:2162]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_5 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi_1, regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_lo_hi_7 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_5, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_5};
  wire [31:0]        regroupV0_lo_hi_lo_lo_lo_lo_7 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_7, regroupV0_lo_hi_lo_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo_1 = {regroupV0_lo_6[2187:2186], regroupV0_lo_6[2179:2178]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi_1 = {regroupV0_lo_6[2203:2202], regroupV0_lo_6[2195:2194]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_5 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi_1, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo_1 = {regroupV0_lo_6[2219:2218], regroupV0_lo_6[2211:2210]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi_1 = {regroupV0_lo_6[2235:2234], regroupV0_lo_6[2227:2226]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_5 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi_1, regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_hi_lo_7 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_5, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_5};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo_1 = {regroupV0_lo_6[2251:2250], regroupV0_lo_6[2243:2242]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi_1 = {regroupV0_lo_6[2267:2266], regroupV0_lo_6[2259:2258]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_5 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi_1, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo_1 = {regroupV0_lo_6[2283:2282], regroupV0_lo_6[2275:2274]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi_1 = {regroupV0_lo_6[2299:2298], regroupV0_lo_6[2291:2290]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_5 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi_1, regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_hi_hi_7 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_5, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_5};
  wire [31:0]        regroupV0_lo_hi_lo_lo_lo_hi_7 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_7, regroupV0_lo_hi_lo_lo_lo_hi_lo_7};
  wire [63:0]        regroupV0_lo_hi_lo_lo_lo_7 = {regroupV0_lo_hi_lo_lo_lo_hi_7, regroupV0_lo_hi_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo_1 = {regroupV0_lo_6[2315:2314], regroupV0_lo_6[2307:2306]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi_1 = {regroupV0_lo_6[2331:2330], regroupV0_lo_6[2323:2322]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_5 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi_1, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo_1 = {regroupV0_lo_6[2347:2346], regroupV0_lo_6[2339:2338]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi_1 = {regroupV0_lo_6[2363:2362], regroupV0_lo_6[2355:2354]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_5 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi_1, regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_lo_lo_7 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_5, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_5};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo_1 = {regroupV0_lo_6[2379:2378], regroupV0_lo_6[2371:2370]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi_1 = {regroupV0_lo_6[2395:2394], regroupV0_lo_6[2387:2386]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_5 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi_1, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo_1 = {regroupV0_lo_6[2411:2410], regroupV0_lo_6[2403:2402]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi_1 = {regroupV0_lo_6[2427:2426], regroupV0_lo_6[2419:2418]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_5 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi_1, regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_lo_hi_7 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_5, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_5};
  wire [31:0]        regroupV0_lo_hi_lo_lo_hi_lo_7 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_7, regroupV0_lo_hi_lo_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo_1 = {regroupV0_lo_6[2443:2442], regroupV0_lo_6[2435:2434]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi_1 = {regroupV0_lo_6[2459:2458], regroupV0_lo_6[2451:2450]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_5 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi_1, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo_1 = {regroupV0_lo_6[2475:2474], regroupV0_lo_6[2467:2466]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi_1 = {regroupV0_lo_6[2491:2490], regroupV0_lo_6[2483:2482]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_5 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi_1, regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_hi_lo_7 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_5, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_5};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo_1 = {regroupV0_lo_6[2507:2506], regroupV0_lo_6[2499:2498]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi_1 = {regroupV0_lo_6[2523:2522], regroupV0_lo_6[2515:2514]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_5 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi_1, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo_1 = {regroupV0_lo_6[2539:2538], regroupV0_lo_6[2531:2530]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi_1 = {regroupV0_lo_6[2555:2554], regroupV0_lo_6[2547:2546]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_5 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi_1, regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_hi_hi_7 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_5, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_5};
  wire [31:0]        regroupV0_lo_hi_lo_lo_hi_hi_7 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_7, regroupV0_lo_hi_lo_lo_hi_hi_lo_7};
  wire [63:0]        regroupV0_lo_hi_lo_lo_hi_7 = {regroupV0_lo_hi_lo_lo_hi_hi_7, regroupV0_lo_hi_lo_lo_hi_lo_7};
  wire [127:0]       regroupV0_lo_hi_lo_lo_7 = {regroupV0_lo_hi_lo_lo_hi_7, regroupV0_lo_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo_1 = {regroupV0_lo_6[2571:2570], regroupV0_lo_6[2563:2562]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi_1 = {regroupV0_lo_6[2587:2586], regroupV0_lo_6[2579:2578]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_5 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi_1, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo_1 = {regroupV0_lo_6[2603:2602], regroupV0_lo_6[2595:2594]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi_1 = {regroupV0_lo_6[2619:2618], regroupV0_lo_6[2611:2610]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_5 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi_1, regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_lo_lo_7 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_5, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_5};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo_1 = {regroupV0_lo_6[2635:2634], regroupV0_lo_6[2627:2626]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi_1 = {regroupV0_lo_6[2651:2650], regroupV0_lo_6[2643:2642]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_5 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi_1, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo_1 = {regroupV0_lo_6[2667:2666], regroupV0_lo_6[2659:2658]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi_1 = {regroupV0_lo_6[2683:2682], regroupV0_lo_6[2675:2674]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_5 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi_1, regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_lo_hi_7 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_5, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_5};
  wire [31:0]        regroupV0_lo_hi_lo_hi_lo_lo_7 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_7, regroupV0_lo_hi_lo_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo_1 = {regroupV0_lo_6[2699:2698], regroupV0_lo_6[2691:2690]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi_1 = {regroupV0_lo_6[2715:2714], regroupV0_lo_6[2707:2706]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_5 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi_1, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo_1 = {regroupV0_lo_6[2731:2730], regroupV0_lo_6[2723:2722]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi_1 = {regroupV0_lo_6[2747:2746], regroupV0_lo_6[2739:2738]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_5 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi_1, regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_hi_lo_7 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_5, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_5};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo_1 = {regroupV0_lo_6[2763:2762], regroupV0_lo_6[2755:2754]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi_1 = {regroupV0_lo_6[2779:2778], regroupV0_lo_6[2771:2770]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_5 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi_1, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo_1 = {regroupV0_lo_6[2795:2794], regroupV0_lo_6[2787:2786]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi_1 = {regroupV0_lo_6[2811:2810], regroupV0_lo_6[2803:2802]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_5 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi_1, regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_hi_hi_7 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_5, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_5};
  wire [31:0]        regroupV0_lo_hi_lo_hi_lo_hi_7 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_7, regroupV0_lo_hi_lo_hi_lo_hi_lo_7};
  wire [63:0]        regroupV0_lo_hi_lo_hi_lo_7 = {regroupV0_lo_hi_lo_hi_lo_hi_7, regroupV0_lo_hi_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo_1 = {regroupV0_lo_6[2827:2826], regroupV0_lo_6[2819:2818]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi_1 = {regroupV0_lo_6[2843:2842], regroupV0_lo_6[2835:2834]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_5 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi_1, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo_1 = {regroupV0_lo_6[2859:2858], regroupV0_lo_6[2851:2850]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi_1 = {regroupV0_lo_6[2875:2874], regroupV0_lo_6[2867:2866]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_5 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi_1, regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_lo_lo_7 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_5, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_5};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo_1 = {regroupV0_lo_6[2891:2890], regroupV0_lo_6[2883:2882]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi_1 = {regroupV0_lo_6[2907:2906], regroupV0_lo_6[2899:2898]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_5 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi_1, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo_1 = {regroupV0_lo_6[2923:2922], regroupV0_lo_6[2915:2914]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi_1 = {regroupV0_lo_6[2939:2938], regroupV0_lo_6[2931:2930]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_5 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi_1, regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_lo_hi_7 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_5, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_5};
  wire [31:0]        regroupV0_lo_hi_lo_hi_hi_lo_7 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_7, regroupV0_lo_hi_lo_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo_1 = {regroupV0_lo_6[2955:2954], regroupV0_lo_6[2947:2946]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi_1 = {regroupV0_lo_6[2971:2970], regroupV0_lo_6[2963:2962]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_5 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi_1, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo_1 = {regroupV0_lo_6[2987:2986], regroupV0_lo_6[2979:2978]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi_1 = {regroupV0_lo_6[3003:3002], regroupV0_lo_6[2995:2994]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_5 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi_1, regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_hi_lo_7 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_5, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_5};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo_1 = {regroupV0_lo_6[3019:3018], regroupV0_lo_6[3011:3010]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi_1 = {regroupV0_lo_6[3035:3034], regroupV0_lo_6[3027:3026]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_5 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi_1, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo_1 = {regroupV0_lo_6[3051:3050], regroupV0_lo_6[3043:3042]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi_1 = {regroupV0_lo_6[3067:3066], regroupV0_lo_6[3059:3058]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_5 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi_1, regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_hi_hi_7 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_5, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_5};
  wire [31:0]        regroupV0_lo_hi_lo_hi_hi_hi_7 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_7, regroupV0_lo_hi_lo_hi_hi_hi_lo_7};
  wire [63:0]        regroupV0_lo_hi_lo_hi_hi_7 = {regroupV0_lo_hi_lo_hi_hi_hi_7, regroupV0_lo_hi_lo_hi_hi_lo_7};
  wire [127:0]       regroupV0_lo_hi_lo_hi_7 = {regroupV0_lo_hi_lo_hi_hi_7, regroupV0_lo_hi_lo_hi_lo_7};
  wire [255:0]       regroupV0_lo_hi_lo_7 = {regroupV0_lo_hi_lo_hi_7, regroupV0_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo_1 = {regroupV0_lo_6[3083:3082], regroupV0_lo_6[3075:3074]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi_1 = {regroupV0_lo_6[3099:3098], regroupV0_lo_6[3091:3090]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_5 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi_1, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo_1 = {regroupV0_lo_6[3115:3114], regroupV0_lo_6[3107:3106]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi_1 = {regroupV0_lo_6[3131:3130], regroupV0_lo_6[3123:3122]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_5 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi_1, regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_lo_lo_7 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_5, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_5};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo_1 = {regroupV0_lo_6[3147:3146], regroupV0_lo_6[3139:3138]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi_1 = {regroupV0_lo_6[3163:3162], regroupV0_lo_6[3155:3154]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_5 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi_1, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo_1 = {regroupV0_lo_6[3179:3178], regroupV0_lo_6[3171:3170]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi_1 = {regroupV0_lo_6[3195:3194], regroupV0_lo_6[3187:3186]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_5 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi_1, regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_lo_hi_7 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_5, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_5};
  wire [31:0]        regroupV0_lo_hi_hi_lo_lo_lo_7 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_7, regroupV0_lo_hi_hi_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo_1 = {regroupV0_lo_6[3211:3210], regroupV0_lo_6[3203:3202]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi_1 = {regroupV0_lo_6[3227:3226], regroupV0_lo_6[3219:3218]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_5 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi_1, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo_1 = {regroupV0_lo_6[3243:3242], regroupV0_lo_6[3235:3234]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi_1 = {regroupV0_lo_6[3259:3258], regroupV0_lo_6[3251:3250]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_5 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi_1, regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_hi_lo_7 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_5, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_5};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo_1 = {regroupV0_lo_6[3275:3274], regroupV0_lo_6[3267:3266]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi_1 = {regroupV0_lo_6[3291:3290], regroupV0_lo_6[3283:3282]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_5 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi_1, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo_1 = {regroupV0_lo_6[3307:3306], regroupV0_lo_6[3299:3298]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi_1 = {regroupV0_lo_6[3323:3322], regroupV0_lo_6[3315:3314]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_5 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi_1, regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_hi_hi_7 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_5, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_5};
  wire [31:0]        regroupV0_lo_hi_hi_lo_lo_hi_7 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_7, regroupV0_lo_hi_hi_lo_lo_hi_lo_7};
  wire [63:0]        regroupV0_lo_hi_hi_lo_lo_7 = {regroupV0_lo_hi_hi_lo_lo_hi_7, regroupV0_lo_hi_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo_1 = {regroupV0_lo_6[3339:3338], regroupV0_lo_6[3331:3330]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi_1 = {regroupV0_lo_6[3355:3354], regroupV0_lo_6[3347:3346]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_5 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi_1, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo_1 = {regroupV0_lo_6[3371:3370], regroupV0_lo_6[3363:3362]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi_1 = {regroupV0_lo_6[3387:3386], regroupV0_lo_6[3379:3378]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_5 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi_1, regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_lo_lo_7 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_5, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_5};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo_1 = {regroupV0_lo_6[3403:3402], regroupV0_lo_6[3395:3394]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi_1 = {regroupV0_lo_6[3419:3418], regroupV0_lo_6[3411:3410]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_5 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi_1, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo_1 = {regroupV0_lo_6[3435:3434], regroupV0_lo_6[3427:3426]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi_1 = {regroupV0_lo_6[3451:3450], regroupV0_lo_6[3443:3442]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_5 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi_1, regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_lo_hi_7 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_5, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_5};
  wire [31:0]        regroupV0_lo_hi_hi_lo_hi_lo_7 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_7, regroupV0_lo_hi_hi_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo_1 = {regroupV0_lo_6[3467:3466], regroupV0_lo_6[3459:3458]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi_1 = {regroupV0_lo_6[3483:3482], regroupV0_lo_6[3475:3474]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_5 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi_1, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo_1 = {regroupV0_lo_6[3499:3498], regroupV0_lo_6[3491:3490]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi_1 = {regroupV0_lo_6[3515:3514], regroupV0_lo_6[3507:3506]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_5 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi_1, regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_hi_lo_7 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_5, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_5};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo_1 = {regroupV0_lo_6[3531:3530], regroupV0_lo_6[3523:3522]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi_1 = {regroupV0_lo_6[3547:3546], regroupV0_lo_6[3539:3538]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_5 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi_1, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo_1 = {regroupV0_lo_6[3563:3562], regroupV0_lo_6[3555:3554]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi_1 = {regroupV0_lo_6[3579:3578], regroupV0_lo_6[3571:3570]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_5 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi_1, regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_hi_hi_7 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_5, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_5};
  wire [31:0]        regroupV0_lo_hi_hi_lo_hi_hi_7 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_7, regroupV0_lo_hi_hi_lo_hi_hi_lo_7};
  wire [63:0]        regroupV0_lo_hi_hi_lo_hi_7 = {regroupV0_lo_hi_hi_lo_hi_hi_7, regroupV0_lo_hi_hi_lo_hi_lo_7};
  wire [127:0]       regroupV0_lo_hi_hi_lo_7 = {regroupV0_lo_hi_hi_lo_hi_7, regroupV0_lo_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo_1 = {regroupV0_lo_6[3595:3594], regroupV0_lo_6[3587:3586]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi_1 = {regroupV0_lo_6[3611:3610], regroupV0_lo_6[3603:3602]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_5 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi_1, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo_1 = {regroupV0_lo_6[3627:3626], regroupV0_lo_6[3619:3618]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi_1 = {regroupV0_lo_6[3643:3642], regroupV0_lo_6[3635:3634]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_5 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi_1, regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_lo_lo_7 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_5, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_5};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo_1 = {regroupV0_lo_6[3659:3658], regroupV0_lo_6[3651:3650]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi_1 = {regroupV0_lo_6[3675:3674], regroupV0_lo_6[3667:3666]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_5 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi_1, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo_1 = {regroupV0_lo_6[3691:3690], regroupV0_lo_6[3683:3682]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi_1 = {regroupV0_lo_6[3707:3706], regroupV0_lo_6[3699:3698]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_5 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi_1, regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_lo_hi_7 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_5, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_5};
  wire [31:0]        regroupV0_lo_hi_hi_hi_lo_lo_7 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_7, regroupV0_lo_hi_hi_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo_1 = {regroupV0_lo_6[3723:3722], regroupV0_lo_6[3715:3714]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi_1 = {regroupV0_lo_6[3739:3738], regroupV0_lo_6[3731:3730]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_5 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi_1, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo_1 = {regroupV0_lo_6[3755:3754], regroupV0_lo_6[3747:3746]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi_1 = {regroupV0_lo_6[3771:3770], regroupV0_lo_6[3763:3762]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_5 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi_1, regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_hi_lo_7 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_5, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_5};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo_1 = {regroupV0_lo_6[3787:3786], regroupV0_lo_6[3779:3778]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi_1 = {regroupV0_lo_6[3803:3802], regroupV0_lo_6[3795:3794]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_5 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi_1, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo_1 = {regroupV0_lo_6[3819:3818], regroupV0_lo_6[3811:3810]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi_1 = {regroupV0_lo_6[3835:3834], regroupV0_lo_6[3827:3826]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_5 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi_1, regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_hi_hi_7 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_5, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_5};
  wire [31:0]        regroupV0_lo_hi_hi_hi_lo_hi_7 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_7, regroupV0_lo_hi_hi_hi_lo_hi_lo_7};
  wire [63:0]        regroupV0_lo_hi_hi_hi_lo_7 = {regroupV0_lo_hi_hi_hi_lo_hi_7, regroupV0_lo_hi_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo_1 = {regroupV0_lo_6[3851:3850], regroupV0_lo_6[3843:3842]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi_1 = {regroupV0_lo_6[3867:3866], regroupV0_lo_6[3859:3858]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_5 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi_1, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo_1 = {regroupV0_lo_6[3883:3882], regroupV0_lo_6[3875:3874]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi_1 = {regroupV0_lo_6[3899:3898], regroupV0_lo_6[3891:3890]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_5 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi_1, regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_lo_lo_7 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_5, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_5};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo_1 = {regroupV0_lo_6[3915:3914], regroupV0_lo_6[3907:3906]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi_1 = {regroupV0_lo_6[3931:3930], regroupV0_lo_6[3923:3922]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_5 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi_1, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo_1 = {regroupV0_lo_6[3947:3946], regroupV0_lo_6[3939:3938]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi_1 = {regroupV0_lo_6[3963:3962], regroupV0_lo_6[3955:3954]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_5 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi_1, regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_lo_hi_7 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_5, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_5};
  wire [31:0]        regroupV0_lo_hi_hi_hi_hi_lo_7 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_7, regroupV0_lo_hi_hi_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo_1 = {regroupV0_lo_6[3979:3978], regroupV0_lo_6[3971:3970]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi_1 = {regroupV0_lo_6[3995:3994], regroupV0_lo_6[3987:3986]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_5 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi_1, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo_1 = {regroupV0_lo_6[4011:4010], regroupV0_lo_6[4003:4002]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi_1 = {regroupV0_lo_6[4027:4026], regroupV0_lo_6[4019:4018]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_5 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi_1, regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_hi_lo_7 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_5, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_5};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo_1 = {regroupV0_lo_6[4043:4042], regroupV0_lo_6[4035:4034]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi_1 = {regroupV0_lo_6[4059:4058], regroupV0_lo_6[4051:4050]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_5 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi_1, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo_1 = {regroupV0_lo_6[4075:4074], regroupV0_lo_6[4067:4066]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi_1 = {regroupV0_lo_6[4091:4090], regroupV0_lo_6[4083:4082]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_5 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi_1, regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_hi_hi_7 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_5, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_5};
  wire [31:0]        regroupV0_lo_hi_hi_hi_hi_hi_7 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_7, regroupV0_lo_hi_hi_hi_hi_hi_lo_7};
  wire [63:0]        regroupV0_lo_hi_hi_hi_hi_7 = {regroupV0_lo_hi_hi_hi_hi_hi_7, regroupV0_lo_hi_hi_hi_hi_lo_7};
  wire [127:0]       regroupV0_lo_hi_hi_hi_7 = {regroupV0_lo_hi_hi_hi_hi_7, regroupV0_lo_hi_hi_hi_lo_7};
  wire [255:0]       regroupV0_lo_hi_hi_7 = {regroupV0_lo_hi_hi_hi_7, regroupV0_lo_hi_hi_lo_7};
  wire [511:0]       regroupV0_lo_hi_7 = {regroupV0_lo_hi_hi_7, regroupV0_lo_hi_lo_7};
  wire [1023:0]      regroupV0_lo_8 = {regroupV0_lo_hi_7, regroupV0_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo_1 = {regroupV0_hi_6[11:10], regroupV0_hi_6[3:2]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi_1 = {regroupV0_hi_6[27:26], regroupV0_hi_6[19:18]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_5 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo_1 = {regroupV0_hi_6[43:42], regroupV0_hi_6[35:34]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi_1 = {regroupV0_hi_6[59:58], regroupV0_hi_6[51:50]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_5 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi_1, regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_lo_lo_7 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_5, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_5};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo_1 = {regroupV0_hi_6[75:74], regroupV0_hi_6[67:66]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi_1 = {regroupV0_hi_6[91:90], regroupV0_hi_6[83:82]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_5 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi_1, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo_1 = {regroupV0_hi_6[107:106], regroupV0_hi_6[99:98]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi_1 = {regroupV0_hi_6[123:122], regroupV0_hi_6[115:114]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_5 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi_1, regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_lo_hi_7 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_5, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_5};
  wire [31:0]        regroupV0_hi_lo_lo_lo_lo_lo_7 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_7, regroupV0_hi_lo_lo_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo_1 = {regroupV0_hi_6[139:138], regroupV0_hi_6[131:130]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi_1 = {regroupV0_hi_6[155:154], regroupV0_hi_6[147:146]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_5 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo_1 = {regroupV0_hi_6[171:170], regroupV0_hi_6[163:162]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi_1 = {regroupV0_hi_6[187:186], regroupV0_hi_6[179:178]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_5 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi_1, regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_hi_lo_7 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_5, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_5};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo_1 = {regroupV0_hi_6[203:202], regroupV0_hi_6[195:194]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi_1 = {regroupV0_hi_6[219:218], regroupV0_hi_6[211:210]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_5 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi_1, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo_1 = {regroupV0_hi_6[235:234], regroupV0_hi_6[227:226]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi_1 = {regroupV0_hi_6[251:250], regroupV0_hi_6[243:242]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_5 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi_1, regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_hi_hi_7 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_5, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_5};
  wire [31:0]        regroupV0_hi_lo_lo_lo_lo_hi_7 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_7, regroupV0_hi_lo_lo_lo_lo_hi_lo_7};
  wire [63:0]        regroupV0_hi_lo_lo_lo_lo_7 = {regroupV0_hi_lo_lo_lo_lo_hi_7, regroupV0_hi_lo_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo_1 = {regroupV0_hi_6[267:266], regroupV0_hi_6[259:258]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi_1 = {regroupV0_hi_6[283:282], regroupV0_hi_6[275:274]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_5 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo_1 = {regroupV0_hi_6[299:298], regroupV0_hi_6[291:290]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi_1 = {regroupV0_hi_6[315:314], regroupV0_hi_6[307:306]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_5 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi_1, regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_lo_lo_7 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_5, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_5};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo_1 = {regroupV0_hi_6[331:330], regroupV0_hi_6[323:322]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi_1 = {regroupV0_hi_6[347:346], regroupV0_hi_6[339:338]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_5 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi_1, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo_1 = {regroupV0_hi_6[363:362], regroupV0_hi_6[355:354]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi_1 = {regroupV0_hi_6[379:378], regroupV0_hi_6[371:370]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_5 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi_1, regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_lo_hi_7 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_5, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_5};
  wire [31:0]        regroupV0_hi_lo_lo_lo_hi_lo_7 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_7, regroupV0_hi_lo_lo_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo_1 = {regroupV0_hi_6[395:394], regroupV0_hi_6[387:386]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi_1 = {regroupV0_hi_6[411:410], regroupV0_hi_6[403:402]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_5 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo_1 = {regroupV0_hi_6[427:426], regroupV0_hi_6[419:418]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi_1 = {regroupV0_hi_6[443:442], regroupV0_hi_6[435:434]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_5 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi_1, regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_hi_lo_7 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_5, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_5};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo_1 = {regroupV0_hi_6[459:458], regroupV0_hi_6[451:450]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi_1 = {regroupV0_hi_6[475:474], regroupV0_hi_6[467:466]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_5 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi_1, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo_1 = {regroupV0_hi_6[491:490], regroupV0_hi_6[483:482]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi_1 = {regroupV0_hi_6[507:506], regroupV0_hi_6[499:498]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_5 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi_1, regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_hi_hi_7 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_5, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_5};
  wire [31:0]        regroupV0_hi_lo_lo_lo_hi_hi_7 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_7, regroupV0_hi_lo_lo_lo_hi_hi_lo_7};
  wire [63:0]        regroupV0_hi_lo_lo_lo_hi_7 = {regroupV0_hi_lo_lo_lo_hi_hi_7, regroupV0_hi_lo_lo_lo_hi_lo_7};
  wire [127:0]       regroupV0_hi_lo_lo_lo_7 = {regroupV0_hi_lo_lo_lo_hi_7, regroupV0_hi_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo_1 = {regroupV0_hi_6[523:522], regroupV0_hi_6[515:514]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi_1 = {regroupV0_hi_6[539:538], regroupV0_hi_6[531:530]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_5 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi_1, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo_1 = {regroupV0_hi_6[555:554], regroupV0_hi_6[547:546]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi_1 = {regroupV0_hi_6[571:570], regroupV0_hi_6[563:562]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_5 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi_1, regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_lo_lo_7 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_5, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_5};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo_1 = {regroupV0_hi_6[587:586], regroupV0_hi_6[579:578]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi_1 = {regroupV0_hi_6[603:602], regroupV0_hi_6[595:594]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_5 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi_1, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo_1 = {regroupV0_hi_6[619:618], regroupV0_hi_6[611:610]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi_1 = {regroupV0_hi_6[635:634], regroupV0_hi_6[627:626]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_5 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi_1, regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_lo_hi_7 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_5, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_5};
  wire [31:0]        regroupV0_hi_lo_lo_hi_lo_lo_7 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_7, regroupV0_hi_lo_lo_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo_1 = {regroupV0_hi_6[651:650], regroupV0_hi_6[643:642]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi_1 = {regroupV0_hi_6[667:666], regroupV0_hi_6[659:658]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_5 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi_1, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo_1 = {regroupV0_hi_6[683:682], regroupV0_hi_6[675:674]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi_1 = {regroupV0_hi_6[699:698], regroupV0_hi_6[691:690]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_5 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi_1, regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_hi_lo_7 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_5, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_5};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo_1 = {regroupV0_hi_6[715:714], regroupV0_hi_6[707:706]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi_1 = {regroupV0_hi_6[731:730], regroupV0_hi_6[723:722]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_5 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi_1, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo_1 = {regroupV0_hi_6[747:746], regroupV0_hi_6[739:738]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi_1 = {regroupV0_hi_6[763:762], regroupV0_hi_6[755:754]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_5 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi_1, regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_hi_hi_7 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_5, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_5};
  wire [31:0]        regroupV0_hi_lo_lo_hi_lo_hi_7 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_7, regroupV0_hi_lo_lo_hi_lo_hi_lo_7};
  wire [63:0]        regroupV0_hi_lo_lo_hi_lo_7 = {regroupV0_hi_lo_lo_hi_lo_hi_7, regroupV0_hi_lo_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo_1 = {regroupV0_hi_6[779:778], regroupV0_hi_6[771:770]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi_1 = {regroupV0_hi_6[795:794], regroupV0_hi_6[787:786]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_5 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi_1, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo_1 = {regroupV0_hi_6[811:810], regroupV0_hi_6[803:802]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi_1 = {regroupV0_hi_6[827:826], regroupV0_hi_6[819:818]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_5 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi_1, regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_lo_lo_7 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_5, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_5};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo_1 = {regroupV0_hi_6[843:842], regroupV0_hi_6[835:834]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi_1 = {regroupV0_hi_6[859:858], regroupV0_hi_6[851:850]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_5 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi_1, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo_1 = {regroupV0_hi_6[875:874], regroupV0_hi_6[867:866]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi_1 = {regroupV0_hi_6[891:890], regroupV0_hi_6[883:882]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_5 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi_1, regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_lo_hi_7 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_5, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_5};
  wire [31:0]        regroupV0_hi_lo_lo_hi_hi_lo_7 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_7, regroupV0_hi_lo_lo_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo_1 = {regroupV0_hi_6[907:906], regroupV0_hi_6[899:898]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi_1 = {regroupV0_hi_6[923:922], regroupV0_hi_6[915:914]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_5 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi_1, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo_1 = {regroupV0_hi_6[939:938], regroupV0_hi_6[931:930]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi_1 = {regroupV0_hi_6[955:954], regroupV0_hi_6[947:946]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_5 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi_1, regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_hi_lo_7 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_5, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_5};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo_1 = {regroupV0_hi_6[971:970], regroupV0_hi_6[963:962]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi_1 = {regroupV0_hi_6[987:986], regroupV0_hi_6[979:978]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_5 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi_1, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo_1 = {regroupV0_hi_6[1003:1002], regroupV0_hi_6[995:994]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi_1 = {regroupV0_hi_6[1019:1018], regroupV0_hi_6[1011:1010]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_5 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi_1, regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_hi_hi_7 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_5, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_5};
  wire [31:0]        regroupV0_hi_lo_lo_hi_hi_hi_7 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_7, regroupV0_hi_lo_lo_hi_hi_hi_lo_7};
  wire [63:0]        regroupV0_hi_lo_lo_hi_hi_7 = {regroupV0_hi_lo_lo_hi_hi_hi_7, regroupV0_hi_lo_lo_hi_hi_lo_7};
  wire [127:0]       regroupV0_hi_lo_lo_hi_7 = {regroupV0_hi_lo_lo_hi_hi_7, regroupV0_hi_lo_lo_hi_lo_7};
  wire [255:0]       regroupV0_hi_lo_lo_7 = {regroupV0_hi_lo_lo_hi_7, regroupV0_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo_1 = {regroupV0_hi_6[1035:1034], regroupV0_hi_6[1027:1026]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi_1 = {regroupV0_hi_6[1051:1050], regroupV0_hi_6[1043:1042]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_5 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi_1, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo_1 = {regroupV0_hi_6[1067:1066], regroupV0_hi_6[1059:1058]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi_1 = {regroupV0_hi_6[1083:1082], regroupV0_hi_6[1075:1074]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_5 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi_1, regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_lo_lo_7 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_5, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_5};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo_1 = {regroupV0_hi_6[1099:1098], regroupV0_hi_6[1091:1090]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi_1 = {regroupV0_hi_6[1115:1114], regroupV0_hi_6[1107:1106]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_5 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi_1, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo_1 = {regroupV0_hi_6[1131:1130], regroupV0_hi_6[1123:1122]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi_1 = {regroupV0_hi_6[1147:1146], regroupV0_hi_6[1139:1138]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_5 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi_1, regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_lo_hi_7 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_5, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_5};
  wire [31:0]        regroupV0_hi_lo_hi_lo_lo_lo_7 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_7, regroupV0_hi_lo_hi_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo_1 = {regroupV0_hi_6[1163:1162], regroupV0_hi_6[1155:1154]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi_1 = {regroupV0_hi_6[1179:1178], regroupV0_hi_6[1171:1170]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_5 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi_1, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo_1 = {regroupV0_hi_6[1195:1194], regroupV0_hi_6[1187:1186]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi_1 = {regroupV0_hi_6[1211:1210], regroupV0_hi_6[1203:1202]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_5 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi_1, regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_hi_lo_7 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_5, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_5};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo_1 = {regroupV0_hi_6[1227:1226], regroupV0_hi_6[1219:1218]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi_1 = {regroupV0_hi_6[1243:1242], regroupV0_hi_6[1235:1234]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_5 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi_1, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo_1 = {regroupV0_hi_6[1259:1258], regroupV0_hi_6[1251:1250]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi_1 = {regroupV0_hi_6[1275:1274], regroupV0_hi_6[1267:1266]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_5 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi_1, regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_hi_hi_7 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_5, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_5};
  wire [31:0]        regroupV0_hi_lo_hi_lo_lo_hi_7 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_7, regroupV0_hi_lo_hi_lo_lo_hi_lo_7};
  wire [63:0]        regroupV0_hi_lo_hi_lo_lo_7 = {regroupV0_hi_lo_hi_lo_lo_hi_7, regroupV0_hi_lo_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo_1 = {regroupV0_hi_6[1291:1290], regroupV0_hi_6[1283:1282]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi_1 = {regroupV0_hi_6[1307:1306], regroupV0_hi_6[1299:1298]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_5 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi_1, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo_1 = {regroupV0_hi_6[1323:1322], regroupV0_hi_6[1315:1314]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi_1 = {regroupV0_hi_6[1339:1338], regroupV0_hi_6[1331:1330]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_5 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi_1, regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_lo_lo_7 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_5, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_5};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo_1 = {regroupV0_hi_6[1355:1354], regroupV0_hi_6[1347:1346]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi_1 = {regroupV0_hi_6[1371:1370], regroupV0_hi_6[1363:1362]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_5 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi_1, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo_1 = {regroupV0_hi_6[1387:1386], regroupV0_hi_6[1379:1378]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi_1 = {regroupV0_hi_6[1403:1402], regroupV0_hi_6[1395:1394]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_5 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi_1, regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_lo_hi_7 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_5, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_5};
  wire [31:0]        regroupV0_hi_lo_hi_lo_hi_lo_7 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_7, regroupV0_hi_lo_hi_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo_1 = {regroupV0_hi_6[1419:1418], regroupV0_hi_6[1411:1410]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi_1 = {regroupV0_hi_6[1435:1434], regroupV0_hi_6[1427:1426]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_5 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi_1, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo_1 = {regroupV0_hi_6[1451:1450], regroupV0_hi_6[1443:1442]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi_1 = {regroupV0_hi_6[1467:1466], regroupV0_hi_6[1459:1458]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_5 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi_1, regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_hi_lo_7 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_5, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_5};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo_1 = {regroupV0_hi_6[1483:1482], regroupV0_hi_6[1475:1474]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi_1 = {regroupV0_hi_6[1499:1498], regroupV0_hi_6[1491:1490]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_5 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi_1, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo_1 = {regroupV0_hi_6[1515:1514], regroupV0_hi_6[1507:1506]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi_1 = {regroupV0_hi_6[1531:1530], regroupV0_hi_6[1523:1522]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_5 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi_1, regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_hi_hi_7 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_5, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_5};
  wire [31:0]        regroupV0_hi_lo_hi_lo_hi_hi_7 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_7, regroupV0_hi_lo_hi_lo_hi_hi_lo_7};
  wire [63:0]        regroupV0_hi_lo_hi_lo_hi_7 = {regroupV0_hi_lo_hi_lo_hi_hi_7, regroupV0_hi_lo_hi_lo_hi_lo_7};
  wire [127:0]       regroupV0_hi_lo_hi_lo_7 = {regroupV0_hi_lo_hi_lo_hi_7, regroupV0_hi_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo_1 = {regroupV0_hi_6[1547:1546], regroupV0_hi_6[1539:1538]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi_1 = {regroupV0_hi_6[1563:1562], regroupV0_hi_6[1555:1554]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_5 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi_1, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo_1 = {regroupV0_hi_6[1579:1578], regroupV0_hi_6[1571:1570]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi_1 = {regroupV0_hi_6[1595:1594], regroupV0_hi_6[1587:1586]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_5 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi_1, regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_lo_lo_7 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_5, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_5};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo_1 = {regroupV0_hi_6[1611:1610], regroupV0_hi_6[1603:1602]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi_1 = {regroupV0_hi_6[1627:1626], regroupV0_hi_6[1619:1618]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_5 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi_1, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo_1 = {regroupV0_hi_6[1643:1642], regroupV0_hi_6[1635:1634]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi_1 = {regroupV0_hi_6[1659:1658], regroupV0_hi_6[1651:1650]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_5 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi_1, regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_lo_hi_7 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_5, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_5};
  wire [31:0]        regroupV0_hi_lo_hi_hi_lo_lo_7 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_7, regroupV0_hi_lo_hi_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo_1 = {regroupV0_hi_6[1675:1674], regroupV0_hi_6[1667:1666]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi_1 = {regroupV0_hi_6[1691:1690], regroupV0_hi_6[1683:1682]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_5 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi_1, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo_1 = {regroupV0_hi_6[1707:1706], regroupV0_hi_6[1699:1698]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi_1 = {regroupV0_hi_6[1723:1722], regroupV0_hi_6[1715:1714]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_5 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi_1, regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_hi_lo_7 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_5, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_5};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo_1 = {regroupV0_hi_6[1739:1738], regroupV0_hi_6[1731:1730]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi_1 = {regroupV0_hi_6[1755:1754], regroupV0_hi_6[1747:1746]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_5 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi_1, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo_1 = {regroupV0_hi_6[1771:1770], regroupV0_hi_6[1763:1762]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi_1 = {regroupV0_hi_6[1787:1786], regroupV0_hi_6[1779:1778]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_5 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi_1, regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_hi_hi_7 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_5, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_5};
  wire [31:0]        regroupV0_hi_lo_hi_hi_lo_hi_7 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_7, regroupV0_hi_lo_hi_hi_lo_hi_lo_7};
  wire [63:0]        regroupV0_hi_lo_hi_hi_lo_7 = {regroupV0_hi_lo_hi_hi_lo_hi_7, regroupV0_hi_lo_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo_1 = {regroupV0_hi_6[1803:1802], regroupV0_hi_6[1795:1794]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi_1 = {regroupV0_hi_6[1819:1818], regroupV0_hi_6[1811:1810]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_5 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi_1, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo_1 = {regroupV0_hi_6[1835:1834], regroupV0_hi_6[1827:1826]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi_1 = {regroupV0_hi_6[1851:1850], regroupV0_hi_6[1843:1842]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_5 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi_1, regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_lo_lo_7 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_5, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_5};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo_1 = {regroupV0_hi_6[1867:1866], regroupV0_hi_6[1859:1858]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi_1 = {regroupV0_hi_6[1883:1882], regroupV0_hi_6[1875:1874]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_5 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi_1, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo_1 = {regroupV0_hi_6[1899:1898], regroupV0_hi_6[1891:1890]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi_1 = {regroupV0_hi_6[1915:1914], regroupV0_hi_6[1907:1906]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_5 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi_1, regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_lo_hi_7 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_5, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_5};
  wire [31:0]        regroupV0_hi_lo_hi_hi_hi_lo_7 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_7, regroupV0_hi_lo_hi_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo_1 = {regroupV0_hi_6[1931:1930], regroupV0_hi_6[1923:1922]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi_1 = {regroupV0_hi_6[1947:1946], regroupV0_hi_6[1939:1938]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_5 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi_1, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo_1 = {regroupV0_hi_6[1963:1962], regroupV0_hi_6[1955:1954]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi_1 = {regroupV0_hi_6[1979:1978], regroupV0_hi_6[1971:1970]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_5 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi_1, regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_hi_lo_7 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_5, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_5};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo_1 = {regroupV0_hi_6[1995:1994], regroupV0_hi_6[1987:1986]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi_1 = {regroupV0_hi_6[2011:2010], regroupV0_hi_6[2003:2002]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_5 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi_1, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo_1 = {regroupV0_hi_6[2027:2026], regroupV0_hi_6[2019:2018]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi_1 = {regroupV0_hi_6[2043:2042], regroupV0_hi_6[2035:2034]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_5 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi_1, regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_hi_hi_7 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_5, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_5};
  wire [31:0]        regroupV0_hi_lo_hi_hi_hi_hi_7 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_7, regroupV0_hi_lo_hi_hi_hi_hi_lo_7};
  wire [63:0]        regroupV0_hi_lo_hi_hi_hi_7 = {regroupV0_hi_lo_hi_hi_hi_hi_7, regroupV0_hi_lo_hi_hi_hi_lo_7};
  wire [127:0]       regroupV0_hi_lo_hi_hi_7 = {regroupV0_hi_lo_hi_hi_hi_7, regroupV0_hi_lo_hi_hi_lo_7};
  wire [255:0]       regroupV0_hi_lo_hi_7 = {regroupV0_hi_lo_hi_hi_7, regroupV0_hi_lo_hi_lo_7};
  wire [511:0]       regroupV0_hi_lo_7 = {regroupV0_hi_lo_hi_7, regroupV0_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo_1 = {regroupV0_hi_6[2059:2058], regroupV0_hi_6[2051:2050]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi_1 = {regroupV0_hi_6[2075:2074], regroupV0_hi_6[2067:2066]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_5 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi_1, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo_1 = {regroupV0_hi_6[2091:2090], regroupV0_hi_6[2083:2082]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi_1 = {regroupV0_hi_6[2107:2106], regroupV0_hi_6[2099:2098]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_5 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi_1, regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_lo_lo_7 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_5, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_5};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo_1 = {regroupV0_hi_6[2123:2122], regroupV0_hi_6[2115:2114]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi_1 = {regroupV0_hi_6[2139:2138], regroupV0_hi_6[2131:2130]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_5 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi_1, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo_1 = {regroupV0_hi_6[2155:2154], regroupV0_hi_6[2147:2146]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi_1 = {regroupV0_hi_6[2171:2170], regroupV0_hi_6[2163:2162]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_5 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi_1, regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_lo_hi_7 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_5, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_5};
  wire [31:0]        regroupV0_hi_hi_lo_lo_lo_lo_7 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_7, regroupV0_hi_hi_lo_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo_1 = {regroupV0_hi_6[2187:2186], regroupV0_hi_6[2179:2178]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi_1 = {regroupV0_hi_6[2203:2202], regroupV0_hi_6[2195:2194]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_5 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi_1, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo_1 = {regroupV0_hi_6[2219:2218], regroupV0_hi_6[2211:2210]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi_1 = {regroupV0_hi_6[2235:2234], regroupV0_hi_6[2227:2226]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_5 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi_1, regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_hi_lo_7 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_5, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_5};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo_1 = {regroupV0_hi_6[2251:2250], regroupV0_hi_6[2243:2242]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi_1 = {regroupV0_hi_6[2267:2266], regroupV0_hi_6[2259:2258]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_5 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi_1, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo_1 = {regroupV0_hi_6[2283:2282], regroupV0_hi_6[2275:2274]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi_1 = {regroupV0_hi_6[2299:2298], regroupV0_hi_6[2291:2290]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_5 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi_1, regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_hi_hi_7 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_5, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_5};
  wire [31:0]        regroupV0_hi_hi_lo_lo_lo_hi_7 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_7, regroupV0_hi_hi_lo_lo_lo_hi_lo_7};
  wire [63:0]        regroupV0_hi_hi_lo_lo_lo_7 = {regroupV0_hi_hi_lo_lo_lo_hi_7, regroupV0_hi_hi_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo_1 = {regroupV0_hi_6[2315:2314], regroupV0_hi_6[2307:2306]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi_1 = {regroupV0_hi_6[2331:2330], regroupV0_hi_6[2323:2322]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_5 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi_1, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo_1 = {regroupV0_hi_6[2347:2346], regroupV0_hi_6[2339:2338]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi_1 = {regroupV0_hi_6[2363:2362], regroupV0_hi_6[2355:2354]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_5 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi_1, regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_lo_lo_7 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_5, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_5};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo_1 = {regroupV0_hi_6[2379:2378], regroupV0_hi_6[2371:2370]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi_1 = {regroupV0_hi_6[2395:2394], regroupV0_hi_6[2387:2386]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_5 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi_1, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo_1 = {regroupV0_hi_6[2411:2410], regroupV0_hi_6[2403:2402]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi_1 = {regroupV0_hi_6[2427:2426], regroupV0_hi_6[2419:2418]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_5 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi_1, regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_lo_hi_7 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_5, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_5};
  wire [31:0]        regroupV0_hi_hi_lo_lo_hi_lo_7 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_7, regroupV0_hi_hi_lo_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo_1 = {regroupV0_hi_6[2443:2442], regroupV0_hi_6[2435:2434]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi_1 = {regroupV0_hi_6[2459:2458], regroupV0_hi_6[2451:2450]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_5 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi_1, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo_1 = {regroupV0_hi_6[2475:2474], regroupV0_hi_6[2467:2466]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi_1 = {regroupV0_hi_6[2491:2490], regroupV0_hi_6[2483:2482]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_5 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi_1, regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_hi_lo_7 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_5, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_5};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo_1 = {regroupV0_hi_6[2507:2506], regroupV0_hi_6[2499:2498]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi_1 = {regroupV0_hi_6[2523:2522], regroupV0_hi_6[2515:2514]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_5 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi_1, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo_1 = {regroupV0_hi_6[2539:2538], regroupV0_hi_6[2531:2530]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi_1 = {regroupV0_hi_6[2555:2554], regroupV0_hi_6[2547:2546]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_5 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi_1, regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_hi_hi_7 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_5, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_5};
  wire [31:0]        regroupV0_hi_hi_lo_lo_hi_hi_7 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_7, regroupV0_hi_hi_lo_lo_hi_hi_lo_7};
  wire [63:0]        regroupV0_hi_hi_lo_lo_hi_7 = {regroupV0_hi_hi_lo_lo_hi_hi_7, regroupV0_hi_hi_lo_lo_hi_lo_7};
  wire [127:0]       regroupV0_hi_hi_lo_lo_7 = {regroupV0_hi_hi_lo_lo_hi_7, regroupV0_hi_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo_1 = {regroupV0_hi_6[2571:2570], regroupV0_hi_6[2563:2562]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi_1 = {regroupV0_hi_6[2587:2586], regroupV0_hi_6[2579:2578]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_5 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi_1, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo_1 = {regroupV0_hi_6[2603:2602], regroupV0_hi_6[2595:2594]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi_1 = {regroupV0_hi_6[2619:2618], regroupV0_hi_6[2611:2610]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_5 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi_1, regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_lo_lo_7 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_5, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_5};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo_1 = {regroupV0_hi_6[2635:2634], regroupV0_hi_6[2627:2626]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi_1 = {regroupV0_hi_6[2651:2650], regroupV0_hi_6[2643:2642]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_5 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi_1, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo_1 = {regroupV0_hi_6[2667:2666], regroupV0_hi_6[2659:2658]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi_1 = {regroupV0_hi_6[2683:2682], regroupV0_hi_6[2675:2674]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_5 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi_1, regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_lo_hi_7 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_5, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_5};
  wire [31:0]        regroupV0_hi_hi_lo_hi_lo_lo_7 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_7, regroupV0_hi_hi_lo_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo_1 = {regroupV0_hi_6[2699:2698], regroupV0_hi_6[2691:2690]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi_1 = {regroupV0_hi_6[2715:2714], regroupV0_hi_6[2707:2706]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_5 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi_1, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo_1 = {regroupV0_hi_6[2731:2730], regroupV0_hi_6[2723:2722]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi_1 = {regroupV0_hi_6[2747:2746], regroupV0_hi_6[2739:2738]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_5 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi_1, regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_hi_lo_7 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_5, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_5};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo_1 = {regroupV0_hi_6[2763:2762], regroupV0_hi_6[2755:2754]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi_1 = {regroupV0_hi_6[2779:2778], regroupV0_hi_6[2771:2770]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_5 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi_1, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo_1 = {regroupV0_hi_6[2795:2794], regroupV0_hi_6[2787:2786]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi_1 = {regroupV0_hi_6[2811:2810], regroupV0_hi_6[2803:2802]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_5 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi_1, regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_hi_hi_7 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_5, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_5};
  wire [31:0]        regroupV0_hi_hi_lo_hi_lo_hi_7 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_7, regroupV0_hi_hi_lo_hi_lo_hi_lo_7};
  wire [63:0]        regroupV0_hi_hi_lo_hi_lo_7 = {regroupV0_hi_hi_lo_hi_lo_hi_7, regroupV0_hi_hi_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo_1 = {regroupV0_hi_6[2827:2826], regroupV0_hi_6[2819:2818]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi_1 = {regroupV0_hi_6[2843:2842], regroupV0_hi_6[2835:2834]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_5 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi_1, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo_1 = {regroupV0_hi_6[2859:2858], regroupV0_hi_6[2851:2850]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi_1 = {regroupV0_hi_6[2875:2874], regroupV0_hi_6[2867:2866]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_5 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi_1, regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_lo_lo_7 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_5, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_5};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo_1 = {regroupV0_hi_6[2891:2890], regroupV0_hi_6[2883:2882]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi_1 = {regroupV0_hi_6[2907:2906], regroupV0_hi_6[2899:2898]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_5 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi_1, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo_1 = {regroupV0_hi_6[2923:2922], regroupV0_hi_6[2915:2914]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi_1 = {regroupV0_hi_6[2939:2938], regroupV0_hi_6[2931:2930]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_5 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi_1, regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_lo_hi_7 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_5, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_5};
  wire [31:0]        regroupV0_hi_hi_lo_hi_hi_lo_7 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_7, regroupV0_hi_hi_lo_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo_1 = {regroupV0_hi_6[2955:2954], regroupV0_hi_6[2947:2946]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi_1 = {regroupV0_hi_6[2971:2970], regroupV0_hi_6[2963:2962]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_5 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi_1, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo_1 = {regroupV0_hi_6[2987:2986], regroupV0_hi_6[2979:2978]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi_1 = {regroupV0_hi_6[3003:3002], regroupV0_hi_6[2995:2994]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_5 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi_1, regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_hi_lo_7 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_5, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_5};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo_1 = {regroupV0_hi_6[3019:3018], regroupV0_hi_6[3011:3010]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi_1 = {regroupV0_hi_6[3035:3034], regroupV0_hi_6[3027:3026]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_5 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi_1, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo_1 = {regroupV0_hi_6[3051:3050], regroupV0_hi_6[3043:3042]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi_1 = {regroupV0_hi_6[3067:3066], regroupV0_hi_6[3059:3058]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_5 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi_1, regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_hi_hi_7 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_5, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_5};
  wire [31:0]        regroupV0_hi_hi_lo_hi_hi_hi_7 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_7, regroupV0_hi_hi_lo_hi_hi_hi_lo_7};
  wire [63:0]        regroupV0_hi_hi_lo_hi_hi_7 = {regroupV0_hi_hi_lo_hi_hi_hi_7, regroupV0_hi_hi_lo_hi_hi_lo_7};
  wire [127:0]       regroupV0_hi_hi_lo_hi_7 = {regroupV0_hi_hi_lo_hi_hi_7, regroupV0_hi_hi_lo_hi_lo_7};
  wire [255:0]       regroupV0_hi_hi_lo_7 = {regroupV0_hi_hi_lo_hi_7, regroupV0_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo_1 = {regroupV0_hi_6[3083:3082], regroupV0_hi_6[3075:3074]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi_1 = {regroupV0_hi_6[3099:3098], regroupV0_hi_6[3091:3090]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_5 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi_1, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo_1 = {regroupV0_hi_6[3115:3114], regroupV0_hi_6[3107:3106]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi_1 = {regroupV0_hi_6[3131:3130], regroupV0_hi_6[3123:3122]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_5 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi_1, regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_lo_lo_7 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_5, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_5};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo_1 = {regroupV0_hi_6[3147:3146], regroupV0_hi_6[3139:3138]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi_1 = {regroupV0_hi_6[3163:3162], regroupV0_hi_6[3155:3154]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_5 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi_1, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo_1 = {regroupV0_hi_6[3179:3178], regroupV0_hi_6[3171:3170]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi_1 = {regroupV0_hi_6[3195:3194], regroupV0_hi_6[3187:3186]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_5 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi_1, regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_lo_hi_7 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_5, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_5};
  wire [31:0]        regroupV0_hi_hi_hi_lo_lo_lo_7 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_7, regroupV0_hi_hi_hi_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo_1 = {regroupV0_hi_6[3211:3210], regroupV0_hi_6[3203:3202]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi_1 = {regroupV0_hi_6[3227:3226], regroupV0_hi_6[3219:3218]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_5 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi_1, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo_1 = {regroupV0_hi_6[3243:3242], regroupV0_hi_6[3235:3234]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi_1 = {regroupV0_hi_6[3259:3258], regroupV0_hi_6[3251:3250]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_5 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi_1, regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_hi_lo_7 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_5, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_5};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo_1 = {regroupV0_hi_6[3275:3274], regroupV0_hi_6[3267:3266]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi_1 = {regroupV0_hi_6[3291:3290], regroupV0_hi_6[3283:3282]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_5 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi_1, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo_1 = {regroupV0_hi_6[3307:3306], regroupV0_hi_6[3299:3298]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi_1 = {regroupV0_hi_6[3323:3322], regroupV0_hi_6[3315:3314]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_5 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_hi_hi_7 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_5, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_5};
  wire [31:0]        regroupV0_hi_hi_hi_lo_lo_hi_7 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_7, regroupV0_hi_hi_hi_lo_lo_hi_lo_7};
  wire [63:0]        regroupV0_hi_hi_hi_lo_lo_7 = {regroupV0_hi_hi_hi_lo_lo_hi_7, regroupV0_hi_hi_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo_1 = {regroupV0_hi_6[3339:3338], regroupV0_hi_6[3331:3330]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi_1 = {regroupV0_hi_6[3355:3354], regroupV0_hi_6[3347:3346]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_5 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi_1, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo_1 = {regroupV0_hi_6[3371:3370], regroupV0_hi_6[3363:3362]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi_1 = {regroupV0_hi_6[3387:3386], regroupV0_hi_6[3379:3378]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_5 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi_1, regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_lo_lo_7 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_5, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_5};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo_1 = {regroupV0_hi_6[3403:3402], regroupV0_hi_6[3395:3394]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi_1 = {regroupV0_hi_6[3419:3418], regroupV0_hi_6[3411:3410]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_5 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi_1, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo_1 = {regroupV0_hi_6[3435:3434], regroupV0_hi_6[3427:3426]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi_1 = {regroupV0_hi_6[3451:3450], regroupV0_hi_6[3443:3442]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_5 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi_1, regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_lo_hi_7 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_5, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_5};
  wire [31:0]        regroupV0_hi_hi_hi_lo_hi_lo_7 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_7, regroupV0_hi_hi_hi_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo_1 = {regroupV0_hi_6[3467:3466], regroupV0_hi_6[3459:3458]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi_1 = {regroupV0_hi_6[3483:3482], regroupV0_hi_6[3475:3474]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_5 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi_1, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo_1 = {regroupV0_hi_6[3499:3498], regroupV0_hi_6[3491:3490]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi_1 = {regroupV0_hi_6[3515:3514], regroupV0_hi_6[3507:3506]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_5 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi_1, regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_hi_lo_7 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_5, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_5};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo_1 = {regroupV0_hi_6[3531:3530], regroupV0_hi_6[3523:3522]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi_1 = {regroupV0_hi_6[3547:3546], regroupV0_hi_6[3539:3538]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_5 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi_1, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo_1 = {regroupV0_hi_6[3563:3562], regroupV0_hi_6[3555:3554]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi_1 = {regroupV0_hi_6[3579:3578], regroupV0_hi_6[3571:3570]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_5 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_hi_hi_7 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_5, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_5};
  wire [31:0]        regroupV0_hi_hi_hi_lo_hi_hi_7 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_7, regroupV0_hi_hi_hi_lo_hi_hi_lo_7};
  wire [63:0]        regroupV0_hi_hi_hi_lo_hi_7 = {regroupV0_hi_hi_hi_lo_hi_hi_7, regroupV0_hi_hi_hi_lo_hi_lo_7};
  wire [127:0]       regroupV0_hi_hi_hi_lo_7 = {regroupV0_hi_hi_hi_lo_hi_7, regroupV0_hi_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo_1 = {regroupV0_hi_6[3595:3594], regroupV0_hi_6[3587:3586]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi_1 = {regroupV0_hi_6[3611:3610], regroupV0_hi_6[3603:3602]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_5 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi_1, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo_1 = {regroupV0_hi_6[3627:3626], regroupV0_hi_6[3619:3618]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi_1 = {regroupV0_hi_6[3643:3642], regroupV0_hi_6[3635:3634]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_5 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi_1, regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_lo_lo_7 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_5, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_5};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo_1 = {regroupV0_hi_6[3659:3658], regroupV0_hi_6[3651:3650]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi_1 = {regroupV0_hi_6[3675:3674], regroupV0_hi_6[3667:3666]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_5 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi_1, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo_1 = {regroupV0_hi_6[3691:3690], regroupV0_hi_6[3683:3682]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi_1 = {regroupV0_hi_6[3707:3706], regroupV0_hi_6[3699:3698]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_5 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi_1, regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_lo_hi_7 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_5, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_5};
  wire [31:0]        regroupV0_hi_hi_hi_hi_lo_lo_7 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_7, regroupV0_hi_hi_hi_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo_1 = {regroupV0_hi_6[3723:3722], regroupV0_hi_6[3715:3714]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi_1 = {regroupV0_hi_6[3739:3738], regroupV0_hi_6[3731:3730]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_5 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi_1, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo_1 = {regroupV0_hi_6[3755:3754], regroupV0_hi_6[3747:3746]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi_1 = {regroupV0_hi_6[3771:3770], regroupV0_hi_6[3763:3762]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_5 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi_1, regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_hi_lo_7 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_5, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_5};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo_1 = {regroupV0_hi_6[3787:3786], regroupV0_hi_6[3779:3778]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi_1 = {regroupV0_hi_6[3803:3802], regroupV0_hi_6[3795:3794]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_5 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi_1, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo_1 = {regroupV0_hi_6[3819:3818], regroupV0_hi_6[3811:3810]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi_1 = {regroupV0_hi_6[3835:3834], regroupV0_hi_6[3827:3826]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_5 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_hi_hi_7 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_5, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_5};
  wire [31:0]        regroupV0_hi_hi_hi_hi_lo_hi_7 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_7, regroupV0_hi_hi_hi_hi_lo_hi_lo_7};
  wire [63:0]        regroupV0_hi_hi_hi_hi_lo_7 = {regroupV0_hi_hi_hi_hi_lo_hi_7, regroupV0_hi_hi_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo_1 = {regroupV0_hi_6[3851:3850], regroupV0_hi_6[3843:3842]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi_1 = {regroupV0_hi_6[3867:3866], regroupV0_hi_6[3859:3858]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_5 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi_1, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo_1 = {regroupV0_hi_6[3883:3882], regroupV0_hi_6[3875:3874]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi_1 = {regroupV0_hi_6[3899:3898], regroupV0_hi_6[3891:3890]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_5 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi_1, regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_lo_lo_7 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_5, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_5};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo_1 = {regroupV0_hi_6[3915:3914], regroupV0_hi_6[3907:3906]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi_1 = {regroupV0_hi_6[3931:3930], regroupV0_hi_6[3923:3922]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_5 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi_1, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo_1 = {regroupV0_hi_6[3947:3946], regroupV0_hi_6[3939:3938]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi_1 = {regroupV0_hi_6[3963:3962], regroupV0_hi_6[3955:3954]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_5 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi_1, regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_lo_hi_7 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_5, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_5};
  wire [31:0]        regroupV0_hi_hi_hi_hi_hi_lo_7 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_7, regroupV0_hi_hi_hi_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo_1 = {regroupV0_hi_6[3979:3978], regroupV0_hi_6[3971:3970]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi_1 = {regroupV0_hi_6[3995:3994], regroupV0_hi_6[3987:3986]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_5 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi_1, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo_1 = {regroupV0_hi_6[4011:4010], regroupV0_hi_6[4003:4002]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi_1 = {regroupV0_hi_6[4027:4026], regroupV0_hi_6[4019:4018]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_5 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi_1, regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_hi_lo_7 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_5, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_5};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo_1 = {regroupV0_hi_6[4043:4042], regroupV0_hi_6[4035:4034]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi_1 = {regroupV0_hi_6[4059:4058], regroupV0_hi_6[4051:4050]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_5 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi_1, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo_1 = {regroupV0_hi_6[4075:4074], regroupV0_hi_6[4067:4066]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi_1 = {regroupV0_hi_6[4091:4090], regroupV0_hi_6[4083:4082]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_5 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_hi_hi_7 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_5, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_5};
  wire [31:0]        regroupV0_hi_hi_hi_hi_hi_hi_7 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_7, regroupV0_hi_hi_hi_hi_hi_hi_lo_7};
  wire [63:0]        regroupV0_hi_hi_hi_hi_hi_7 = {regroupV0_hi_hi_hi_hi_hi_hi_7, regroupV0_hi_hi_hi_hi_hi_lo_7};
  wire [127:0]       regroupV0_hi_hi_hi_hi_7 = {regroupV0_hi_hi_hi_hi_hi_7, regroupV0_hi_hi_hi_hi_lo_7};
  wire [255:0]       regroupV0_hi_hi_hi_7 = {regroupV0_hi_hi_hi_hi_7, regroupV0_hi_hi_hi_lo_7};
  wire [511:0]       regroupV0_hi_hi_7 = {regroupV0_hi_hi_hi_7, regroupV0_hi_hi_lo_7};
  wire [1023:0]      regroupV0_hi_8 = {regroupV0_hi_hi_7, regroupV0_hi_lo_7};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo_2 = {regroupV0_lo_6[13:12], regroupV0_lo_6[5:4]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi_2 = {regroupV0_lo_6[29:28], regroupV0_lo_6[21:20]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_6 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo_2 = {regroupV0_lo_6[45:44], regroupV0_lo_6[37:36]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi_2 = {regroupV0_lo_6[61:60], regroupV0_lo_6[53:52]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_6 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi_2, regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_lo_lo_8 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_6, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo_2 = {regroupV0_lo_6[77:76], regroupV0_lo_6[69:68]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi_2 = {regroupV0_lo_6[93:92], regroupV0_lo_6[85:84]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_6 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi_2, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo_2 = {regroupV0_lo_6[109:108], regroupV0_lo_6[101:100]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi_2 = {regroupV0_lo_6[125:124], regroupV0_lo_6[117:116]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_6 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi_2, regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_lo_hi_8 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_6, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_6};
  wire [31:0]        regroupV0_lo_lo_lo_lo_lo_lo_8 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_8, regroupV0_lo_lo_lo_lo_lo_lo_lo_8};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo_2 = {regroupV0_lo_6[141:140], regroupV0_lo_6[133:132]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi_2 = {regroupV0_lo_6[157:156], regroupV0_lo_6[149:148]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_6 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo_2 = {regroupV0_lo_6[173:172], regroupV0_lo_6[165:164]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi_2 = {regroupV0_lo_6[189:188], regroupV0_lo_6[181:180]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_6 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi_2, regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_hi_lo_8 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_6, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo_2 = {regroupV0_lo_6[205:204], regroupV0_lo_6[197:196]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi_2 = {regroupV0_lo_6[221:220], regroupV0_lo_6[213:212]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_6 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi_2, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo_2 = {regroupV0_lo_6[237:236], regroupV0_lo_6[229:228]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi_2 = {regroupV0_lo_6[253:252], regroupV0_lo_6[245:244]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_6 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi_2, regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_hi_hi_8 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_6, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_6};
  wire [31:0]        regroupV0_lo_lo_lo_lo_lo_hi_8 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_8, regroupV0_lo_lo_lo_lo_lo_hi_lo_8};
  wire [63:0]        regroupV0_lo_lo_lo_lo_lo_8 = {regroupV0_lo_lo_lo_lo_lo_hi_8, regroupV0_lo_lo_lo_lo_lo_lo_8};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo_2 = {regroupV0_lo_6[269:268], regroupV0_lo_6[261:260]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi_2 = {regroupV0_lo_6[285:284], regroupV0_lo_6[277:276]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_6 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo_2 = {regroupV0_lo_6[301:300], regroupV0_lo_6[293:292]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi_2 = {regroupV0_lo_6[317:316], regroupV0_lo_6[309:308]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_6 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi_2, regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_lo_lo_8 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_6, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo_2 = {regroupV0_lo_6[333:332], regroupV0_lo_6[325:324]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi_2 = {regroupV0_lo_6[349:348], regroupV0_lo_6[341:340]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_6 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi_2, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo_2 = {regroupV0_lo_6[365:364], regroupV0_lo_6[357:356]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi_2 = {regroupV0_lo_6[381:380], regroupV0_lo_6[373:372]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_6 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi_2, regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_lo_hi_8 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_6, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_6};
  wire [31:0]        regroupV0_lo_lo_lo_lo_hi_lo_8 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_8, regroupV0_lo_lo_lo_lo_hi_lo_lo_8};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo_2 = {regroupV0_lo_6[397:396], regroupV0_lo_6[389:388]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi_2 = {regroupV0_lo_6[413:412], regroupV0_lo_6[405:404]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_6 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo_2 = {regroupV0_lo_6[429:428], regroupV0_lo_6[421:420]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi_2 = {regroupV0_lo_6[445:444], regroupV0_lo_6[437:436]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_6 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi_2, regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_hi_lo_8 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_6, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo_2 = {regroupV0_lo_6[461:460], regroupV0_lo_6[453:452]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi_2 = {regroupV0_lo_6[477:476], regroupV0_lo_6[469:468]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_6 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi_2, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo_2 = {regroupV0_lo_6[493:492], regroupV0_lo_6[485:484]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi_2 = {regroupV0_lo_6[509:508], regroupV0_lo_6[501:500]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_6 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi_2, regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_hi_hi_8 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_6, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_6};
  wire [31:0]        regroupV0_lo_lo_lo_lo_hi_hi_8 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_8, regroupV0_lo_lo_lo_lo_hi_hi_lo_8};
  wire [63:0]        regroupV0_lo_lo_lo_lo_hi_8 = {regroupV0_lo_lo_lo_lo_hi_hi_8, regroupV0_lo_lo_lo_lo_hi_lo_8};
  wire [127:0]       regroupV0_lo_lo_lo_lo_8 = {regroupV0_lo_lo_lo_lo_hi_8, regroupV0_lo_lo_lo_lo_lo_8};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo_2 = {regroupV0_lo_6[525:524], regroupV0_lo_6[517:516]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi_2 = {regroupV0_lo_6[541:540], regroupV0_lo_6[533:532]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_6 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo_2 = {regroupV0_lo_6[557:556], regroupV0_lo_6[549:548]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi_2 = {regroupV0_lo_6[573:572], regroupV0_lo_6[565:564]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_6 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi_2, regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_lo_lo_8 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_6, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo_2 = {regroupV0_lo_6[589:588], regroupV0_lo_6[581:580]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi_2 = {regroupV0_lo_6[605:604], regroupV0_lo_6[597:596]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_6 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi_2, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo_2 = {regroupV0_lo_6[621:620], regroupV0_lo_6[613:612]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi_2 = {regroupV0_lo_6[637:636], regroupV0_lo_6[629:628]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_6 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi_2, regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_lo_hi_8 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_6, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_6};
  wire [31:0]        regroupV0_lo_lo_lo_hi_lo_lo_8 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_8, regroupV0_lo_lo_lo_hi_lo_lo_lo_8};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo_2 = {regroupV0_lo_6[653:652], regroupV0_lo_6[645:644]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi_2 = {regroupV0_lo_6[669:668], regroupV0_lo_6[661:660]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_6 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi_2, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo_2 = {regroupV0_lo_6[685:684], regroupV0_lo_6[677:676]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi_2 = {regroupV0_lo_6[701:700], regroupV0_lo_6[693:692]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_6 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi_2, regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_hi_lo_8 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_6, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo_2 = {regroupV0_lo_6[717:716], regroupV0_lo_6[709:708]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi_2 = {regroupV0_lo_6[733:732], regroupV0_lo_6[725:724]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_6 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi_2, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo_2 = {regroupV0_lo_6[749:748], regroupV0_lo_6[741:740]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi_2 = {regroupV0_lo_6[765:764], regroupV0_lo_6[757:756]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_6 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi_2, regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_hi_hi_8 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_6, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_6};
  wire [31:0]        regroupV0_lo_lo_lo_hi_lo_hi_8 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_8, regroupV0_lo_lo_lo_hi_lo_hi_lo_8};
  wire [63:0]        regroupV0_lo_lo_lo_hi_lo_8 = {regroupV0_lo_lo_lo_hi_lo_hi_8, regroupV0_lo_lo_lo_hi_lo_lo_8};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo_2 = {regroupV0_lo_6[781:780], regroupV0_lo_6[773:772]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi_2 = {regroupV0_lo_6[797:796], regroupV0_lo_6[789:788]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_6 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo_2 = {regroupV0_lo_6[813:812], regroupV0_lo_6[805:804]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi_2 = {regroupV0_lo_6[829:828], regroupV0_lo_6[821:820]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_6 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi_2, regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_lo_lo_8 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_6, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo_2 = {regroupV0_lo_6[845:844], regroupV0_lo_6[837:836]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi_2 = {regroupV0_lo_6[861:860], regroupV0_lo_6[853:852]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_6 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi_2, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo_2 = {regroupV0_lo_6[877:876], regroupV0_lo_6[869:868]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi_2 = {regroupV0_lo_6[893:892], regroupV0_lo_6[885:884]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_6 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi_2, regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_lo_hi_8 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_6, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_6};
  wire [31:0]        regroupV0_lo_lo_lo_hi_hi_lo_8 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_8, regroupV0_lo_lo_lo_hi_hi_lo_lo_8};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo_2 = {regroupV0_lo_6[909:908], regroupV0_lo_6[901:900]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi_2 = {regroupV0_lo_6[925:924], regroupV0_lo_6[917:916]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_6 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi_2, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo_2 = {regroupV0_lo_6[941:940], regroupV0_lo_6[933:932]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi_2 = {regroupV0_lo_6[957:956], regroupV0_lo_6[949:948]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_6 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi_2, regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_hi_lo_8 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_6, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo_2 = {regroupV0_lo_6[973:972], regroupV0_lo_6[965:964]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi_2 = {regroupV0_lo_6[989:988], regroupV0_lo_6[981:980]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_6 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi_2, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo_2 = {regroupV0_lo_6[1005:1004], regroupV0_lo_6[997:996]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi_2 = {regroupV0_lo_6[1021:1020], regroupV0_lo_6[1013:1012]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_6 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi_2, regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_hi_hi_8 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_6, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_6};
  wire [31:0]        regroupV0_lo_lo_lo_hi_hi_hi_8 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_8, regroupV0_lo_lo_lo_hi_hi_hi_lo_8};
  wire [63:0]        regroupV0_lo_lo_lo_hi_hi_8 = {regroupV0_lo_lo_lo_hi_hi_hi_8, regroupV0_lo_lo_lo_hi_hi_lo_8};
  wire [127:0]       regroupV0_lo_lo_lo_hi_8 = {regroupV0_lo_lo_lo_hi_hi_8, regroupV0_lo_lo_lo_hi_lo_8};
  wire [255:0]       regroupV0_lo_lo_lo_8 = {regroupV0_lo_lo_lo_hi_8, regroupV0_lo_lo_lo_lo_8};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo_2 = {regroupV0_lo_6[1037:1036], regroupV0_lo_6[1029:1028]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi_2 = {regroupV0_lo_6[1053:1052], regroupV0_lo_6[1045:1044]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_6 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi_2, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo_2 = {regroupV0_lo_6[1069:1068], regroupV0_lo_6[1061:1060]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi_2 = {regroupV0_lo_6[1085:1084], regroupV0_lo_6[1077:1076]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_6 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi_2, regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_lo_lo_8 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_6, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo_2 = {regroupV0_lo_6[1101:1100], regroupV0_lo_6[1093:1092]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi_2 = {regroupV0_lo_6[1117:1116], regroupV0_lo_6[1109:1108]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_6 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi_2, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo_2 = {regroupV0_lo_6[1133:1132], regroupV0_lo_6[1125:1124]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi_2 = {regroupV0_lo_6[1149:1148], regroupV0_lo_6[1141:1140]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_6 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi_2, regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_lo_hi_8 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_6, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_6};
  wire [31:0]        regroupV0_lo_lo_hi_lo_lo_lo_8 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_8, regroupV0_lo_lo_hi_lo_lo_lo_lo_8};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo_2 = {regroupV0_lo_6[1165:1164], regroupV0_lo_6[1157:1156]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi_2 = {regroupV0_lo_6[1181:1180], regroupV0_lo_6[1173:1172]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_6 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi_2, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo_2 = {regroupV0_lo_6[1197:1196], regroupV0_lo_6[1189:1188]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi_2 = {regroupV0_lo_6[1213:1212], regroupV0_lo_6[1205:1204]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_6 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi_2, regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_hi_lo_8 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_6, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo_2 = {regroupV0_lo_6[1229:1228], regroupV0_lo_6[1221:1220]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi_2 = {regroupV0_lo_6[1245:1244], regroupV0_lo_6[1237:1236]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_6 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi_2, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo_2 = {regroupV0_lo_6[1261:1260], regroupV0_lo_6[1253:1252]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi_2 = {regroupV0_lo_6[1277:1276], regroupV0_lo_6[1269:1268]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_6 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi_2, regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_hi_hi_8 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_6, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_6};
  wire [31:0]        regroupV0_lo_lo_hi_lo_lo_hi_8 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_8, regroupV0_lo_lo_hi_lo_lo_hi_lo_8};
  wire [63:0]        regroupV0_lo_lo_hi_lo_lo_8 = {regroupV0_lo_lo_hi_lo_lo_hi_8, regroupV0_lo_lo_hi_lo_lo_lo_8};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo_2 = {regroupV0_lo_6[1293:1292], regroupV0_lo_6[1285:1284]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi_2 = {regroupV0_lo_6[1309:1308], regroupV0_lo_6[1301:1300]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_6 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi_2, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo_2 = {regroupV0_lo_6[1325:1324], regroupV0_lo_6[1317:1316]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi_2 = {regroupV0_lo_6[1341:1340], regroupV0_lo_6[1333:1332]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_6 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi_2, regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_lo_lo_8 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_6, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo_2 = {regroupV0_lo_6[1357:1356], regroupV0_lo_6[1349:1348]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi_2 = {regroupV0_lo_6[1373:1372], regroupV0_lo_6[1365:1364]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_6 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi_2, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo_2 = {regroupV0_lo_6[1389:1388], regroupV0_lo_6[1381:1380]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi_2 = {regroupV0_lo_6[1405:1404], regroupV0_lo_6[1397:1396]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_6 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi_2, regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_lo_hi_8 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_6, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_6};
  wire [31:0]        regroupV0_lo_lo_hi_lo_hi_lo_8 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_8, regroupV0_lo_lo_hi_lo_hi_lo_lo_8};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo_2 = {regroupV0_lo_6[1421:1420], regroupV0_lo_6[1413:1412]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi_2 = {regroupV0_lo_6[1437:1436], regroupV0_lo_6[1429:1428]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_6 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi_2, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo_2 = {regroupV0_lo_6[1453:1452], regroupV0_lo_6[1445:1444]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi_2 = {regroupV0_lo_6[1469:1468], regroupV0_lo_6[1461:1460]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_6 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi_2, regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_hi_lo_8 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_6, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo_2 = {regroupV0_lo_6[1485:1484], regroupV0_lo_6[1477:1476]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi_2 = {regroupV0_lo_6[1501:1500], regroupV0_lo_6[1493:1492]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_6 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi_2, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo_2 = {regroupV0_lo_6[1517:1516], regroupV0_lo_6[1509:1508]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi_2 = {regroupV0_lo_6[1533:1532], regroupV0_lo_6[1525:1524]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_6 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi_2, regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_hi_hi_8 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_6, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_6};
  wire [31:0]        regroupV0_lo_lo_hi_lo_hi_hi_8 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_8, regroupV0_lo_lo_hi_lo_hi_hi_lo_8};
  wire [63:0]        regroupV0_lo_lo_hi_lo_hi_8 = {regroupV0_lo_lo_hi_lo_hi_hi_8, regroupV0_lo_lo_hi_lo_hi_lo_8};
  wire [127:0]       regroupV0_lo_lo_hi_lo_8 = {regroupV0_lo_lo_hi_lo_hi_8, regroupV0_lo_lo_hi_lo_lo_8};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo_2 = {regroupV0_lo_6[1549:1548], regroupV0_lo_6[1541:1540]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi_2 = {regroupV0_lo_6[1565:1564], regroupV0_lo_6[1557:1556]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_6 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi_2, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo_2 = {regroupV0_lo_6[1581:1580], regroupV0_lo_6[1573:1572]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi_2 = {regroupV0_lo_6[1597:1596], regroupV0_lo_6[1589:1588]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_6 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi_2, regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_lo_lo_8 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_6, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo_2 = {regroupV0_lo_6[1613:1612], regroupV0_lo_6[1605:1604]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi_2 = {regroupV0_lo_6[1629:1628], regroupV0_lo_6[1621:1620]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_6 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi_2, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo_2 = {regroupV0_lo_6[1645:1644], regroupV0_lo_6[1637:1636]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi_2 = {regroupV0_lo_6[1661:1660], regroupV0_lo_6[1653:1652]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_6 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi_2, regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_lo_hi_8 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_6, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_6};
  wire [31:0]        regroupV0_lo_lo_hi_hi_lo_lo_8 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_8, regroupV0_lo_lo_hi_hi_lo_lo_lo_8};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo_2 = {regroupV0_lo_6[1677:1676], regroupV0_lo_6[1669:1668]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi_2 = {regroupV0_lo_6[1693:1692], regroupV0_lo_6[1685:1684]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_6 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi_2, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo_2 = {regroupV0_lo_6[1709:1708], regroupV0_lo_6[1701:1700]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi_2 = {regroupV0_lo_6[1725:1724], regroupV0_lo_6[1717:1716]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_6 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi_2, regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_hi_lo_8 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_6, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo_2 = {regroupV0_lo_6[1741:1740], regroupV0_lo_6[1733:1732]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi_2 = {regroupV0_lo_6[1757:1756], regroupV0_lo_6[1749:1748]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_6 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi_2, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo_2 = {regroupV0_lo_6[1773:1772], regroupV0_lo_6[1765:1764]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi_2 = {regroupV0_lo_6[1789:1788], regroupV0_lo_6[1781:1780]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_6 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi_2, regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_hi_hi_8 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_6, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_6};
  wire [31:0]        regroupV0_lo_lo_hi_hi_lo_hi_8 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_8, regroupV0_lo_lo_hi_hi_lo_hi_lo_8};
  wire [63:0]        regroupV0_lo_lo_hi_hi_lo_8 = {regroupV0_lo_lo_hi_hi_lo_hi_8, regroupV0_lo_lo_hi_hi_lo_lo_8};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo_2 = {regroupV0_lo_6[1805:1804], regroupV0_lo_6[1797:1796]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi_2 = {regroupV0_lo_6[1821:1820], regroupV0_lo_6[1813:1812]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_6 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi_2, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo_2 = {regroupV0_lo_6[1837:1836], regroupV0_lo_6[1829:1828]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi_2 = {regroupV0_lo_6[1853:1852], regroupV0_lo_6[1845:1844]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_6 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi_2, regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_lo_lo_8 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_6, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo_2 = {regroupV0_lo_6[1869:1868], regroupV0_lo_6[1861:1860]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi_2 = {regroupV0_lo_6[1885:1884], regroupV0_lo_6[1877:1876]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_6 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi_2, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo_2 = {regroupV0_lo_6[1901:1900], regroupV0_lo_6[1893:1892]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi_2 = {regroupV0_lo_6[1917:1916], regroupV0_lo_6[1909:1908]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_6 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi_2, regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_lo_hi_8 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_6, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_6};
  wire [31:0]        regroupV0_lo_lo_hi_hi_hi_lo_8 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_8, regroupV0_lo_lo_hi_hi_hi_lo_lo_8};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo_2 = {regroupV0_lo_6[1933:1932], regroupV0_lo_6[1925:1924]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi_2 = {regroupV0_lo_6[1949:1948], regroupV0_lo_6[1941:1940]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_6 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi_2, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo_2 = {regroupV0_lo_6[1965:1964], regroupV0_lo_6[1957:1956]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi_2 = {regroupV0_lo_6[1981:1980], regroupV0_lo_6[1973:1972]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_6 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi_2, regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_hi_lo_8 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_6, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo_2 = {regroupV0_lo_6[1997:1996], regroupV0_lo_6[1989:1988]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi_2 = {regroupV0_lo_6[2013:2012], regroupV0_lo_6[2005:2004]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_6 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi_2, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo_2 = {regroupV0_lo_6[2029:2028], regroupV0_lo_6[2021:2020]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi_2 = {regroupV0_lo_6[2045:2044], regroupV0_lo_6[2037:2036]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_6 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi_2, regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_hi_hi_8 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_6, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_6};
  wire [31:0]        regroupV0_lo_lo_hi_hi_hi_hi_8 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_8, regroupV0_lo_lo_hi_hi_hi_hi_lo_8};
  wire [63:0]        regroupV0_lo_lo_hi_hi_hi_8 = {regroupV0_lo_lo_hi_hi_hi_hi_8, regroupV0_lo_lo_hi_hi_hi_lo_8};
  wire [127:0]       regroupV0_lo_lo_hi_hi_8 = {regroupV0_lo_lo_hi_hi_hi_8, regroupV0_lo_lo_hi_hi_lo_8};
  wire [255:0]       regroupV0_lo_lo_hi_8 = {regroupV0_lo_lo_hi_hi_8, regroupV0_lo_lo_hi_lo_8};
  wire [511:0]       regroupV0_lo_lo_8 = {regroupV0_lo_lo_hi_8, regroupV0_lo_lo_lo_8};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo_2 = {regroupV0_lo_6[2061:2060], regroupV0_lo_6[2053:2052]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi_2 = {regroupV0_lo_6[2077:2076], regroupV0_lo_6[2069:2068]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_6 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi_2, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo_2 = {regroupV0_lo_6[2093:2092], regroupV0_lo_6[2085:2084]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi_2 = {regroupV0_lo_6[2109:2108], regroupV0_lo_6[2101:2100]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_6 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi_2, regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_lo_lo_8 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_6, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo_2 = {regroupV0_lo_6[2125:2124], regroupV0_lo_6[2117:2116]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi_2 = {regroupV0_lo_6[2141:2140], regroupV0_lo_6[2133:2132]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_6 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi_2, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo_2 = {regroupV0_lo_6[2157:2156], regroupV0_lo_6[2149:2148]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi_2 = {regroupV0_lo_6[2173:2172], regroupV0_lo_6[2165:2164]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_6 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi_2, regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_lo_hi_8 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_6, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_6};
  wire [31:0]        regroupV0_lo_hi_lo_lo_lo_lo_8 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_8, regroupV0_lo_hi_lo_lo_lo_lo_lo_8};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo_2 = {regroupV0_lo_6[2189:2188], regroupV0_lo_6[2181:2180]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi_2 = {regroupV0_lo_6[2205:2204], regroupV0_lo_6[2197:2196]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_6 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi_2, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo_2 = {regroupV0_lo_6[2221:2220], regroupV0_lo_6[2213:2212]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi_2 = {regroupV0_lo_6[2237:2236], regroupV0_lo_6[2229:2228]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_6 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi_2, regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_hi_lo_8 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_6, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo_2 = {regroupV0_lo_6[2253:2252], regroupV0_lo_6[2245:2244]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi_2 = {regroupV0_lo_6[2269:2268], regroupV0_lo_6[2261:2260]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_6 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi_2, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo_2 = {regroupV0_lo_6[2285:2284], regroupV0_lo_6[2277:2276]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi_2 = {regroupV0_lo_6[2301:2300], regroupV0_lo_6[2293:2292]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_6 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi_2, regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_hi_hi_8 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_6, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_6};
  wire [31:0]        regroupV0_lo_hi_lo_lo_lo_hi_8 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_8, regroupV0_lo_hi_lo_lo_lo_hi_lo_8};
  wire [63:0]        regroupV0_lo_hi_lo_lo_lo_8 = {regroupV0_lo_hi_lo_lo_lo_hi_8, regroupV0_lo_hi_lo_lo_lo_lo_8};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo_2 = {regroupV0_lo_6[2317:2316], regroupV0_lo_6[2309:2308]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi_2 = {regroupV0_lo_6[2333:2332], regroupV0_lo_6[2325:2324]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_6 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi_2, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo_2 = {regroupV0_lo_6[2349:2348], regroupV0_lo_6[2341:2340]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi_2 = {regroupV0_lo_6[2365:2364], regroupV0_lo_6[2357:2356]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_6 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi_2, regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_lo_lo_8 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_6, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo_2 = {regroupV0_lo_6[2381:2380], regroupV0_lo_6[2373:2372]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi_2 = {regroupV0_lo_6[2397:2396], regroupV0_lo_6[2389:2388]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_6 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi_2, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo_2 = {regroupV0_lo_6[2413:2412], regroupV0_lo_6[2405:2404]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi_2 = {regroupV0_lo_6[2429:2428], regroupV0_lo_6[2421:2420]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_6 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi_2, regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_lo_hi_8 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_6, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_6};
  wire [31:0]        regroupV0_lo_hi_lo_lo_hi_lo_8 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_8, regroupV0_lo_hi_lo_lo_hi_lo_lo_8};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo_2 = {regroupV0_lo_6[2445:2444], regroupV0_lo_6[2437:2436]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi_2 = {regroupV0_lo_6[2461:2460], regroupV0_lo_6[2453:2452]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_6 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi_2, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo_2 = {regroupV0_lo_6[2477:2476], regroupV0_lo_6[2469:2468]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi_2 = {regroupV0_lo_6[2493:2492], regroupV0_lo_6[2485:2484]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_6 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi_2, regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_hi_lo_8 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_6, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo_2 = {regroupV0_lo_6[2509:2508], regroupV0_lo_6[2501:2500]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi_2 = {regroupV0_lo_6[2525:2524], regroupV0_lo_6[2517:2516]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_6 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi_2, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo_2 = {regroupV0_lo_6[2541:2540], regroupV0_lo_6[2533:2532]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi_2 = {regroupV0_lo_6[2557:2556], regroupV0_lo_6[2549:2548]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_6 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi_2, regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_hi_hi_8 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_6, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_6};
  wire [31:0]        regroupV0_lo_hi_lo_lo_hi_hi_8 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_8, regroupV0_lo_hi_lo_lo_hi_hi_lo_8};
  wire [63:0]        regroupV0_lo_hi_lo_lo_hi_8 = {regroupV0_lo_hi_lo_lo_hi_hi_8, regroupV0_lo_hi_lo_lo_hi_lo_8};
  wire [127:0]       regroupV0_lo_hi_lo_lo_8 = {regroupV0_lo_hi_lo_lo_hi_8, regroupV0_lo_hi_lo_lo_lo_8};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo_2 = {regroupV0_lo_6[2573:2572], regroupV0_lo_6[2565:2564]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi_2 = {regroupV0_lo_6[2589:2588], regroupV0_lo_6[2581:2580]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_6 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi_2, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo_2 = {regroupV0_lo_6[2605:2604], regroupV0_lo_6[2597:2596]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi_2 = {regroupV0_lo_6[2621:2620], regroupV0_lo_6[2613:2612]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_6 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi_2, regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_lo_lo_8 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_6, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo_2 = {regroupV0_lo_6[2637:2636], regroupV0_lo_6[2629:2628]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi_2 = {regroupV0_lo_6[2653:2652], regroupV0_lo_6[2645:2644]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_6 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi_2, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo_2 = {regroupV0_lo_6[2669:2668], regroupV0_lo_6[2661:2660]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi_2 = {regroupV0_lo_6[2685:2684], regroupV0_lo_6[2677:2676]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_6 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi_2, regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_lo_hi_8 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_6, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_6};
  wire [31:0]        regroupV0_lo_hi_lo_hi_lo_lo_8 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_8, regroupV0_lo_hi_lo_hi_lo_lo_lo_8};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo_2 = {regroupV0_lo_6[2701:2700], regroupV0_lo_6[2693:2692]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi_2 = {regroupV0_lo_6[2717:2716], regroupV0_lo_6[2709:2708]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_6 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi_2, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo_2 = {regroupV0_lo_6[2733:2732], regroupV0_lo_6[2725:2724]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi_2 = {regroupV0_lo_6[2749:2748], regroupV0_lo_6[2741:2740]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_6 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi_2, regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_hi_lo_8 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_6, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo_2 = {regroupV0_lo_6[2765:2764], regroupV0_lo_6[2757:2756]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi_2 = {regroupV0_lo_6[2781:2780], regroupV0_lo_6[2773:2772]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_6 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi_2, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo_2 = {regroupV0_lo_6[2797:2796], regroupV0_lo_6[2789:2788]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi_2 = {regroupV0_lo_6[2813:2812], regroupV0_lo_6[2805:2804]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_6 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi_2, regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_hi_hi_8 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_6, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_6};
  wire [31:0]        regroupV0_lo_hi_lo_hi_lo_hi_8 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_8, regroupV0_lo_hi_lo_hi_lo_hi_lo_8};
  wire [63:0]        regroupV0_lo_hi_lo_hi_lo_8 = {regroupV0_lo_hi_lo_hi_lo_hi_8, regroupV0_lo_hi_lo_hi_lo_lo_8};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo_2 = {regroupV0_lo_6[2829:2828], regroupV0_lo_6[2821:2820]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi_2 = {regroupV0_lo_6[2845:2844], regroupV0_lo_6[2837:2836]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_6 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi_2, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo_2 = {regroupV0_lo_6[2861:2860], regroupV0_lo_6[2853:2852]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi_2 = {regroupV0_lo_6[2877:2876], regroupV0_lo_6[2869:2868]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_6 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi_2, regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_lo_lo_8 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_6, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo_2 = {regroupV0_lo_6[2893:2892], regroupV0_lo_6[2885:2884]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi_2 = {regroupV0_lo_6[2909:2908], regroupV0_lo_6[2901:2900]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_6 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi_2, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo_2 = {regroupV0_lo_6[2925:2924], regroupV0_lo_6[2917:2916]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi_2 = {regroupV0_lo_6[2941:2940], regroupV0_lo_6[2933:2932]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_6 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi_2, regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_lo_hi_8 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_6, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_6};
  wire [31:0]        regroupV0_lo_hi_lo_hi_hi_lo_8 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_8, regroupV0_lo_hi_lo_hi_hi_lo_lo_8};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo_2 = {regroupV0_lo_6[2957:2956], regroupV0_lo_6[2949:2948]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi_2 = {regroupV0_lo_6[2973:2972], regroupV0_lo_6[2965:2964]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_6 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi_2, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo_2 = {regroupV0_lo_6[2989:2988], regroupV0_lo_6[2981:2980]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi_2 = {regroupV0_lo_6[3005:3004], regroupV0_lo_6[2997:2996]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_6 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi_2, regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_hi_lo_8 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_6, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo_2 = {regroupV0_lo_6[3021:3020], regroupV0_lo_6[3013:3012]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi_2 = {regroupV0_lo_6[3037:3036], regroupV0_lo_6[3029:3028]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_6 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi_2, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo_2 = {regroupV0_lo_6[3053:3052], regroupV0_lo_6[3045:3044]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi_2 = {regroupV0_lo_6[3069:3068], regroupV0_lo_6[3061:3060]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_6 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi_2, regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_hi_hi_8 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_6, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_6};
  wire [31:0]        regroupV0_lo_hi_lo_hi_hi_hi_8 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_8, regroupV0_lo_hi_lo_hi_hi_hi_lo_8};
  wire [63:0]        regroupV0_lo_hi_lo_hi_hi_8 = {regroupV0_lo_hi_lo_hi_hi_hi_8, regroupV0_lo_hi_lo_hi_hi_lo_8};
  wire [127:0]       regroupV0_lo_hi_lo_hi_8 = {regroupV0_lo_hi_lo_hi_hi_8, regroupV0_lo_hi_lo_hi_lo_8};
  wire [255:0]       regroupV0_lo_hi_lo_8 = {regroupV0_lo_hi_lo_hi_8, regroupV0_lo_hi_lo_lo_8};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo_2 = {regroupV0_lo_6[3085:3084], regroupV0_lo_6[3077:3076]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi_2 = {regroupV0_lo_6[3101:3100], regroupV0_lo_6[3093:3092]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_6 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi_2, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo_2 = {regroupV0_lo_6[3117:3116], regroupV0_lo_6[3109:3108]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi_2 = {regroupV0_lo_6[3133:3132], regroupV0_lo_6[3125:3124]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_6 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi_2, regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_lo_lo_8 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_6, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo_2 = {regroupV0_lo_6[3149:3148], regroupV0_lo_6[3141:3140]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi_2 = {regroupV0_lo_6[3165:3164], regroupV0_lo_6[3157:3156]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_6 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi_2, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo_2 = {regroupV0_lo_6[3181:3180], regroupV0_lo_6[3173:3172]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi_2 = {regroupV0_lo_6[3197:3196], regroupV0_lo_6[3189:3188]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_6 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi_2, regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_lo_hi_8 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_6, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_6};
  wire [31:0]        regroupV0_lo_hi_hi_lo_lo_lo_8 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_8, regroupV0_lo_hi_hi_lo_lo_lo_lo_8};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo_2 = {regroupV0_lo_6[3213:3212], regroupV0_lo_6[3205:3204]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi_2 = {regroupV0_lo_6[3229:3228], regroupV0_lo_6[3221:3220]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_6 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi_2, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo_2 = {regroupV0_lo_6[3245:3244], regroupV0_lo_6[3237:3236]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi_2 = {regroupV0_lo_6[3261:3260], regroupV0_lo_6[3253:3252]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_6 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi_2, regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_hi_lo_8 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_6, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo_2 = {regroupV0_lo_6[3277:3276], regroupV0_lo_6[3269:3268]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi_2 = {regroupV0_lo_6[3293:3292], regroupV0_lo_6[3285:3284]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_6 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi_2, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo_2 = {regroupV0_lo_6[3309:3308], regroupV0_lo_6[3301:3300]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi_2 = {regroupV0_lo_6[3325:3324], regroupV0_lo_6[3317:3316]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_6 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi_2, regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_hi_hi_8 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_6, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_6};
  wire [31:0]        regroupV0_lo_hi_hi_lo_lo_hi_8 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_8, regroupV0_lo_hi_hi_lo_lo_hi_lo_8};
  wire [63:0]        regroupV0_lo_hi_hi_lo_lo_8 = {regroupV0_lo_hi_hi_lo_lo_hi_8, regroupV0_lo_hi_hi_lo_lo_lo_8};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo_2 = {regroupV0_lo_6[3341:3340], regroupV0_lo_6[3333:3332]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi_2 = {regroupV0_lo_6[3357:3356], regroupV0_lo_6[3349:3348]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_6 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi_2, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo_2 = {regroupV0_lo_6[3373:3372], regroupV0_lo_6[3365:3364]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi_2 = {regroupV0_lo_6[3389:3388], regroupV0_lo_6[3381:3380]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_6 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi_2, regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_lo_lo_8 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_6, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo_2 = {regroupV0_lo_6[3405:3404], regroupV0_lo_6[3397:3396]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi_2 = {regroupV0_lo_6[3421:3420], regroupV0_lo_6[3413:3412]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_6 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi_2, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo_2 = {regroupV0_lo_6[3437:3436], regroupV0_lo_6[3429:3428]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi_2 = {regroupV0_lo_6[3453:3452], regroupV0_lo_6[3445:3444]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_6 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi_2, regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_lo_hi_8 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_6, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_6};
  wire [31:0]        regroupV0_lo_hi_hi_lo_hi_lo_8 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_8, regroupV0_lo_hi_hi_lo_hi_lo_lo_8};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo_2 = {regroupV0_lo_6[3469:3468], regroupV0_lo_6[3461:3460]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi_2 = {regroupV0_lo_6[3485:3484], regroupV0_lo_6[3477:3476]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_6 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi_2, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo_2 = {regroupV0_lo_6[3501:3500], regroupV0_lo_6[3493:3492]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi_2 = {regroupV0_lo_6[3517:3516], regroupV0_lo_6[3509:3508]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_6 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi_2, regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_hi_lo_8 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_6, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo_2 = {regroupV0_lo_6[3533:3532], regroupV0_lo_6[3525:3524]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi_2 = {regroupV0_lo_6[3549:3548], regroupV0_lo_6[3541:3540]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_6 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi_2, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo_2 = {regroupV0_lo_6[3565:3564], regroupV0_lo_6[3557:3556]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi_2 = {regroupV0_lo_6[3581:3580], regroupV0_lo_6[3573:3572]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_6 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi_2, regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_hi_hi_8 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_6, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_6};
  wire [31:0]        regroupV0_lo_hi_hi_lo_hi_hi_8 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_8, regroupV0_lo_hi_hi_lo_hi_hi_lo_8};
  wire [63:0]        regroupV0_lo_hi_hi_lo_hi_8 = {regroupV0_lo_hi_hi_lo_hi_hi_8, regroupV0_lo_hi_hi_lo_hi_lo_8};
  wire [127:0]       regroupV0_lo_hi_hi_lo_8 = {regroupV0_lo_hi_hi_lo_hi_8, regroupV0_lo_hi_hi_lo_lo_8};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo_2 = {regroupV0_lo_6[3597:3596], regroupV0_lo_6[3589:3588]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi_2 = {regroupV0_lo_6[3613:3612], regroupV0_lo_6[3605:3604]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_6 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi_2, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo_2 = {regroupV0_lo_6[3629:3628], regroupV0_lo_6[3621:3620]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi_2 = {regroupV0_lo_6[3645:3644], regroupV0_lo_6[3637:3636]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_6 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi_2, regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_lo_lo_8 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_6, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo_2 = {regroupV0_lo_6[3661:3660], regroupV0_lo_6[3653:3652]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi_2 = {regroupV0_lo_6[3677:3676], regroupV0_lo_6[3669:3668]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_6 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi_2, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo_2 = {regroupV0_lo_6[3693:3692], regroupV0_lo_6[3685:3684]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi_2 = {regroupV0_lo_6[3709:3708], regroupV0_lo_6[3701:3700]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_6 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi_2, regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_lo_hi_8 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_6, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_6};
  wire [31:0]        regroupV0_lo_hi_hi_hi_lo_lo_8 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_8, regroupV0_lo_hi_hi_hi_lo_lo_lo_8};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo_2 = {regroupV0_lo_6[3725:3724], regroupV0_lo_6[3717:3716]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi_2 = {regroupV0_lo_6[3741:3740], regroupV0_lo_6[3733:3732]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_6 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi_2, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo_2 = {regroupV0_lo_6[3757:3756], regroupV0_lo_6[3749:3748]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi_2 = {regroupV0_lo_6[3773:3772], regroupV0_lo_6[3765:3764]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_6 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi_2, regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_hi_lo_8 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_6, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo_2 = {regroupV0_lo_6[3789:3788], regroupV0_lo_6[3781:3780]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi_2 = {regroupV0_lo_6[3805:3804], regroupV0_lo_6[3797:3796]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_6 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi_2, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo_2 = {regroupV0_lo_6[3821:3820], regroupV0_lo_6[3813:3812]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi_2 = {regroupV0_lo_6[3837:3836], regroupV0_lo_6[3829:3828]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_6 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi_2, regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_hi_hi_8 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_6, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_6};
  wire [31:0]        regroupV0_lo_hi_hi_hi_lo_hi_8 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_8, regroupV0_lo_hi_hi_hi_lo_hi_lo_8};
  wire [63:0]        regroupV0_lo_hi_hi_hi_lo_8 = {regroupV0_lo_hi_hi_hi_lo_hi_8, regroupV0_lo_hi_hi_hi_lo_lo_8};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo_2 = {regroupV0_lo_6[3853:3852], regroupV0_lo_6[3845:3844]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi_2 = {regroupV0_lo_6[3869:3868], regroupV0_lo_6[3861:3860]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_6 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi_2, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo_2 = {regroupV0_lo_6[3885:3884], regroupV0_lo_6[3877:3876]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi_2 = {regroupV0_lo_6[3901:3900], regroupV0_lo_6[3893:3892]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_6 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi_2, regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_lo_lo_8 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_6, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo_2 = {regroupV0_lo_6[3917:3916], regroupV0_lo_6[3909:3908]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi_2 = {regroupV0_lo_6[3933:3932], regroupV0_lo_6[3925:3924]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_6 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi_2, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo_2 = {regroupV0_lo_6[3949:3948], regroupV0_lo_6[3941:3940]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi_2 = {regroupV0_lo_6[3965:3964], regroupV0_lo_6[3957:3956]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_6 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi_2, regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_lo_hi_8 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_6, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_6};
  wire [31:0]        regroupV0_lo_hi_hi_hi_hi_lo_8 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_8, regroupV0_lo_hi_hi_hi_hi_lo_lo_8};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo_2 = {regroupV0_lo_6[3981:3980], regroupV0_lo_6[3973:3972]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi_2 = {regroupV0_lo_6[3997:3996], regroupV0_lo_6[3989:3988]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_6 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi_2, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo_2 = {regroupV0_lo_6[4013:4012], regroupV0_lo_6[4005:4004]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi_2 = {regroupV0_lo_6[4029:4028], regroupV0_lo_6[4021:4020]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_6 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi_2, regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_hi_lo_8 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_6, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo_2 = {regroupV0_lo_6[4045:4044], regroupV0_lo_6[4037:4036]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi_2 = {regroupV0_lo_6[4061:4060], regroupV0_lo_6[4053:4052]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_6 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi_2, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo_2 = {regroupV0_lo_6[4077:4076], regroupV0_lo_6[4069:4068]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi_2 = {regroupV0_lo_6[4093:4092], regroupV0_lo_6[4085:4084]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_6 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi_2, regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_hi_hi_8 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_6, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_6};
  wire [31:0]        regroupV0_lo_hi_hi_hi_hi_hi_8 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_8, regroupV0_lo_hi_hi_hi_hi_hi_lo_8};
  wire [63:0]        regroupV0_lo_hi_hi_hi_hi_8 = {regroupV0_lo_hi_hi_hi_hi_hi_8, regroupV0_lo_hi_hi_hi_hi_lo_8};
  wire [127:0]       regroupV0_lo_hi_hi_hi_8 = {regroupV0_lo_hi_hi_hi_hi_8, regroupV0_lo_hi_hi_hi_lo_8};
  wire [255:0]       regroupV0_lo_hi_hi_8 = {regroupV0_lo_hi_hi_hi_8, regroupV0_lo_hi_hi_lo_8};
  wire [511:0]       regroupV0_lo_hi_8 = {regroupV0_lo_hi_hi_8, regroupV0_lo_hi_lo_8};
  wire [1023:0]      regroupV0_lo_9 = {regroupV0_lo_hi_8, regroupV0_lo_lo_8};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo_2 = {regroupV0_hi_6[13:12], regroupV0_hi_6[5:4]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi_2 = {regroupV0_hi_6[29:28], regroupV0_hi_6[21:20]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_6 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo_2 = {regroupV0_hi_6[45:44], regroupV0_hi_6[37:36]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi_2 = {regroupV0_hi_6[61:60], regroupV0_hi_6[53:52]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_6 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi_2, regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_lo_lo_8 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_6, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo_2 = {regroupV0_hi_6[77:76], regroupV0_hi_6[69:68]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi_2 = {regroupV0_hi_6[93:92], regroupV0_hi_6[85:84]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_6 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi_2, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo_2 = {regroupV0_hi_6[109:108], regroupV0_hi_6[101:100]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi_2 = {regroupV0_hi_6[125:124], regroupV0_hi_6[117:116]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_6 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi_2, regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_lo_hi_8 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_6, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_6};
  wire [31:0]        regroupV0_hi_lo_lo_lo_lo_lo_8 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_8, regroupV0_hi_lo_lo_lo_lo_lo_lo_8};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo_2 = {regroupV0_hi_6[141:140], regroupV0_hi_6[133:132]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi_2 = {regroupV0_hi_6[157:156], regroupV0_hi_6[149:148]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_6 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo_2 = {regroupV0_hi_6[173:172], regroupV0_hi_6[165:164]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi_2 = {regroupV0_hi_6[189:188], regroupV0_hi_6[181:180]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_6 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi_2, regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_hi_lo_8 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_6, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo_2 = {regroupV0_hi_6[205:204], regroupV0_hi_6[197:196]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi_2 = {regroupV0_hi_6[221:220], regroupV0_hi_6[213:212]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_6 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi_2, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo_2 = {regroupV0_hi_6[237:236], regroupV0_hi_6[229:228]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi_2 = {regroupV0_hi_6[253:252], regroupV0_hi_6[245:244]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_6 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi_2, regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_hi_hi_8 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_6, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_6};
  wire [31:0]        regroupV0_hi_lo_lo_lo_lo_hi_8 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_8, regroupV0_hi_lo_lo_lo_lo_hi_lo_8};
  wire [63:0]        regroupV0_hi_lo_lo_lo_lo_8 = {regroupV0_hi_lo_lo_lo_lo_hi_8, regroupV0_hi_lo_lo_lo_lo_lo_8};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo_2 = {regroupV0_hi_6[269:268], regroupV0_hi_6[261:260]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi_2 = {regroupV0_hi_6[285:284], regroupV0_hi_6[277:276]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_6 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo_2 = {regroupV0_hi_6[301:300], regroupV0_hi_6[293:292]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi_2 = {regroupV0_hi_6[317:316], regroupV0_hi_6[309:308]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_6 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi_2, regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_lo_lo_8 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_6, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo_2 = {regroupV0_hi_6[333:332], regroupV0_hi_6[325:324]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi_2 = {regroupV0_hi_6[349:348], regroupV0_hi_6[341:340]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_6 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi_2, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo_2 = {regroupV0_hi_6[365:364], regroupV0_hi_6[357:356]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi_2 = {regroupV0_hi_6[381:380], regroupV0_hi_6[373:372]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_6 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi_2, regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_lo_hi_8 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_6, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_6};
  wire [31:0]        regroupV0_hi_lo_lo_lo_hi_lo_8 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_8, regroupV0_hi_lo_lo_lo_hi_lo_lo_8};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo_2 = {regroupV0_hi_6[397:396], regroupV0_hi_6[389:388]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi_2 = {regroupV0_hi_6[413:412], regroupV0_hi_6[405:404]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_6 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo_2 = {regroupV0_hi_6[429:428], regroupV0_hi_6[421:420]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi_2 = {regroupV0_hi_6[445:444], regroupV0_hi_6[437:436]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_6 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi_2, regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_hi_lo_8 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_6, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo_2 = {regroupV0_hi_6[461:460], regroupV0_hi_6[453:452]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi_2 = {regroupV0_hi_6[477:476], regroupV0_hi_6[469:468]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_6 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi_2, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo_2 = {regroupV0_hi_6[493:492], regroupV0_hi_6[485:484]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi_2 = {regroupV0_hi_6[509:508], regroupV0_hi_6[501:500]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_6 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi_2, regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_hi_hi_8 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_6, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_6};
  wire [31:0]        regroupV0_hi_lo_lo_lo_hi_hi_8 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_8, regroupV0_hi_lo_lo_lo_hi_hi_lo_8};
  wire [63:0]        regroupV0_hi_lo_lo_lo_hi_8 = {regroupV0_hi_lo_lo_lo_hi_hi_8, regroupV0_hi_lo_lo_lo_hi_lo_8};
  wire [127:0]       regroupV0_hi_lo_lo_lo_8 = {regroupV0_hi_lo_lo_lo_hi_8, regroupV0_hi_lo_lo_lo_lo_8};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo_2 = {regroupV0_hi_6[525:524], regroupV0_hi_6[517:516]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi_2 = {regroupV0_hi_6[541:540], regroupV0_hi_6[533:532]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_6 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi_2, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo_2 = {regroupV0_hi_6[557:556], regroupV0_hi_6[549:548]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi_2 = {regroupV0_hi_6[573:572], regroupV0_hi_6[565:564]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_6 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi_2, regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_lo_lo_8 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_6, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo_2 = {regroupV0_hi_6[589:588], regroupV0_hi_6[581:580]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi_2 = {regroupV0_hi_6[605:604], regroupV0_hi_6[597:596]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_6 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi_2, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo_2 = {regroupV0_hi_6[621:620], regroupV0_hi_6[613:612]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi_2 = {regroupV0_hi_6[637:636], regroupV0_hi_6[629:628]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_6 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi_2, regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_lo_hi_8 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_6, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_6};
  wire [31:0]        regroupV0_hi_lo_lo_hi_lo_lo_8 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_8, regroupV0_hi_lo_lo_hi_lo_lo_lo_8};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo_2 = {regroupV0_hi_6[653:652], regroupV0_hi_6[645:644]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi_2 = {regroupV0_hi_6[669:668], regroupV0_hi_6[661:660]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_6 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi_2, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo_2 = {regroupV0_hi_6[685:684], regroupV0_hi_6[677:676]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi_2 = {regroupV0_hi_6[701:700], regroupV0_hi_6[693:692]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_6 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi_2, regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_hi_lo_8 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_6, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo_2 = {regroupV0_hi_6[717:716], regroupV0_hi_6[709:708]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi_2 = {regroupV0_hi_6[733:732], regroupV0_hi_6[725:724]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_6 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi_2, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo_2 = {regroupV0_hi_6[749:748], regroupV0_hi_6[741:740]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi_2 = {regroupV0_hi_6[765:764], regroupV0_hi_6[757:756]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_6 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi_2, regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_hi_hi_8 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_6, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_6};
  wire [31:0]        regroupV0_hi_lo_lo_hi_lo_hi_8 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_8, regroupV0_hi_lo_lo_hi_lo_hi_lo_8};
  wire [63:0]        regroupV0_hi_lo_lo_hi_lo_8 = {regroupV0_hi_lo_lo_hi_lo_hi_8, regroupV0_hi_lo_lo_hi_lo_lo_8};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo_2 = {regroupV0_hi_6[781:780], regroupV0_hi_6[773:772]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi_2 = {regroupV0_hi_6[797:796], regroupV0_hi_6[789:788]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_6 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi_2, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo_2 = {regroupV0_hi_6[813:812], regroupV0_hi_6[805:804]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi_2 = {regroupV0_hi_6[829:828], regroupV0_hi_6[821:820]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_6 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi_2, regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_lo_lo_8 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_6, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo_2 = {regroupV0_hi_6[845:844], regroupV0_hi_6[837:836]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi_2 = {regroupV0_hi_6[861:860], regroupV0_hi_6[853:852]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_6 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi_2, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo_2 = {regroupV0_hi_6[877:876], regroupV0_hi_6[869:868]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi_2 = {regroupV0_hi_6[893:892], regroupV0_hi_6[885:884]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_6 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi_2, regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_lo_hi_8 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_6, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_6};
  wire [31:0]        regroupV0_hi_lo_lo_hi_hi_lo_8 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_8, regroupV0_hi_lo_lo_hi_hi_lo_lo_8};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo_2 = {regroupV0_hi_6[909:908], regroupV0_hi_6[901:900]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi_2 = {regroupV0_hi_6[925:924], regroupV0_hi_6[917:916]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_6 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi_2, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo_2 = {regroupV0_hi_6[941:940], regroupV0_hi_6[933:932]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi_2 = {regroupV0_hi_6[957:956], regroupV0_hi_6[949:948]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_6 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi_2, regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_hi_lo_8 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_6, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo_2 = {regroupV0_hi_6[973:972], regroupV0_hi_6[965:964]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi_2 = {regroupV0_hi_6[989:988], regroupV0_hi_6[981:980]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_6 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi_2, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo_2 = {regroupV0_hi_6[1005:1004], regroupV0_hi_6[997:996]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi_2 = {regroupV0_hi_6[1021:1020], regroupV0_hi_6[1013:1012]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_6 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi_2, regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_hi_hi_8 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_6, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_6};
  wire [31:0]        regroupV0_hi_lo_lo_hi_hi_hi_8 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_8, regroupV0_hi_lo_lo_hi_hi_hi_lo_8};
  wire [63:0]        regroupV0_hi_lo_lo_hi_hi_8 = {regroupV0_hi_lo_lo_hi_hi_hi_8, regroupV0_hi_lo_lo_hi_hi_lo_8};
  wire [127:0]       regroupV0_hi_lo_lo_hi_8 = {regroupV0_hi_lo_lo_hi_hi_8, regroupV0_hi_lo_lo_hi_lo_8};
  wire [255:0]       regroupV0_hi_lo_lo_8 = {regroupV0_hi_lo_lo_hi_8, regroupV0_hi_lo_lo_lo_8};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo_2 = {regroupV0_hi_6[1037:1036], regroupV0_hi_6[1029:1028]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi_2 = {regroupV0_hi_6[1053:1052], regroupV0_hi_6[1045:1044]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_6 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi_2, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo_2 = {regroupV0_hi_6[1069:1068], regroupV0_hi_6[1061:1060]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi_2 = {regroupV0_hi_6[1085:1084], regroupV0_hi_6[1077:1076]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_6 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi_2, regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_lo_lo_8 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_6, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo_2 = {regroupV0_hi_6[1101:1100], regroupV0_hi_6[1093:1092]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi_2 = {regroupV0_hi_6[1117:1116], regroupV0_hi_6[1109:1108]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_6 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi_2, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo_2 = {regroupV0_hi_6[1133:1132], regroupV0_hi_6[1125:1124]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi_2 = {regroupV0_hi_6[1149:1148], regroupV0_hi_6[1141:1140]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_6 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi_2, regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_lo_hi_8 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_6, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_6};
  wire [31:0]        regroupV0_hi_lo_hi_lo_lo_lo_8 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_8, regroupV0_hi_lo_hi_lo_lo_lo_lo_8};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo_2 = {regroupV0_hi_6[1165:1164], regroupV0_hi_6[1157:1156]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi_2 = {regroupV0_hi_6[1181:1180], regroupV0_hi_6[1173:1172]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_6 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi_2, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo_2 = {regroupV0_hi_6[1197:1196], regroupV0_hi_6[1189:1188]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi_2 = {regroupV0_hi_6[1213:1212], regroupV0_hi_6[1205:1204]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_6 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi_2, regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_hi_lo_8 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_6, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo_2 = {regroupV0_hi_6[1229:1228], regroupV0_hi_6[1221:1220]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi_2 = {regroupV0_hi_6[1245:1244], regroupV0_hi_6[1237:1236]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_6 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi_2, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo_2 = {regroupV0_hi_6[1261:1260], regroupV0_hi_6[1253:1252]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi_2 = {regroupV0_hi_6[1277:1276], regroupV0_hi_6[1269:1268]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_6 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi_2, regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_hi_hi_8 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_6, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_6};
  wire [31:0]        regroupV0_hi_lo_hi_lo_lo_hi_8 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_8, regroupV0_hi_lo_hi_lo_lo_hi_lo_8};
  wire [63:0]        regroupV0_hi_lo_hi_lo_lo_8 = {regroupV0_hi_lo_hi_lo_lo_hi_8, regroupV0_hi_lo_hi_lo_lo_lo_8};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo_2 = {regroupV0_hi_6[1293:1292], regroupV0_hi_6[1285:1284]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi_2 = {regroupV0_hi_6[1309:1308], regroupV0_hi_6[1301:1300]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_6 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi_2, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo_2 = {regroupV0_hi_6[1325:1324], regroupV0_hi_6[1317:1316]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi_2 = {regroupV0_hi_6[1341:1340], regroupV0_hi_6[1333:1332]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_6 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi_2, regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_lo_lo_8 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_6, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo_2 = {regroupV0_hi_6[1357:1356], regroupV0_hi_6[1349:1348]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi_2 = {regroupV0_hi_6[1373:1372], regroupV0_hi_6[1365:1364]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_6 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi_2, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo_2 = {regroupV0_hi_6[1389:1388], regroupV0_hi_6[1381:1380]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi_2 = {regroupV0_hi_6[1405:1404], regroupV0_hi_6[1397:1396]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_6 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi_2, regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_lo_hi_8 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_6, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_6};
  wire [31:0]        regroupV0_hi_lo_hi_lo_hi_lo_8 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_8, regroupV0_hi_lo_hi_lo_hi_lo_lo_8};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo_2 = {regroupV0_hi_6[1421:1420], regroupV0_hi_6[1413:1412]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi_2 = {regroupV0_hi_6[1437:1436], regroupV0_hi_6[1429:1428]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_6 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi_2, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo_2 = {regroupV0_hi_6[1453:1452], regroupV0_hi_6[1445:1444]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi_2 = {regroupV0_hi_6[1469:1468], regroupV0_hi_6[1461:1460]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_6 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi_2, regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_hi_lo_8 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_6, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo_2 = {regroupV0_hi_6[1485:1484], regroupV0_hi_6[1477:1476]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi_2 = {regroupV0_hi_6[1501:1500], regroupV0_hi_6[1493:1492]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_6 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi_2, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo_2 = {regroupV0_hi_6[1517:1516], regroupV0_hi_6[1509:1508]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi_2 = {regroupV0_hi_6[1533:1532], regroupV0_hi_6[1525:1524]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_6 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi_2, regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_hi_hi_8 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_6, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_6};
  wire [31:0]        regroupV0_hi_lo_hi_lo_hi_hi_8 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_8, regroupV0_hi_lo_hi_lo_hi_hi_lo_8};
  wire [63:0]        regroupV0_hi_lo_hi_lo_hi_8 = {regroupV0_hi_lo_hi_lo_hi_hi_8, regroupV0_hi_lo_hi_lo_hi_lo_8};
  wire [127:0]       regroupV0_hi_lo_hi_lo_8 = {regroupV0_hi_lo_hi_lo_hi_8, regroupV0_hi_lo_hi_lo_lo_8};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo_2 = {regroupV0_hi_6[1549:1548], regroupV0_hi_6[1541:1540]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi_2 = {regroupV0_hi_6[1565:1564], regroupV0_hi_6[1557:1556]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_6 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi_2, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo_2 = {regroupV0_hi_6[1581:1580], regroupV0_hi_6[1573:1572]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi_2 = {regroupV0_hi_6[1597:1596], regroupV0_hi_6[1589:1588]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_6 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi_2, regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_lo_lo_8 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_6, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo_2 = {regroupV0_hi_6[1613:1612], regroupV0_hi_6[1605:1604]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi_2 = {regroupV0_hi_6[1629:1628], regroupV0_hi_6[1621:1620]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_6 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi_2, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo_2 = {regroupV0_hi_6[1645:1644], regroupV0_hi_6[1637:1636]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi_2 = {regroupV0_hi_6[1661:1660], regroupV0_hi_6[1653:1652]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_6 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi_2, regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_lo_hi_8 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_6, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_6};
  wire [31:0]        regroupV0_hi_lo_hi_hi_lo_lo_8 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_8, regroupV0_hi_lo_hi_hi_lo_lo_lo_8};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo_2 = {regroupV0_hi_6[1677:1676], regroupV0_hi_6[1669:1668]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi_2 = {regroupV0_hi_6[1693:1692], regroupV0_hi_6[1685:1684]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_6 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi_2, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo_2 = {regroupV0_hi_6[1709:1708], regroupV0_hi_6[1701:1700]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi_2 = {regroupV0_hi_6[1725:1724], regroupV0_hi_6[1717:1716]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_6 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi_2, regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_hi_lo_8 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_6, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo_2 = {regroupV0_hi_6[1741:1740], regroupV0_hi_6[1733:1732]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi_2 = {regroupV0_hi_6[1757:1756], regroupV0_hi_6[1749:1748]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_6 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi_2, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo_2 = {regroupV0_hi_6[1773:1772], regroupV0_hi_6[1765:1764]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi_2 = {regroupV0_hi_6[1789:1788], regroupV0_hi_6[1781:1780]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_6 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi_2, regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_hi_hi_8 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_6, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_6};
  wire [31:0]        regroupV0_hi_lo_hi_hi_lo_hi_8 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_8, regroupV0_hi_lo_hi_hi_lo_hi_lo_8};
  wire [63:0]        regroupV0_hi_lo_hi_hi_lo_8 = {regroupV0_hi_lo_hi_hi_lo_hi_8, regroupV0_hi_lo_hi_hi_lo_lo_8};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo_2 = {regroupV0_hi_6[1805:1804], regroupV0_hi_6[1797:1796]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi_2 = {regroupV0_hi_6[1821:1820], regroupV0_hi_6[1813:1812]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_6 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi_2, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo_2 = {regroupV0_hi_6[1837:1836], regroupV0_hi_6[1829:1828]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi_2 = {regroupV0_hi_6[1853:1852], regroupV0_hi_6[1845:1844]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_6 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi_2, regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_lo_lo_8 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_6, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo_2 = {regroupV0_hi_6[1869:1868], regroupV0_hi_6[1861:1860]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi_2 = {regroupV0_hi_6[1885:1884], regroupV0_hi_6[1877:1876]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_6 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi_2, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo_2 = {regroupV0_hi_6[1901:1900], regroupV0_hi_6[1893:1892]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi_2 = {regroupV0_hi_6[1917:1916], regroupV0_hi_6[1909:1908]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_6 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi_2, regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_lo_hi_8 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_6, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_6};
  wire [31:0]        regroupV0_hi_lo_hi_hi_hi_lo_8 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_8, regroupV0_hi_lo_hi_hi_hi_lo_lo_8};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo_2 = {regroupV0_hi_6[1933:1932], regroupV0_hi_6[1925:1924]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi_2 = {regroupV0_hi_6[1949:1948], regroupV0_hi_6[1941:1940]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_6 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi_2, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo_2 = {regroupV0_hi_6[1965:1964], regroupV0_hi_6[1957:1956]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi_2 = {regroupV0_hi_6[1981:1980], regroupV0_hi_6[1973:1972]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_6 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi_2, regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_hi_lo_8 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_6, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo_2 = {regroupV0_hi_6[1997:1996], regroupV0_hi_6[1989:1988]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi_2 = {regroupV0_hi_6[2013:2012], regroupV0_hi_6[2005:2004]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_6 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi_2, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo_2 = {regroupV0_hi_6[2029:2028], regroupV0_hi_6[2021:2020]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi_2 = {regroupV0_hi_6[2045:2044], regroupV0_hi_6[2037:2036]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_6 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi_2, regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_hi_hi_8 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_6, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_6};
  wire [31:0]        regroupV0_hi_lo_hi_hi_hi_hi_8 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_8, regroupV0_hi_lo_hi_hi_hi_hi_lo_8};
  wire [63:0]        regroupV0_hi_lo_hi_hi_hi_8 = {regroupV0_hi_lo_hi_hi_hi_hi_8, regroupV0_hi_lo_hi_hi_hi_lo_8};
  wire [127:0]       regroupV0_hi_lo_hi_hi_8 = {regroupV0_hi_lo_hi_hi_hi_8, regroupV0_hi_lo_hi_hi_lo_8};
  wire [255:0]       regroupV0_hi_lo_hi_8 = {regroupV0_hi_lo_hi_hi_8, regroupV0_hi_lo_hi_lo_8};
  wire [511:0]       regroupV0_hi_lo_8 = {regroupV0_hi_lo_hi_8, regroupV0_hi_lo_lo_8};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo_2 = {regroupV0_hi_6[2061:2060], regroupV0_hi_6[2053:2052]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi_2 = {regroupV0_hi_6[2077:2076], regroupV0_hi_6[2069:2068]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_6 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi_2, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo_2 = {regroupV0_hi_6[2093:2092], regroupV0_hi_6[2085:2084]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi_2 = {regroupV0_hi_6[2109:2108], regroupV0_hi_6[2101:2100]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_6 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi_2, regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_lo_lo_8 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_6, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo_2 = {regroupV0_hi_6[2125:2124], regroupV0_hi_6[2117:2116]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi_2 = {regroupV0_hi_6[2141:2140], regroupV0_hi_6[2133:2132]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_6 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi_2, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo_2 = {regroupV0_hi_6[2157:2156], regroupV0_hi_6[2149:2148]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi_2 = {regroupV0_hi_6[2173:2172], regroupV0_hi_6[2165:2164]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_6 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi_2, regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_lo_hi_8 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_6, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_6};
  wire [31:0]        regroupV0_hi_hi_lo_lo_lo_lo_8 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_8, regroupV0_hi_hi_lo_lo_lo_lo_lo_8};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo_2 = {regroupV0_hi_6[2189:2188], regroupV0_hi_6[2181:2180]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi_2 = {regroupV0_hi_6[2205:2204], regroupV0_hi_6[2197:2196]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_6 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi_2, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo_2 = {regroupV0_hi_6[2221:2220], regroupV0_hi_6[2213:2212]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi_2 = {regroupV0_hi_6[2237:2236], regroupV0_hi_6[2229:2228]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_6 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi_2, regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_hi_lo_8 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_6, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo_2 = {regroupV0_hi_6[2253:2252], regroupV0_hi_6[2245:2244]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi_2 = {regroupV0_hi_6[2269:2268], regroupV0_hi_6[2261:2260]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_6 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi_2, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo_2 = {regroupV0_hi_6[2285:2284], regroupV0_hi_6[2277:2276]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi_2 = {regroupV0_hi_6[2301:2300], regroupV0_hi_6[2293:2292]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_6 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi_2, regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_hi_hi_8 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_6, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_6};
  wire [31:0]        regroupV0_hi_hi_lo_lo_lo_hi_8 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_8, regroupV0_hi_hi_lo_lo_lo_hi_lo_8};
  wire [63:0]        regroupV0_hi_hi_lo_lo_lo_8 = {regroupV0_hi_hi_lo_lo_lo_hi_8, regroupV0_hi_hi_lo_lo_lo_lo_8};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo_2 = {regroupV0_hi_6[2317:2316], regroupV0_hi_6[2309:2308]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi_2 = {regroupV0_hi_6[2333:2332], regroupV0_hi_6[2325:2324]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_6 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi_2, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo_2 = {regroupV0_hi_6[2349:2348], regroupV0_hi_6[2341:2340]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi_2 = {regroupV0_hi_6[2365:2364], regroupV0_hi_6[2357:2356]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_6 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi_2, regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_lo_lo_8 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_6, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo_2 = {regroupV0_hi_6[2381:2380], regroupV0_hi_6[2373:2372]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi_2 = {regroupV0_hi_6[2397:2396], regroupV0_hi_6[2389:2388]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_6 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi_2, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo_2 = {regroupV0_hi_6[2413:2412], regroupV0_hi_6[2405:2404]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi_2 = {regroupV0_hi_6[2429:2428], regroupV0_hi_6[2421:2420]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_6 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi_2, regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_lo_hi_8 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_6, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_6};
  wire [31:0]        regroupV0_hi_hi_lo_lo_hi_lo_8 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_8, regroupV0_hi_hi_lo_lo_hi_lo_lo_8};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo_2 = {regroupV0_hi_6[2445:2444], regroupV0_hi_6[2437:2436]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi_2 = {regroupV0_hi_6[2461:2460], regroupV0_hi_6[2453:2452]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_6 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi_2, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo_2 = {regroupV0_hi_6[2477:2476], regroupV0_hi_6[2469:2468]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi_2 = {regroupV0_hi_6[2493:2492], regroupV0_hi_6[2485:2484]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_6 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi_2, regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_hi_lo_8 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_6, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo_2 = {regroupV0_hi_6[2509:2508], regroupV0_hi_6[2501:2500]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi_2 = {regroupV0_hi_6[2525:2524], regroupV0_hi_6[2517:2516]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_6 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi_2, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo_2 = {regroupV0_hi_6[2541:2540], regroupV0_hi_6[2533:2532]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi_2 = {regroupV0_hi_6[2557:2556], regroupV0_hi_6[2549:2548]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_6 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi_2, regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_hi_hi_8 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_6, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_6};
  wire [31:0]        regroupV0_hi_hi_lo_lo_hi_hi_8 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_8, regroupV0_hi_hi_lo_lo_hi_hi_lo_8};
  wire [63:0]        regroupV0_hi_hi_lo_lo_hi_8 = {regroupV0_hi_hi_lo_lo_hi_hi_8, regroupV0_hi_hi_lo_lo_hi_lo_8};
  wire [127:0]       regroupV0_hi_hi_lo_lo_8 = {regroupV0_hi_hi_lo_lo_hi_8, regroupV0_hi_hi_lo_lo_lo_8};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo_2 = {regroupV0_hi_6[2573:2572], regroupV0_hi_6[2565:2564]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi_2 = {regroupV0_hi_6[2589:2588], regroupV0_hi_6[2581:2580]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_6 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi_2, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo_2 = {regroupV0_hi_6[2605:2604], regroupV0_hi_6[2597:2596]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi_2 = {regroupV0_hi_6[2621:2620], regroupV0_hi_6[2613:2612]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_6 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi_2, regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_lo_lo_8 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_6, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo_2 = {regroupV0_hi_6[2637:2636], regroupV0_hi_6[2629:2628]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi_2 = {regroupV0_hi_6[2653:2652], regroupV0_hi_6[2645:2644]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_6 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi_2, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo_2 = {regroupV0_hi_6[2669:2668], regroupV0_hi_6[2661:2660]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi_2 = {regroupV0_hi_6[2685:2684], regroupV0_hi_6[2677:2676]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_6 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi_2, regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_lo_hi_8 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_6, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_6};
  wire [31:0]        regroupV0_hi_hi_lo_hi_lo_lo_8 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_8, regroupV0_hi_hi_lo_hi_lo_lo_lo_8};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo_2 = {regroupV0_hi_6[2701:2700], regroupV0_hi_6[2693:2692]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi_2 = {regroupV0_hi_6[2717:2716], regroupV0_hi_6[2709:2708]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_6 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi_2, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo_2 = {regroupV0_hi_6[2733:2732], regroupV0_hi_6[2725:2724]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi_2 = {regroupV0_hi_6[2749:2748], regroupV0_hi_6[2741:2740]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_6 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi_2, regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_hi_lo_8 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_6, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo_2 = {regroupV0_hi_6[2765:2764], regroupV0_hi_6[2757:2756]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi_2 = {regroupV0_hi_6[2781:2780], regroupV0_hi_6[2773:2772]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_6 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi_2, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo_2 = {regroupV0_hi_6[2797:2796], regroupV0_hi_6[2789:2788]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi_2 = {regroupV0_hi_6[2813:2812], regroupV0_hi_6[2805:2804]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_6 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi_2, regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_hi_hi_8 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_6, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_6};
  wire [31:0]        regroupV0_hi_hi_lo_hi_lo_hi_8 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_8, regroupV0_hi_hi_lo_hi_lo_hi_lo_8};
  wire [63:0]        regroupV0_hi_hi_lo_hi_lo_8 = {regroupV0_hi_hi_lo_hi_lo_hi_8, regroupV0_hi_hi_lo_hi_lo_lo_8};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo_2 = {regroupV0_hi_6[2829:2828], regroupV0_hi_6[2821:2820]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi_2 = {regroupV0_hi_6[2845:2844], regroupV0_hi_6[2837:2836]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_6 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi_2, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo_2 = {regroupV0_hi_6[2861:2860], regroupV0_hi_6[2853:2852]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi_2 = {regroupV0_hi_6[2877:2876], regroupV0_hi_6[2869:2868]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_6 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi_2, regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_lo_lo_8 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_6, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo_2 = {regroupV0_hi_6[2893:2892], regroupV0_hi_6[2885:2884]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi_2 = {regroupV0_hi_6[2909:2908], regroupV0_hi_6[2901:2900]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_6 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi_2, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo_2 = {regroupV0_hi_6[2925:2924], regroupV0_hi_6[2917:2916]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi_2 = {regroupV0_hi_6[2941:2940], regroupV0_hi_6[2933:2932]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_6 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi_2, regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_lo_hi_8 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_6, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_6};
  wire [31:0]        regroupV0_hi_hi_lo_hi_hi_lo_8 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_8, regroupV0_hi_hi_lo_hi_hi_lo_lo_8};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo_2 = {regroupV0_hi_6[2957:2956], regroupV0_hi_6[2949:2948]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi_2 = {regroupV0_hi_6[2973:2972], regroupV0_hi_6[2965:2964]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_6 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi_2, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo_2 = {regroupV0_hi_6[2989:2988], regroupV0_hi_6[2981:2980]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi_2 = {regroupV0_hi_6[3005:3004], regroupV0_hi_6[2997:2996]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_6 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi_2, regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_hi_lo_8 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_6, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo_2 = {regroupV0_hi_6[3021:3020], regroupV0_hi_6[3013:3012]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi_2 = {regroupV0_hi_6[3037:3036], regroupV0_hi_6[3029:3028]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_6 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi_2, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo_2 = {regroupV0_hi_6[3053:3052], regroupV0_hi_6[3045:3044]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi_2 = {regroupV0_hi_6[3069:3068], regroupV0_hi_6[3061:3060]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_6 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi_2, regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_hi_hi_8 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_6, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_6};
  wire [31:0]        regroupV0_hi_hi_lo_hi_hi_hi_8 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_8, regroupV0_hi_hi_lo_hi_hi_hi_lo_8};
  wire [63:0]        regroupV0_hi_hi_lo_hi_hi_8 = {regroupV0_hi_hi_lo_hi_hi_hi_8, regroupV0_hi_hi_lo_hi_hi_lo_8};
  wire [127:0]       regroupV0_hi_hi_lo_hi_8 = {regroupV0_hi_hi_lo_hi_hi_8, regroupV0_hi_hi_lo_hi_lo_8};
  wire [255:0]       regroupV0_hi_hi_lo_8 = {regroupV0_hi_hi_lo_hi_8, regroupV0_hi_hi_lo_lo_8};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo_2 = {regroupV0_hi_6[3085:3084], regroupV0_hi_6[3077:3076]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi_2 = {regroupV0_hi_6[3101:3100], regroupV0_hi_6[3093:3092]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_6 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi_2, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo_2 = {regroupV0_hi_6[3117:3116], regroupV0_hi_6[3109:3108]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi_2 = {regroupV0_hi_6[3133:3132], regroupV0_hi_6[3125:3124]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_6 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi_2, regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_lo_lo_8 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_6, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo_2 = {regroupV0_hi_6[3149:3148], regroupV0_hi_6[3141:3140]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi_2 = {regroupV0_hi_6[3165:3164], regroupV0_hi_6[3157:3156]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_6 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi_2, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo_2 = {regroupV0_hi_6[3181:3180], regroupV0_hi_6[3173:3172]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi_2 = {regroupV0_hi_6[3197:3196], regroupV0_hi_6[3189:3188]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_6 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi_2, regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_lo_hi_8 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_6, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_6};
  wire [31:0]        regroupV0_hi_hi_hi_lo_lo_lo_8 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_8, regroupV0_hi_hi_hi_lo_lo_lo_lo_8};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo_2 = {regroupV0_hi_6[3213:3212], regroupV0_hi_6[3205:3204]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi_2 = {regroupV0_hi_6[3229:3228], regroupV0_hi_6[3221:3220]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_6 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi_2, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo_2 = {regroupV0_hi_6[3245:3244], regroupV0_hi_6[3237:3236]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi_2 = {regroupV0_hi_6[3261:3260], regroupV0_hi_6[3253:3252]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_6 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi_2, regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_hi_lo_8 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_6, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo_2 = {regroupV0_hi_6[3277:3276], regroupV0_hi_6[3269:3268]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi_2 = {regroupV0_hi_6[3293:3292], regroupV0_hi_6[3285:3284]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_6 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi_2, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo_2 = {regroupV0_hi_6[3309:3308], regroupV0_hi_6[3301:3300]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi_2 = {regroupV0_hi_6[3325:3324], regroupV0_hi_6[3317:3316]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_6 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_hi_hi_8 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_6, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_6};
  wire [31:0]        regroupV0_hi_hi_hi_lo_lo_hi_8 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_8, regroupV0_hi_hi_hi_lo_lo_hi_lo_8};
  wire [63:0]        regroupV0_hi_hi_hi_lo_lo_8 = {regroupV0_hi_hi_hi_lo_lo_hi_8, regroupV0_hi_hi_hi_lo_lo_lo_8};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo_2 = {regroupV0_hi_6[3341:3340], regroupV0_hi_6[3333:3332]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi_2 = {regroupV0_hi_6[3357:3356], regroupV0_hi_6[3349:3348]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_6 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi_2, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo_2 = {regroupV0_hi_6[3373:3372], regroupV0_hi_6[3365:3364]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi_2 = {regroupV0_hi_6[3389:3388], regroupV0_hi_6[3381:3380]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_6 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi_2, regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_lo_lo_8 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_6, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo_2 = {regroupV0_hi_6[3405:3404], regroupV0_hi_6[3397:3396]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi_2 = {regroupV0_hi_6[3421:3420], regroupV0_hi_6[3413:3412]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_6 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi_2, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo_2 = {regroupV0_hi_6[3437:3436], regroupV0_hi_6[3429:3428]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi_2 = {regroupV0_hi_6[3453:3452], regroupV0_hi_6[3445:3444]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_6 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi_2, regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_lo_hi_8 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_6, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_6};
  wire [31:0]        regroupV0_hi_hi_hi_lo_hi_lo_8 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_8, regroupV0_hi_hi_hi_lo_hi_lo_lo_8};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo_2 = {regroupV0_hi_6[3469:3468], regroupV0_hi_6[3461:3460]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi_2 = {regroupV0_hi_6[3485:3484], regroupV0_hi_6[3477:3476]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_6 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi_2, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo_2 = {regroupV0_hi_6[3501:3500], regroupV0_hi_6[3493:3492]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi_2 = {regroupV0_hi_6[3517:3516], regroupV0_hi_6[3509:3508]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_6 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi_2, regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_hi_lo_8 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_6, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo_2 = {regroupV0_hi_6[3533:3532], regroupV0_hi_6[3525:3524]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi_2 = {regroupV0_hi_6[3549:3548], regroupV0_hi_6[3541:3540]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_6 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi_2, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo_2 = {regroupV0_hi_6[3565:3564], regroupV0_hi_6[3557:3556]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi_2 = {regroupV0_hi_6[3581:3580], regroupV0_hi_6[3573:3572]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_6 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_hi_hi_8 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_6, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_6};
  wire [31:0]        regroupV0_hi_hi_hi_lo_hi_hi_8 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_8, regroupV0_hi_hi_hi_lo_hi_hi_lo_8};
  wire [63:0]        regroupV0_hi_hi_hi_lo_hi_8 = {regroupV0_hi_hi_hi_lo_hi_hi_8, regroupV0_hi_hi_hi_lo_hi_lo_8};
  wire [127:0]       regroupV0_hi_hi_hi_lo_8 = {regroupV0_hi_hi_hi_lo_hi_8, regroupV0_hi_hi_hi_lo_lo_8};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo_2 = {regroupV0_hi_6[3597:3596], regroupV0_hi_6[3589:3588]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi_2 = {regroupV0_hi_6[3613:3612], regroupV0_hi_6[3605:3604]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_6 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi_2, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo_2 = {regroupV0_hi_6[3629:3628], regroupV0_hi_6[3621:3620]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi_2 = {regroupV0_hi_6[3645:3644], regroupV0_hi_6[3637:3636]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_6 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi_2, regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_lo_lo_8 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_6, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo_2 = {regroupV0_hi_6[3661:3660], regroupV0_hi_6[3653:3652]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi_2 = {regroupV0_hi_6[3677:3676], regroupV0_hi_6[3669:3668]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_6 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi_2, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo_2 = {regroupV0_hi_6[3693:3692], regroupV0_hi_6[3685:3684]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi_2 = {regroupV0_hi_6[3709:3708], regroupV0_hi_6[3701:3700]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_6 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi_2, regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_lo_hi_8 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_6, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_6};
  wire [31:0]        regroupV0_hi_hi_hi_hi_lo_lo_8 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_8, regroupV0_hi_hi_hi_hi_lo_lo_lo_8};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo_2 = {regroupV0_hi_6[3725:3724], regroupV0_hi_6[3717:3716]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi_2 = {regroupV0_hi_6[3741:3740], regroupV0_hi_6[3733:3732]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_6 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi_2, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo_2 = {regroupV0_hi_6[3757:3756], regroupV0_hi_6[3749:3748]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi_2 = {regroupV0_hi_6[3773:3772], regroupV0_hi_6[3765:3764]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_6 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi_2, regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_hi_lo_8 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_6, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo_2 = {regroupV0_hi_6[3789:3788], regroupV0_hi_6[3781:3780]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi_2 = {regroupV0_hi_6[3805:3804], regroupV0_hi_6[3797:3796]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_6 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi_2, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo_2 = {regroupV0_hi_6[3821:3820], regroupV0_hi_6[3813:3812]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi_2 = {regroupV0_hi_6[3837:3836], regroupV0_hi_6[3829:3828]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_6 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_hi_hi_8 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_6, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_6};
  wire [31:0]        regroupV0_hi_hi_hi_hi_lo_hi_8 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_8, regroupV0_hi_hi_hi_hi_lo_hi_lo_8};
  wire [63:0]        regroupV0_hi_hi_hi_hi_lo_8 = {regroupV0_hi_hi_hi_hi_lo_hi_8, regroupV0_hi_hi_hi_hi_lo_lo_8};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo_2 = {regroupV0_hi_6[3853:3852], regroupV0_hi_6[3845:3844]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi_2 = {regroupV0_hi_6[3869:3868], regroupV0_hi_6[3861:3860]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_6 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi_2, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo_2 = {regroupV0_hi_6[3885:3884], regroupV0_hi_6[3877:3876]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi_2 = {regroupV0_hi_6[3901:3900], regroupV0_hi_6[3893:3892]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_6 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi_2, regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_lo_lo_8 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_6, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo_2 = {regroupV0_hi_6[3917:3916], regroupV0_hi_6[3909:3908]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi_2 = {regroupV0_hi_6[3933:3932], regroupV0_hi_6[3925:3924]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_6 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi_2, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo_2 = {regroupV0_hi_6[3949:3948], regroupV0_hi_6[3941:3940]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi_2 = {regroupV0_hi_6[3965:3964], regroupV0_hi_6[3957:3956]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_6 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi_2, regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_lo_hi_8 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_6, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_6};
  wire [31:0]        regroupV0_hi_hi_hi_hi_hi_lo_8 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_8, regroupV0_hi_hi_hi_hi_hi_lo_lo_8};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo_2 = {regroupV0_hi_6[3981:3980], regroupV0_hi_6[3973:3972]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi_2 = {regroupV0_hi_6[3997:3996], regroupV0_hi_6[3989:3988]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_6 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi_2, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo_2 = {regroupV0_hi_6[4013:4012], regroupV0_hi_6[4005:4004]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi_2 = {regroupV0_hi_6[4029:4028], regroupV0_hi_6[4021:4020]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_6 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi_2, regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_hi_lo_8 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_6, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo_2 = {regroupV0_hi_6[4045:4044], regroupV0_hi_6[4037:4036]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi_2 = {regroupV0_hi_6[4061:4060], regroupV0_hi_6[4053:4052]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_6 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi_2, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo_2 = {regroupV0_hi_6[4077:4076], regroupV0_hi_6[4069:4068]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi_2 = {regroupV0_hi_6[4093:4092], regroupV0_hi_6[4085:4084]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_6 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_hi_hi_8 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_6, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_6};
  wire [31:0]        regroupV0_hi_hi_hi_hi_hi_hi_8 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_8, regroupV0_hi_hi_hi_hi_hi_hi_lo_8};
  wire [63:0]        regroupV0_hi_hi_hi_hi_hi_8 = {regroupV0_hi_hi_hi_hi_hi_hi_8, regroupV0_hi_hi_hi_hi_hi_lo_8};
  wire [127:0]       regroupV0_hi_hi_hi_hi_8 = {regroupV0_hi_hi_hi_hi_hi_8, regroupV0_hi_hi_hi_hi_lo_8};
  wire [255:0]       regroupV0_hi_hi_hi_8 = {regroupV0_hi_hi_hi_hi_8, regroupV0_hi_hi_hi_lo_8};
  wire [511:0]       regroupV0_hi_hi_8 = {regroupV0_hi_hi_hi_8, regroupV0_hi_hi_lo_8};
  wire [1023:0]      regroupV0_hi_9 = {regroupV0_hi_hi_8, regroupV0_hi_lo_8};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo_3 = {regroupV0_lo_6[15:14], regroupV0_lo_6[7:6]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi_3 = {regroupV0_lo_6[31:30], regroupV0_lo_6[23:22]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_7 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo_3 = {regroupV0_lo_6[47:46], regroupV0_lo_6[39:38]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi_3 = {regroupV0_lo_6[63:62], regroupV0_lo_6[55:54]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_7 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi_3, regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_lo_lo_9 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_7, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo_3 = {regroupV0_lo_6[79:78], regroupV0_lo_6[71:70]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi_3 = {regroupV0_lo_6[95:94], regroupV0_lo_6[87:86]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_7 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi_3, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo_3 = {regroupV0_lo_6[111:110], regroupV0_lo_6[103:102]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi_3 = {regroupV0_lo_6[127:126], regroupV0_lo_6[119:118]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_7 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi_3, regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_lo_hi_9 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_7, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_7};
  wire [31:0]        regroupV0_lo_lo_lo_lo_lo_lo_9 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_9, regroupV0_lo_lo_lo_lo_lo_lo_lo_9};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo_3 = {regroupV0_lo_6[143:142], regroupV0_lo_6[135:134]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi_3 = {regroupV0_lo_6[159:158], regroupV0_lo_6[151:150]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_7 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo_3 = {regroupV0_lo_6[175:174], regroupV0_lo_6[167:166]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi_3 = {regroupV0_lo_6[191:190], regroupV0_lo_6[183:182]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_7 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi_3, regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_hi_lo_9 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_7, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo_3 = {regroupV0_lo_6[207:206], regroupV0_lo_6[199:198]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi_3 = {regroupV0_lo_6[223:222], regroupV0_lo_6[215:214]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_7 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi_3, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo_3 = {regroupV0_lo_6[239:238], regroupV0_lo_6[231:230]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi_3 = {regroupV0_lo_6[255:254], regroupV0_lo_6[247:246]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_7 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi_3, regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_hi_hi_9 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_7, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_7};
  wire [31:0]        regroupV0_lo_lo_lo_lo_lo_hi_9 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_9, regroupV0_lo_lo_lo_lo_lo_hi_lo_9};
  wire [63:0]        regroupV0_lo_lo_lo_lo_lo_9 = {regroupV0_lo_lo_lo_lo_lo_hi_9, regroupV0_lo_lo_lo_lo_lo_lo_9};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo_3 = {regroupV0_lo_6[271:270], regroupV0_lo_6[263:262]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi_3 = {regroupV0_lo_6[287:286], regroupV0_lo_6[279:278]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_7 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo_3 = {regroupV0_lo_6[303:302], regroupV0_lo_6[295:294]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi_3 = {regroupV0_lo_6[319:318], regroupV0_lo_6[311:310]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_7 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi_3, regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_lo_lo_9 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_7, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo_3 = {regroupV0_lo_6[335:334], regroupV0_lo_6[327:326]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi_3 = {regroupV0_lo_6[351:350], regroupV0_lo_6[343:342]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_7 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi_3, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo_3 = {regroupV0_lo_6[367:366], regroupV0_lo_6[359:358]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi_3 = {regroupV0_lo_6[383:382], regroupV0_lo_6[375:374]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_7 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi_3, regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_lo_hi_9 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_7, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_7};
  wire [31:0]        regroupV0_lo_lo_lo_lo_hi_lo_9 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_9, regroupV0_lo_lo_lo_lo_hi_lo_lo_9};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo_3 = {regroupV0_lo_6[399:398], regroupV0_lo_6[391:390]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi_3 = {regroupV0_lo_6[415:414], regroupV0_lo_6[407:406]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_7 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo_3 = {regroupV0_lo_6[431:430], regroupV0_lo_6[423:422]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi_3 = {regroupV0_lo_6[447:446], regroupV0_lo_6[439:438]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_7 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi_3, regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_hi_lo_9 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_7, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo_3 = {regroupV0_lo_6[463:462], regroupV0_lo_6[455:454]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi_3 = {regroupV0_lo_6[479:478], regroupV0_lo_6[471:470]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_7 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi_3, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo_3 = {regroupV0_lo_6[495:494], regroupV0_lo_6[487:486]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi_3 = {regroupV0_lo_6[511:510], regroupV0_lo_6[503:502]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_7 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi_3, regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_hi_hi_9 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_7, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_7};
  wire [31:0]        regroupV0_lo_lo_lo_lo_hi_hi_9 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_9, regroupV0_lo_lo_lo_lo_hi_hi_lo_9};
  wire [63:0]        regroupV0_lo_lo_lo_lo_hi_9 = {regroupV0_lo_lo_lo_lo_hi_hi_9, regroupV0_lo_lo_lo_lo_hi_lo_9};
  wire [127:0]       regroupV0_lo_lo_lo_lo_9 = {regroupV0_lo_lo_lo_lo_hi_9, regroupV0_lo_lo_lo_lo_lo_9};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo_3 = {regroupV0_lo_6[527:526], regroupV0_lo_6[519:518]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi_3 = {regroupV0_lo_6[543:542], regroupV0_lo_6[535:534]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_7 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo_3 = {regroupV0_lo_6[559:558], regroupV0_lo_6[551:550]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi_3 = {regroupV0_lo_6[575:574], regroupV0_lo_6[567:566]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_7 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi_3, regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_lo_lo_9 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_7, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo_3 = {regroupV0_lo_6[591:590], regroupV0_lo_6[583:582]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi_3 = {regroupV0_lo_6[607:606], regroupV0_lo_6[599:598]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_7 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi_3, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo_3 = {regroupV0_lo_6[623:622], regroupV0_lo_6[615:614]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi_3 = {regroupV0_lo_6[639:638], regroupV0_lo_6[631:630]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_7 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi_3, regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_lo_hi_9 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_7, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_7};
  wire [31:0]        regroupV0_lo_lo_lo_hi_lo_lo_9 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_9, regroupV0_lo_lo_lo_hi_lo_lo_lo_9};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo_3 = {regroupV0_lo_6[655:654], regroupV0_lo_6[647:646]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi_3 = {regroupV0_lo_6[671:670], regroupV0_lo_6[663:662]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_7 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi_3, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo_3 = {regroupV0_lo_6[687:686], regroupV0_lo_6[679:678]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi_3 = {regroupV0_lo_6[703:702], regroupV0_lo_6[695:694]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_7 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi_3, regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_hi_lo_9 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_7, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo_3 = {regroupV0_lo_6[719:718], regroupV0_lo_6[711:710]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi_3 = {regroupV0_lo_6[735:734], regroupV0_lo_6[727:726]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_7 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi_3, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo_3 = {regroupV0_lo_6[751:750], regroupV0_lo_6[743:742]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi_3 = {regroupV0_lo_6[767:766], regroupV0_lo_6[759:758]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_7 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi_3, regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_hi_hi_9 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_7, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_7};
  wire [31:0]        regroupV0_lo_lo_lo_hi_lo_hi_9 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_9, regroupV0_lo_lo_lo_hi_lo_hi_lo_9};
  wire [63:0]        regroupV0_lo_lo_lo_hi_lo_9 = {regroupV0_lo_lo_lo_hi_lo_hi_9, regroupV0_lo_lo_lo_hi_lo_lo_9};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo_3 = {regroupV0_lo_6[783:782], regroupV0_lo_6[775:774]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi_3 = {regroupV0_lo_6[799:798], regroupV0_lo_6[791:790]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_7 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo_3 = {regroupV0_lo_6[815:814], regroupV0_lo_6[807:806]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi_3 = {regroupV0_lo_6[831:830], regroupV0_lo_6[823:822]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_7 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi_3, regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_lo_lo_9 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_7, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo_3 = {regroupV0_lo_6[847:846], regroupV0_lo_6[839:838]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi_3 = {regroupV0_lo_6[863:862], regroupV0_lo_6[855:854]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_7 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi_3, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo_3 = {regroupV0_lo_6[879:878], regroupV0_lo_6[871:870]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi_3 = {regroupV0_lo_6[895:894], regroupV0_lo_6[887:886]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_7 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi_3, regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_lo_hi_9 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_7, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_7};
  wire [31:0]        regroupV0_lo_lo_lo_hi_hi_lo_9 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_9, regroupV0_lo_lo_lo_hi_hi_lo_lo_9};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo_3 = {regroupV0_lo_6[911:910], regroupV0_lo_6[903:902]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi_3 = {regroupV0_lo_6[927:926], regroupV0_lo_6[919:918]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_7 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi_3, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo_3 = {regroupV0_lo_6[943:942], regroupV0_lo_6[935:934]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi_3 = {regroupV0_lo_6[959:958], regroupV0_lo_6[951:950]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_7 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi_3, regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_hi_lo_9 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_7, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo_3 = {regroupV0_lo_6[975:974], regroupV0_lo_6[967:966]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi_3 = {regroupV0_lo_6[991:990], regroupV0_lo_6[983:982]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_7 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi_3, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo_3 = {regroupV0_lo_6[1007:1006], regroupV0_lo_6[999:998]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi_3 = {regroupV0_lo_6[1023:1022], regroupV0_lo_6[1015:1014]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_7 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi_3, regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_hi_hi_9 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_7, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_7};
  wire [31:0]        regroupV0_lo_lo_lo_hi_hi_hi_9 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_9, regroupV0_lo_lo_lo_hi_hi_hi_lo_9};
  wire [63:0]        regroupV0_lo_lo_lo_hi_hi_9 = {regroupV0_lo_lo_lo_hi_hi_hi_9, regroupV0_lo_lo_lo_hi_hi_lo_9};
  wire [127:0]       regroupV0_lo_lo_lo_hi_9 = {regroupV0_lo_lo_lo_hi_hi_9, regroupV0_lo_lo_lo_hi_lo_9};
  wire [255:0]       regroupV0_lo_lo_lo_9 = {regroupV0_lo_lo_lo_hi_9, regroupV0_lo_lo_lo_lo_9};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo_3 = {regroupV0_lo_6[1039:1038], regroupV0_lo_6[1031:1030]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi_3 = {regroupV0_lo_6[1055:1054], regroupV0_lo_6[1047:1046]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_7 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi_3, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo_3 = {regroupV0_lo_6[1071:1070], regroupV0_lo_6[1063:1062]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi_3 = {regroupV0_lo_6[1087:1086], regroupV0_lo_6[1079:1078]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_7 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi_3, regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_lo_lo_9 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_7, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo_3 = {regroupV0_lo_6[1103:1102], regroupV0_lo_6[1095:1094]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi_3 = {regroupV0_lo_6[1119:1118], regroupV0_lo_6[1111:1110]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_7 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi_3, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo_3 = {regroupV0_lo_6[1135:1134], regroupV0_lo_6[1127:1126]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi_3 = {regroupV0_lo_6[1151:1150], regroupV0_lo_6[1143:1142]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_7 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi_3, regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_lo_hi_9 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_7, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_7};
  wire [31:0]        regroupV0_lo_lo_hi_lo_lo_lo_9 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_9, regroupV0_lo_lo_hi_lo_lo_lo_lo_9};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo_3 = {regroupV0_lo_6[1167:1166], regroupV0_lo_6[1159:1158]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi_3 = {regroupV0_lo_6[1183:1182], regroupV0_lo_6[1175:1174]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_7 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi_3, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo_3 = {regroupV0_lo_6[1199:1198], regroupV0_lo_6[1191:1190]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi_3 = {regroupV0_lo_6[1215:1214], regroupV0_lo_6[1207:1206]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_7 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi_3, regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_hi_lo_9 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_7, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo_3 = {regroupV0_lo_6[1231:1230], regroupV0_lo_6[1223:1222]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi_3 = {regroupV0_lo_6[1247:1246], regroupV0_lo_6[1239:1238]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_7 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi_3, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo_3 = {regroupV0_lo_6[1263:1262], regroupV0_lo_6[1255:1254]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi_3 = {regroupV0_lo_6[1279:1278], regroupV0_lo_6[1271:1270]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_7 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi_3, regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_hi_hi_9 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_7, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_7};
  wire [31:0]        regroupV0_lo_lo_hi_lo_lo_hi_9 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_9, regroupV0_lo_lo_hi_lo_lo_hi_lo_9};
  wire [63:0]        regroupV0_lo_lo_hi_lo_lo_9 = {regroupV0_lo_lo_hi_lo_lo_hi_9, regroupV0_lo_lo_hi_lo_lo_lo_9};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo_3 = {regroupV0_lo_6[1295:1294], regroupV0_lo_6[1287:1286]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi_3 = {regroupV0_lo_6[1311:1310], regroupV0_lo_6[1303:1302]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_7 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi_3, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo_3 = {regroupV0_lo_6[1327:1326], regroupV0_lo_6[1319:1318]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi_3 = {regroupV0_lo_6[1343:1342], regroupV0_lo_6[1335:1334]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_7 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi_3, regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_lo_lo_9 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_7, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo_3 = {regroupV0_lo_6[1359:1358], regroupV0_lo_6[1351:1350]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi_3 = {regroupV0_lo_6[1375:1374], regroupV0_lo_6[1367:1366]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_7 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi_3, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo_3 = {regroupV0_lo_6[1391:1390], regroupV0_lo_6[1383:1382]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi_3 = {regroupV0_lo_6[1407:1406], regroupV0_lo_6[1399:1398]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_7 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi_3, regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_lo_hi_9 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_7, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_7};
  wire [31:0]        regroupV0_lo_lo_hi_lo_hi_lo_9 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_9, regroupV0_lo_lo_hi_lo_hi_lo_lo_9};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo_3 = {regroupV0_lo_6[1423:1422], regroupV0_lo_6[1415:1414]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi_3 = {regroupV0_lo_6[1439:1438], regroupV0_lo_6[1431:1430]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_7 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi_3, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo_3 = {regroupV0_lo_6[1455:1454], regroupV0_lo_6[1447:1446]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi_3 = {regroupV0_lo_6[1471:1470], regroupV0_lo_6[1463:1462]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_7 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi_3, regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_hi_lo_9 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_7, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo_3 = {regroupV0_lo_6[1487:1486], regroupV0_lo_6[1479:1478]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi_3 = {regroupV0_lo_6[1503:1502], regroupV0_lo_6[1495:1494]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_7 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi_3, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo_3 = {regroupV0_lo_6[1519:1518], regroupV0_lo_6[1511:1510]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi_3 = {regroupV0_lo_6[1535:1534], regroupV0_lo_6[1527:1526]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_7 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi_3, regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_hi_hi_9 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_7, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_7};
  wire [31:0]        regroupV0_lo_lo_hi_lo_hi_hi_9 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_9, regroupV0_lo_lo_hi_lo_hi_hi_lo_9};
  wire [63:0]        regroupV0_lo_lo_hi_lo_hi_9 = {regroupV0_lo_lo_hi_lo_hi_hi_9, regroupV0_lo_lo_hi_lo_hi_lo_9};
  wire [127:0]       regroupV0_lo_lo_hi_lo_9 = {regroupV0_lo_lo_hi_lo_hi_9, regroupV0_lo_lo_hi_lo_lo_9};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo_3 = {regroupV0_lo_6[1551:1550], regroupV0_lo_6[1543:1542]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi_3 = {regroupV0_lo_6[1567:1566], regroupV0_lo_6[1559:1558]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_7 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi_3, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo_3 = {regroupV0_lo_6[1583:1582], regroupV0_lo_6[1575:1574]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi_3 = {regroupV0_lo_6[1599:1598], regroupV0_lo_6[1591:1590]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_7 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi_3, regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_lo_lo_9 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_7, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo_3 = {regroupV0_lo_6[1615:1614], regroupV0_lo_6[1607:1606]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi_3 = {regroupV0_lo_6[1631:1630], regroupV0_lo_6[1623:1622]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_7 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi_3, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo_3 = {regroupV0_lo_6[1647:1646], regroupV0_lo_6[1639:1638]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi_3 = {regroupV0_lo_6[1663:1662], regroupV0_lo_6[1655:1654]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_7 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi_3, regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_lo_hi_9 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_7, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_7};
  wire [31:0]        regroupV0_lo_lo_hi_hi_lo_lo_9 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_9, regroupV0_lo_lo_hi_hi_lo_lo_lo_9};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo_3 = {regroupV0_lo_6[1679:1678], regroupV0_lo_6[1671:1670]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi_3 = {regroupV0_lo_6[1695:1694], regroupV0_lo_6[1687:1686]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_7 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi_3, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo_3 = {regroupV0_lo_6[1711:1710], regroupV0_lo_6[1703:1702]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi_3 = {regroupV0_lo_6[1727:1726], regroupV0_lo_6[1719:1718]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_7 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi_3, regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_hi_lo_9 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_7, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo_3 = {regroupV0_lo_6[1743:1742], regroupV0_lo_6[1735:1734]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi_3 = {regroupV0_lo_6[1759:1758], regroupV0_lo_6[1751:1750]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_7 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi_3, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo_3 = {regroupV0_lo_6[1775:1774], regroupV0_lo_6[1767:1766]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi_3 = {regroupV0_lo_6[1791:1790], regroupV0_lo_6[1783:1782]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_7 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi_3, regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_hi_hi_9 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_7, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_7};
  wire [31:0]        regroupV0_lo_lo_hi_hi_lo_hi_9 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_9, regroupV0_lo_lo_hi_hi_lo_hi_lo_9};
  wire [63:0]        regroupV0_lo_lo_hi_hi_lo_9 = {regroupV0_lo_lo_hi_hi_lo_hi_9, regroupV0_lo_lo_hi_hi_lo_lo_9};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo_3 = {regroupV0_lo_6[1807:1806], regroupV0_lo_6[1799:1798]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi_3 = {regroupV0_lo_6[1823:1822], regroupV0_lo_6[1815:1814]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_7 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi_3, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo_3 = {regroupV0_lo_6[1839:1838], regroupV0_lo_6[1831:1830]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi_3 = {regroupV0_lo_6[1855:1854], regroupV0_lo_6[1847:1846]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_7 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi_3, regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_lo_lo_9 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_7, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo_3 = {regroupV0_lo_6[1871:1870], regroupV0_lo_6[1863:1862]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi_3 = {regroupV0_lo_6[1887:1886], regroupV0_lo_6[1879:1878]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_7 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi_3, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo_3 = {regroupV0_lo_6[1903:1902], regroupV0_lo_6[1895:1894]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi_3 = {regroupV0_lo_6[1919:1918], regroupV0_lo_6[1911:1910]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_7 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi_3, regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_lo_hi_9 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_7, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_7};
  wire [31:0]        regroupV0_lo_lo_hi_hi_hi_lo_9 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_9, regroupV0_lo_lo_hi_hi_hi_lo_lo_9};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo_3 = {regroupV0_lo_6[1935:1934], regroupV0_lo_6[1927:1926]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi_3 = {regroupV0_lo_6[1951:1950], regroupV0_lo_6[1943:1942]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_7 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi_3, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo_3 = {regroupV0_lo_6[1967:1966], regroupV0_lo_6[1959:1958]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi_3 = {regroupV0_lo_6[1983:1982], regroupV0_lo_6[1975:1974]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_7 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi_3, regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_hi_lo_9 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_7, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo_3 = {regroupV0_lo_6[1999:1998], regroupV0_lo_6[1991:1990]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi_3 = {regroupV0_lo_6[2015:2014], regroupV0_lo_6[2007:2006]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_7 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi_3, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo_3 = {regroupV0_lo_6[2031:2030], regroupV0_lo_6[2023:2022]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi_3 = {regroupV0_lo_6[2047:2046], regroupV0_lo_6[2039:2038]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_7 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi_3, regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_hi_hi_9 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_7, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_7};
  wire [31:0]        regroupV0_lo_lo_hi_hi_hi_hi_9 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_9, regroupV0_lo_lo_hi_hi_hi_hi_lo_9};
  wire [63:0]        regroupV0_lo_lo_hi_hi_hi_9 = {regroupV0_lo_lo_hi_hi_hi_hi_9, regroupV0_lo_lo_hi_hi_hi_lo_9};
  wire [127:0]       regroupV0_lo_lo_hi_hi_9 = {regroupV0_lo_lo_hi_hi_hi_9, regroupV0_lo_lo_hi_hi_lo_9};
  wire [255:0]       regroupV0_lo_lo_hi_9 = {regroupV0_lo_lo_hi_hi_9, regroupV0_lo_lo_hi_lo_9};
  wire [511:0]       regroupV0_lo_lo_9 = {regroupV0_lo_lo_hi_9, regroupV0_lo_lo_lo_9};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo_3 = {regroupV0_lo_6[2063:2062], regroupV0_lo_6[2055:2054]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi_3 = {regroupV0_lo_6[2079:2078], regroupV0_lo_6[2071:2070]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_7 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi_3, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo_3 = {regroupV0_lo_6[2095:2094], regroupV0_lo_6[2087:2086]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi_3 = {regroupV0_lo_6[2111:2110], regroupV0_lo_6[2103:2102]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_7 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi_3, regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_lo_lo_9 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_7, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo_3 = {regroupV0_lo_6[2127:2126], regroupV0_lo_6[2119:2118]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi_3 = {regroupV0_lo_6[2143:2142], regroupV0_lo_6[2135:2134]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_7 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi_3, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo_3 = {regroupV0_lo_6[2159:2158], regroupV0_lo_6[2151:2150]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi_3 = {regroupV0_lo_6[2175:2174], regroupV0_lo_6[2167:2166]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_7 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi_3, regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_lo_hi_9 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_7, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_7};
  wire [31:0]        regroupV0_lo_hi_lo_lo_lo_lo_9 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_9, regroupV0_lo_hi_lo_lo_lo_lo_lo_9};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo_3 = {regroupV0_lo_6[2191:2190], regroupV0_lo_6[2183:2182]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi_3 = {regroupV0_lo_6[2207:2206], regroupV0_lo_6[2199:2198]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_7 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi_3, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo_3 = {regroupV0_lo_6[2223:2222], regroupV0_lo_6[2215:2214]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi_3 = {regroupV0_lo_6[2239:2238], regroupV0_lo_6[2231:2230]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_7 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi_3, regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_hi_lo_9 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_7, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo_3 = {regroupV0_lo_6[2255:2254], regroupV0_lo_6[2247:2246]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi_3 = {regroupV0_lo_6[2271:2270], regroupV0_lo_6[2263:2262]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_7 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi_3, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo_3 = {regroupV0_lo_6[2287:2286], regroupV0_lo_6[2279:2278]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi_3 = {regroupV0_lo_6[2303:2302], regroupV0_lo_6[2295:2294]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_7 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi_3, regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_hi_hi_9 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_7, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_7};
  wire [31:0]        regroupV0_lo_hi_lo_lo_lo_hi_9 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_9, regroupV0_lo_hi_lo_lo_lo_hi_lo_9};
  wire [63:0]        regroupV0_lo_hi_lo_lo_lo_9 = {regroupV0_lo_hi_lo_lo_lo_hi_9, regroupV0_lo_hi_lo_lo_lo_lo_9};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo_3 = {regroupV0_lo_6[2319:2318], regroupV0_lo_6[2311:2310]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi_3 = {regroupV0_lo_6[2335:2334], regroupV0_lo_6[2327:2326]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_7 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi_3, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo_3 = {regroupV0_lo_6[2351:2350], regroupV0_lo_6[2343:2342]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi_3 = {regroupV0_lo_6[2367:2366], regroupV0_lo_6[2359:2358]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_7 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi_3, regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_lo_lo_9 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_7, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo_3 = {regroupV0_lo_6[2383:2382], regroupV0_lo_6[2375:2374]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi_3 = {regroupV0_lo_6[2399:2398], regroupV0_lo_6[2391:2390]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_7 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi_3, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo_3 = {regroupV0_lo_6[2415:2414], regroupV0_lo_6[2407:2406]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi_3 = {regroupV0_lo_6[2431:2430], regroupV0_lo_6[2423:2422]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_7 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi_3, regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_lo_hi_9 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_7, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_7};
  wire [31:0]        regroupV0_lo_hi_lo_lo_hi_lo_9 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_9, regroupV0_lo_hi_lo_lo_hi_lo_lo_9};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo_3 = {regroupV0_lo_6[2447:2446], regroupV0_lo_6[2439:2438]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi_3 = {regroupV0_lo_6[2463:2462], regroupV0_lo_6[2455:2454]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_7 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi_3, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo_3 = {regroupV0_lo_6[2479:2478], regroupV0_lo_6[2471:2470]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi_3 = {regroupV0_lo_6[2495:2494], regroupV0_lo_6[2487:2486]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_7 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi_3, regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_hi_lo_9 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_7, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo_3 = {regroupV0_lo_6[2511:2510], regroupV0_lo_6[2503:2502]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi_3 = {regroupV0_lo_6[2527:2526], regroupV0_lo_6[2519:2518]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_7 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi_3, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo_3 = {regroupV0_lo_6[2543:2542], regroupV0_lo_6[2535:2534]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi_3 = {regroupV0_lo_6[2559:2558], regroupV0_lo_6[2551:2550]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_7 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi_3, regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_hi_hi_9 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_7, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_7};
  wire [31:0]        regroupV0_lo_hi_lo_lo_hi_hi_9 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_9, regroupV0_lo_hi_lo_lo_hi_hi_lo_9};
  wire [63:0]        regroupV0_lo_hi_lo_lo_hi_9 = {regroupV0_lo_hi_lo_lo_hi_hi_9, regroupV0_lo_hi_lo_lo_hi_lo_9};
  wire [127:0]       regroupV0_lo_hi_lo_lo_9 = {regroupV0_lo_hi_lo_lo_hi_9, regroupV0_lo_hi_lo_lo_lo_9};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo_3 = {regroupV0_lo_6[2575:2574], regroupV0_lo_6[2567:2566]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi_3 = {regroupV0_lo_6[2591:2590], regroupV0_lo_6[2583:2582]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_7 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi_3, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo_3 = {regroupV0_lo_6[2607:2606], regroupV0_lo_6[2599:2598]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi_3 = {regroupV0_lo_6[2623:2622], regroupV0_lo_6[2615:2614]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_7 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi_3, regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_lo_lo_9 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_7, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo_3 = {regroupV0_lo_6[2639:2638], regroupV0_lo_6[2631:2630]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi_3 = {regroupV0_lo_6[2655:2654], regroupV0_lo_6[2647:2646]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_7 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi_3, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo_3 = {regroupV0_lo_6[2671:2670], regroupV0_lo_6[2663:2662]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi_3 = {regroupV0_lo_6[2687:2686], regroupV0_lo_6[2679:2678]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_7 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi_3, regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_lo_hi_9 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_7, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_7};
  wire [31:0]        regroupV0_lo_hi_lo_hi_lo_lo_9 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_9, regroupV0_lo_hi_lo_hi_lo_lo_lo_9};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo_3 = {regroupV0_lo_6[2703:2702], regroupV0_lo_6[2695:2694]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi_3 = {regroupV0_lo_6[2719:2718], regroupV0_lo_6[2711:2710]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_7 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi_3, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo_3 = {regroupV0_lo_6[2735:2734], regroupV0_lo_6[2727:2726]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi_3 = {regroupV0_lo_6[2751:2750], regroupV0_lo_6[2743:2742]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_7 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi_3, regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_hi_lo_9 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_7, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo_3 = {regroupV0_lo_6[2767:2766], regroupV0_lo_6[2759:2758]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi_3 = {regroupV0_lo_6[2783:2782], regroupV0_lo_6[2775:2774]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_7 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi_3, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo_3 = {regroupV0_lo_6[2799:2798], regroupV0_lo_6[2791:2790]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi_3 = {regroupV0_lo_6[2815:2814], regroupV0_lo_6[2807:2806]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_7 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi_3, regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_hi_hi_9 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_7, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_7};
  wire [31:0]        regroupV0_lo_hi_lo_hi_lo_hi_9 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_9, regroupV0_lo_hi_lo_hi_lo_hi_lo_9};
  wire [63:0]        regroupV0_lo_hi_lo_hi_lo_9 = {regroupV0_lo_hi_lo_hi_lo_hi_9, regroupV0_lo_hi_lo_hi_lo_lo_9};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo_3 = {regroupV0_lo_6[2831:2830], regroupV0_lo_6[2823:2822]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi_3 = {regroupV0_lo_6[2847:2846], regroupV0_lo_6[2839:2838]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_7 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi_3, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo_3 = {regroupV0_lo_6[2863:2862], regroupV0_lo_6[2855:2854]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi_3 = {regroupV0_lo_6[2879:2878], regroupV0_lo_6[2871:2870]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_7 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi_3, regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_lo_lo_9 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_7, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo_3 = {regroupV0_lo_6[2895:2894], regroupV0_lo_6[2887:2886]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi_3 = {regroupV0_lo_6[2911:2910], regroupV0_lo_6[2903:2902]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_7 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi_3, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo_3 = {regroupV0_lo_6[2927:2926], regroupV0_lo_6[2919:2918]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi_3 = {regroupV0_lo_6[2943:2942], regroupV0_lo_6[2935:2934]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_7 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi_3, regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_lo_hi_9 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_7, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_7};
  wire [31:0]        regroupV0_lo_hi_lo_hi_hi_lo_9 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_9, regroupV0_lo_hi_lo_hi_hi_lo_lo_9};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo_3 = {regroupV0_lo_6[2959:2958], regroupV0_lo_6[2951:2950]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi_3 = {regroupV0_lo_6[2975:2974], regroupV0_lo_6[2967:2966]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_7 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi_3, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo_3 = {regroupV0_lo_6[2991:2990], regroupV0_lo_6[2983:2982]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi_3 = {regroupV0_lo_6[3007:3006], regroupV0_lo_6[2999:2998]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_7 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi_3, regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_hi_lo_9 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_7, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo_3 = {regroupV0_lo_6[3023:3022], regroupV0_lo_6[3015:3014]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi_3 = {regroupV0_lo_6[3039:3038], regroupV0_lo_6[3031:3030]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_7 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi_3, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo_3 = {regroupV0_lo_6[3055:3054], regroupV0_lo_6[3047:3046]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi_3 = {regroupV0_lo_6[3071:3070], regroupV0_lo_6[3063:3062]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_7 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi_3, regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_hi_hi_9 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_7, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_7};
  wire [31:0]        regroupV0_lo_hi_lo_hi_hi_hi_9 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_9, regroupV0_lo_hi_lo_hi_hi_hi_lo_9};
  wire [63:0]        regroupV0_lo_hi_lo_hi_hi_9 = {regroupV0_lo_hi_lo_hi_hi_hi_9, regroupV0_lo_hi_lo_hi_hi_lo_9};
  wire [127:0]       regroupV0_lo_hi_lo_hi_9 = {regroupV0_lo_hi_lo_hi_hi_9, regroupV0_lo_hi_lo_hi_lo_9};
  wire [255:0]       regroupV0_lo_hi_lo_9 = {regroupV0_lo_hi_lo_hi_9, regroupV0_lo_hi_lo_lo_9};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo_3 = {regroupV0_lo_6[3087:3086], regroupV0_lo_6[3079:3078]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi_3 = {regroupV0_lo_6[3103:3102], regroupV0_lo_6[3095:3094]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_7 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi_3, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo_3 = {regroupV0_lo_6[3119:3118], regroupV0_lo_6[3111:3110]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi_3 = {regroupV0_lo_6[3135:3134], regroupV0_lo_6[3127:3126]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_7 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi_3, regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_lo_lo_9 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_7, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo_3 = {regroupV0_lo_6[3151:3150], regroupV0_lo_6[3143:3142]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi_3 = {regroupV0_lo_6[3167:3166], regroupV0_lo_6[3159:3158]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_7 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi_3, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo_3 = {regroupV0_lo_6[3183:3182], regroupV0_lo_6[3175:3174]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi_3 = {regroupV0_lo_6[3199:3198], regroupV0_lo_6[3191:3190]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_7 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi_3, regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_lo_hi_9 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_7, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_7};
  wire [31:0]        regroupV0_lo_hi_hi_lo_lo_lo_9 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_9, regroupV0_lo_hi_hi_lo_lo_lo_lo_9};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo_3 = {regroupV0_lo_6[3215:3214], regroupV0_lo_6[3207:3206]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi_3 = {regroupV0_lo_6[3231:3230], regroupV0_lo_6[3223:3222]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_7 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi_3, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo_3 = {regroupV0_lo_6[3247:3246], regroupV0_lo_6[3239:3238]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi_3 = {regroupV0_lo_6[3263:3262], regroupV0_lo_6[3255:3254]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_7 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi_3, regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_hi_lo_9 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_7, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo_3 = {regroupV0_lo_6[3279:3278], regroupV0_lo_6[3271:3270]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi_3 = {regroupV0_lo_6[3295:3294], regroupV0_lo_6[3287:3286]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_7 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi_3, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo_3 = {regroupV0_lo_6[3311:3310], regroupV0_lo_6[3303:3302]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi_3 = {regroupV0_lo_6[3327:3326], regroupV0_lo_6[3319:3318]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_7 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi_3, regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_hi_hi_9 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_7, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_7};
  wire [31:0]        regroupV0_lo_hi_hi_lo_lo_hi_9 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_9, regroupV0_lo_hi_hi_lo_lo_hi_lo_9};
  wire [63:0]        regroupV0_lo_hi_hi_lo_lo_9 = {regroupV0_lo_hi_hi_lo_lo_hi_9, regroupV0_lo_hi_hi_lo_lo_lo_9};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo_3 = {regroupV0_lo_6[3343:3342], regroupV0_lo_6[3335:3334]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi_3 = {regroupV0_lo_6[3359:3358], regroupV0_lo_6[3351:3350]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_7 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi_3, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo_3 = {regroupV0_lo_6[3375:3374], regroupV0_lo_6[3367:3366]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi_3 = {regroupV0_lo_6[3391:3390], regroupV0_lo_6[3383:3382]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_7 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi_3, regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_lo_lo_9 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_7, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo_3 = {regroupV0_lo_6[3407:3406], regroupV0_lo_6[3399:3398]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi_3 = {regroupV0_lo_6[3423:3422], regroupV0_lo_6[3415:3414]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_7 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi_3, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo_3 = {regroupV0_lo_6[3439:3438], regroupV0_lo_6[3431:3430]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi_3 = {regroupV0_lo_6[3455:3454], regroupV0_lo_6[3447:3446]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_7 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi_3, regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_lo_hi_9 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_7, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_7};
  wire [31:0]        regroupV0_lo_hi_hi_lo_hi_lo_9 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_9, regroupV0_lo_hi_hi_lo_hi_lo_lo_9};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo_3 = {regroupV0_lo_6[3471:3470], regroupV0_lo_6[3463:3462]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi_3 = {regroupV0_lo_6[3487:3486], regroupV0_lo_6[3479:3478]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_7 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi_3, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo_3 = {regroupV0_lo_6[3503:3502], regroupV0_lo_6[3495:3494]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi_3 = {regroupV0_lo_6[3519:3518], regroupV0_lo_6[3511:3510]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_7 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi_3, regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_hi_lo_9 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_7, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo_3 = {regroupV0_lo_6[3535:3534], regroupV0_lo_6[3527:3526]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi_3 = {regroupV0_lo_6[3551:3550], regroupV0_lo_6[3543:3542]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_7 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi_3, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo_3 = {regroupV0_lo_6[3567:3566], regroupV0_lo_6[3559:3558]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi_3 = {regroupV0_lo_6[3583:3582], regroupV0_lo_6[3575:3574]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_7 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi_3, regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_hi_hi_9 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_7, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_7};
  wire [31:0]        regroupV0_lo_hi_hi_lo_hi_hi_9 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_9, regroupV0_lo_hi_hi_lo_hi_hi_lo_9};
  wire [63:0]        regroupV0_lo_hi_hi_lo_hi_9 = {regroupV0_lo_hi_hi_lo_hi_hi_9, regroupV0_lo_hi_hi_lo_hi_lo_9};
  wire [127:0]       regroupV0_lo_hi_hi_lo_9 = {regroupV0_lo_hi_hi_lo_hi_9, regroupV0_lo_hi_hi_lo_lo_9};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo_3 = {regroupV0_lo_6[3599:3598], regroupV0_lo_6[3591:3590]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi_3 = {regroupV0_lo_6[3615:3614], regroupV0_lo_6[3607:3606]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_7 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi_3, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo_3 = {regroupV0_lo_6[3631:3630], regroupV0_lo_6[3623:3622]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi_3 = {regroupV0_lo_6[3647:3646], regroupV0_lo_6[3639:3638]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_7 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi_3, regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_lo_lo_9 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_7, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo_3 = {regroupV0_lo_6[3663:3662], regroupV0_lo_6[3655:3654]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi_3 = {regroupV0_lo_6[3679:3678], regroupV0_lo_6[3671:3670]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_7 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi_3, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo_3 = {regroupV0_lo_6[3695:3694], regroupV0_lo_6[3687:3686]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi_3 = {regroupV0_lo_6[3711:3710], regroupV0_lo_6[3703:3702]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_7 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi_3, regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_lo_hi_9 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_7, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_7};
  wire [31:0]        regroupV0_lo_hi_hi_hi_lo_lo_9 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_9, regroupV0_lo_hi_hi_hi_lo_lo_lo_9};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo_3 = {regroupV0_lo_6[3727:3726], regroupV0_lo_6[3719:3718]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi_3 = {regroupV0_lo_6[3743:3742], regroupV0_lo_6[3735:3734]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_7 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi_3, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo_3 = {regroupV0_lo_6[3759:3758], regroupV0_lo_6[3751:3750]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi_3 = {regroupV0_lo_6[3775:3774], regroupV0_lo_6[3767:3766]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_7 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi_3, regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_hi_lo_9 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_7, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo_3 = {regroupV0_lo_6[3791:3790], regroupV0_lo_6[3783:3782]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi_3 = {regroupV0_lo_6[3807:3806], regroupV0_lo_6[3799:3798]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_7 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi_3, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo_3 = {regroupV0_lo_6[3823:3822], regroupV0_lo_6[3815:3814]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi_3 = {regroupV0_lo_6[3839:3838], regroupV0_lo_6[3831:3830]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_7 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi_3, regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_hi_hi_9 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_7, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_7};
  wire [31:0]        regroupV0_lo_hi_hi_hi_lo_hi_9 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_9, regroupV0_lo_hi_hi_hi_lo_hi_lo_9};
  wire [63:0]        regroupV0_lo_hi_hi_hi_lo_9 = {regroupV0_lo_hi_hi_hi_lo_hi_9, regroupV0_lo_hi_hi_hi_lo_lo_9};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo_3 = {regroupV0_lo_6[3855:3854], regroupV0_lo_6[3847:3846]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi_3 = {regroupV0_lo_6[3871:3870], regroupV0_lo_6[3863:3862]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_7 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi_3, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo_3 = {regroupV0_lo_6[3887:3886], regroupV0_lo_6[3879:3878]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi_3 = {regroupV0_lo_6[3903:3902], regroupV0_lo_6[3895:3894]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_7 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi_3, regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_lo_lo_9 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_7, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo_3 = {regroupV0_lo_6[3919:3918], regroupV0_lo_6[3911:3910]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi_3 = {regroupV0_lo_6[3935:3934], regroupV0_lo_6[3927:3926]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_7 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi_3, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo_3 = {regroupV0_lo_6[3951:3950], regroupV0_lo_6[3943:3942]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi_3 = {regroupV0_lo_6[3967:3966], regroupV0_lo_6[3959:3958]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_7 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi_3, regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_lo_hi_9 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_7, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_7};
  wire [31:0]        regroupV0_lo_hi_hi_hi_hi_lo_9 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_9, regroupV0_lo_hi_hi_hi_hi_lo_lo_9};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo_3 = {regroupV0_lo_6[3983:3982], regroupV0_lo_6[3975:3974]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi_3 = {regroupV0_lo_6[3999:3998], regroupV0_lo_6[3991:3990]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_7 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi_3, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo_3 = {regroupV0_lo_6[4015:4014], regroupV0_lo_6[4007:4006]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi_3 = {regroupV0_lo_6[4031:4030], regroupV0_lo_6[4023:4022]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_7 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi_3, regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_hi_lo_9 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_7, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo_3 = {regroupV0_lo_6[4047:4046], regroupV0_lo_6[4039:4038]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi_3 = {regroupV0_lo_6[4063:4062], regroupV0_lo_6[4055:4054]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_7 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi_3, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo_3 = {regroupV0_lo_6[4079:4078], regroupV0_lo_6[4071:4070]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi_3 = {regroupV0_lo_6[4095:4094], regroupV0_lo_6[4087:4086]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_7 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi_3, regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_hi_hi_9 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_7, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_7};
  wire [31:0]        regroupV0_lo_hi_hi_hi_hi_hi_9 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_9, regroupV0_lo_hi_hi_hi_hi_hi_lo_9};
  wire [63:0]        regroupV0_lo_hi_hi_hi_hi_9 = {regroupV0_lo_hi_hi_hi_hi_hi_9, regroupV0_lo_hi_hi_hi_hi_lo_9};
  wire [127:0]       regroupV0_lo_hi_hi_hi_9 = {regroupV0_lo_hi_hi_hi_hi_9, regroupV0_lo_hi_hi_hi_lo_9};
  wire [255:0]       regroupV0_lo_hi_hi_9 = {regroupV0_lo_hi_hi_hi_9, regroupV0_lo_hi_hi_lo_9};
  wire [511:0]       regroupV0_lo_hi_9 = {regroupV0_lo_hi_hi_9, regroupV0_lo_hi_lo_9};
  wire [1023:0]      regroupV0_lo_10 = {regroupV0_lo_hi_9, regroupV0_lo_lo_9};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo_3 = {regroupV0_hi_6[15:14], regroupV0_hi_6[7:6]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi_3 = {regroupV0_hi_6[31:30], regroupV0_hi_6[23:22]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_7 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo_3 = {regroupV0_hi_6[47:46], regroupV0_hi_6[39:38]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi_3 = {regroupV0_hi_6[63:62], regroupV0_hi_6[55:54]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_7 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi_3, regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_lo_lo_9 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_7, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo_3 = {regroupV0_hi_6[79:78], regroupV0_hi_6[71:70]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi_3 = {regroupV0_hi_6[95:94], regroupV0_hi_6[87:86]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_7 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi_3, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo_3 = {regroupV0_hi_6[111:110], regroupV0_hi_6[103:102]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi_3 = {regroupV0_hi_6[127:126], regroupV0_hi_6[119:118]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_7 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi_3, regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_lo_hi_9 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_7, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_7};
  wire [31:0]        regroupV0_hi_lo_lo_lo_lo_lo_9 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_9, regroupV0_hi_lo_lo_lo_lo_lo_lo_9};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo_3 = {regroupV0_hi_6[143:142], regroupV0_hi_6[135:134]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi_3 = {regroupV0_hi_6[159:158], regroupV0_hi_6[151:150]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_7 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo_3 = {regroupV0_hi_6[175:174], regroupV0_hi_6[167:166]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi_3 = {regroupV0_hi_6[191:190], regroupV0_hi_6[183:182]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_7 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi_3, regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_hi_lo_9 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_7, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo_3 = {regroupV0_hi_6[207:206], regroupV0_hi_6[199:198]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi_3 = {regroupV0_hi_6[223:222], regroupV0_hi_6[215:214]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_7 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi_3, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo_3 = {regroupV0_hi_6[239:238], regroupV0_hi_6[231:230]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi_3 = {regroupV0_hi_6[255:254], regroupV0_hi_6[247:246]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_7 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi_3, regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_hi_hi_9 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_7, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_7};
  wire [31:0]        regroupV0_hi_lo_lo_lo_lo_hi_9 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_9, regroupV0_hi_lo_lo_lo_lo_hi_lo_9};
  wire [63:0]        regroupV0_hi_lo_lo_lo_lo_9 = {regroupV0_hi_lo_lo_lo_lo_hi_9, regroupV0_hi_lo_lo_lo_lo_lo_9};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo_3 = {regroupV0_hi_6[271:270], regroupV0_hi_6[263:262]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi_3 = {regroupV0_hi_6[287:286], regroupV0_hi_6[279:278]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_7 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo_3 = {regroupV0_hi_6[303:302], regroupV0_hi_6[295:294]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi_3 = {regroupV0_hi_6[319:318], regroupV0_hi_6[311:310]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_7 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi_3, regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_lo_lo_9 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_7, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo_3 = {regroupV0_hi_6[335:334], regroupV0_hi_6[327:326]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi_3 = {regroupV0_hi_6[351:350], regroupV0_hi_6[343:342]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_7 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi_3, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo_3 = {regroupV0_hi_6[367:366], regroupV0_hi_6[359:358]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi_3 = {regroupV0_hi_6[383:382], regroupV0_hi_6[375:374]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_7 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi_3, regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_lo_hi_9 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_7, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_7};
  wire [31:0]        regroupV0_hi_lo_lo_lo_hi_lo_9 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_9, regroupV0_hi_lo_lo_lo_hi_lo_lo_9};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo_3 = {regroupV0_hi_6[399:398], regroupV0_hi_6[391:390]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi_3 = {regroupV0_hi_6[415:414], regroupV0_hi_6[407:406]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_7 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo_3 = {regroupV0_hi_6[431:430], regroupV0_hi_6[423:422]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi_3 = {regroupV0_hi_6[447:446], regroupV0_hi_6[439:438]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_7 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi_3, regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_hi_lo_9 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_7, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo_3 = {regroupV0_hi_6[463:462], regroupV0_hi_6[455:454]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi_3 = {regroupV0_hi_6[479:478], regroupV0_hi_6[471:470]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_7 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi_3, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo_3 = {regroupV0_hi_6[495:494], regroupV0_hi_6[487:486]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi_3 = {regroupV0_hi_6[511:510], regroupV0_hi_6[503:502]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_7 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi_3, regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_hi_hi_9 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_7, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_7};
  wire [31:0]        regroupV0_hi_lo_lo_lo_hi_hi_9 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_9, regroupV0_hi_lo_lo_lo_hi_hi_lo_9};
  wire [63:0]        regroupV0_hi_lo_lo_lo_hi_9 = {regroupV0_hi_lo_lo_lo_hi_hi_9, regroupV0_hi_lo_lo_lo_hi_lo_9};
  wire [127:0]       regroupV0_hi_lo_lo_lo_9 = {regroupV0_hi_lo_lo_lo_hi_9, regroupV0_hi_lo_lo_lo_lo_9};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo_3 = {regroupV0_hi_6[527:526], regroupV0_hi_6[519:518]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi_3 = {regroupV0_hi_6[543:542], regroupV0_hi_6[535:534]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_7 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi_3, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo_3 = {regroupV0_hi_6[559:558], regroupV0_hi_6[551:550]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi_3 = {regroupV0_hi_6[575:574], regroupV0_hi_6[567:566]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_7 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi_3, regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_lo_lo_9 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_7, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo_3 = {regroupV0_hi_6[591:590], regroupV0_hi_6[583:582]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi_3 = {regroupV0_hi_6[607:606], regroupV0_hi_6[599:598]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_7 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi_3, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo_3 = {regroupV0_hi_6[623:622], regroupV0_hi_6[615:614]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi_3 = {regroupV0_hi_6[639:638], regroupV0_hi_6[631:630]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_7 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi_3, regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_lo_hi_9 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_7, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_7};
  wire [31:0]        regroupV0_hi_lo_lo_hi_lo_lo_9 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_9, regroupV0_hi_lo_lo_hi_lo_lo_lo_9};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo_3 = {regroupV0_hi_6[655:654], regroupV0_hi_6[647:646]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi_3 = {regroupV0_hi_6[671:670], regroupV0_hi_6[663:662]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_7 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi_3, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo_3 = {regroupV0_hi_6[687:686], regroupV0_hi_6[679:678]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi_3 = {regroupV0_hi_6[703:702], regroupV0_hi_6[695:694]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_7 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi_3, regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_hi_lo_9 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_7, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo_3 = {regroupV0_hi_6[719:718], regroupV0_hi_6[711:710]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi_3 = {regroupV0_hi_6[735:734], regroupV0_hi_6[727:726]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_7 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi_3, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo_3 = {regroupV0_hi_6[751:750], regroupV0_hi_6[743:742]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi_3 = {regroupV0_hi_6[767:766], regroupV0_hi_6[759:758]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_7 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi_3, regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_hi_hi_9 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_7, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_7};
  wire [31:0]        regroupV0_hi_lo_lo_hi_lo_hi_9 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_9, regroupV0_hi_lo_lo_hi_lo_hi_lo_9};
  wire [63:0]        regroupV0_hi_lo_lo_hi_lo_9 = {regroupV0_hi_lo_lo_hi_lo_hi_9, regroupV0_hi_lo_lo_hi_lo_lo_9};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo_3 = {regroupV0_hi_6[783:782], regroupV0_hi_6[775:774]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi_3 = {regroupV0_hi_6[799:798], regroupV0_hi_6[791:790]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_7 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi_3, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo_3 = {regroupV0_hi_6[815:814], regroupV0_hi_6[807:806]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi_3 = {regroupV0_hi_6[831:830], regroupV0_hi_6[823:822]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_7 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi_3, regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_lo_lo_9 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_7, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo_3 = {regroupV0_hi_6[847:846], regroupV0_hi_6[839:838]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi_3 = {regroupV0_hi_6[863:862], regroupV0_hi_6[855:854]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_7 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi_3, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo_3 = {regroupV0_hi_6[879:878], regroupV0_hi_6[871:870]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi_3 = {regroupV0_hi_6[895:894], regroupV0_hi_6[887:886]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_7 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi_3, regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_lo_hi_9 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_7, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_7};
  wire [31:0]        regroupV0_hi_lo_lo_hi_hi_lo_9 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_9, regroupV0_hi_lo_lo_hi_hi_lo_lo_9};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo_3 = {regroupV0_hi_6[911:910], regroupV0_hi_6[903:902]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi_3 = {regroupV0_hi_6[927:926], regroupV0_hi_6[919:918]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_7 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi_3, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo_3 = {regroupV0_hi_6[943:942], regroupV0_hi_6[935:934]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi_3 = {regroupV0_hi_6[959:958], regroupV0_hi_6[951:950]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_7 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi_3, regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_hi_lo_9 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_7, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo_3 = {regroupV0_hi_6[975:974], regroupV0_hi_6[967:966]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi_3 = {regroupV0_hi_6[991:990], regroupV0_hi_6[983:982]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_7 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi_3, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo_3 = {regroupV0_hi_6[1007:1006], regroupV0_hi_6[999:998]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi_3 = {regroupV0_hi_6[1023:1022], regroupV0_hi_6[1015:1014]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_7 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi_3, regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_hi_hi_9 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_7, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_7};
  wire [31:0]        regroupV0_hi_lo_lo_hi_hi_hi_9 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_9, regroupV0_hi_lo_lo_hi_hi_hi_lo_9};
  wire [63:0]        regroupV0_hi_lo_lo_hi_hi_9 = {regroupV0_hi_lo_lo_hi_hi_hi_9, regroupV0_hi_lo_lo_hi_hi_lo_9};
  wire [127:0]       regroupV0_hi_lo_lo_hi_9 = {regroupV0_hi_lo_lo_hi_hi_9, regroupV0_hi_lo_lo_hi_lo_9};
  wire [255:0]       regroupV0_hi_lo_lo_9 = {regroupV0_hi_lo_lo_hi_9, regroupV0_hi_lo_lo_lo_9};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo_3 = {regroupV0_hi_6[1039:1038], regroupV0_hi_6[1031:1030]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi_3 = {regroupV0_hi_6[1055:1054], regroupV0_hi_6[1047:1046]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_7 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi_3, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo_3 = {regroupV0_hi_6[1071:1070], regroupV0_hi_6[1063:1062]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi_3 = {regroupV0_hi_6[1087:1086], regroupV0_hi_6[1079:1078]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_7 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi_3, regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_lo_lo_9 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_7, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo_3 = {regroupV0_hi_6[1103:1102], regroupV0_hi_6[1095:1094]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi_3 = {regroupV0_hi_6[1119:1118], regroupV0_hi_6[1111:1110]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_7 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi_3, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo_3 = {regroupV0_hi_6[1135:1134], regroupV0_hi_6[1127:1126]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi_3 = {regroupV0_hi_6[1151:1150], regroupV0_hi_6[1143:1142]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_7 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi_3, regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_lo_hi_9 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_7, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_7};
  wire [31:0]        regroupV0_hi_lo_hi_lo_lo_lo_9 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_9, regroupV0_hi_lo_hi_lo_lo_lo_lo_9};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo_3 = {regroupV0_hi_6[1167:1166], regroupV0_hi_6[1159:1158]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi_3 = {regroupV0_hi_6[1183:1182], regroupV0_hi_6[1175:1174]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_7 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi_3, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo_3 = {regroupV0_hi_6[1199:1198], regroupV0_hi_6[1191:1190]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi_3 = {regroupV0_hi_6[1215:1214], regroupV0_hi_6[1207:1206]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_7 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi_3, regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_hi_lo_9 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_7, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo_3 = {regroupV0_hi_6[1231:1230], regroupV0_hi_6[1223:1222]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi_3 = {regroupV0_hi_6[1247:1246], regroupV0_hi_6[1239:1238]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_7 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi_3, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo_3 = {regroupV0_hi_6[1263:1262], regroupV0_hi_6[1255:1254]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi_3 = {regroupV0_hi_6[1279:1278], regroupV0_hi_6[1271:1270]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_7 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi_3, regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_hi_hi_9 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_7, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_7};
  wire [31:0]        regroupV0_hi_lo_hi_lo_lo_hi_9 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_9, regroupV0_hi_lo_hi_lo_lo_hi_lo_9};
  wire [63:0]        regroupV0_hi_lo_hi_lo_lo_9 = {regroupV0_hi_lo_hi_lo_lo_hi_9, regroupV0_hi_lo_hi_lo_lo_lo_9};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo_3 = {regroupV0_hi_6[1295:1294], regroupV0_hi_6[1287:1286]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi_3 = {regroupV0_hi_6[1311:1310], regroupV0_hi_6[1303:1302]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_7 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi_3, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo_3 = {regroupV0_hi_6[1327:1326], regroupV0_hi_6[1319:1318]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi_3 = {regroupV0_hi_6[1343:1342], regroupV0_hi_6[1335:1334]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_7 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi_3, regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_lo_lo_9 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_7, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo_3 = {regroupV0_hi_6[1359:1358], regroupV0_hi_6[1351:1350]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi_3 = {regroupV0_hi_6[1375:1374], regroupV0_hi_6[1367:1366]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_7 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi_3, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo_3 = {regroupV0_hi_6[1391:1390], regroupV0_hi_6[1383:1382]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi_3 = {regroupV0_hi_6[1407:1406], regroupV0_hi_6[1399:1398]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_7 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi_3, regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_lo_hi_9 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_7, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_7};
  wire [31:0]        regroupV0_hi_lo_hi_lo_hi_lo_9 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_9, regroupV0_hi_lo_hi_lo_hi_lo_lo_9};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo_3 = {regroupV0_hi_6[1423:1422], regroupV0_hi_6[1415:1414]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi_3 = {regroupV0_hi_6[1439:1438], regroupV0_hi_6[1431:1430]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_7 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi_3, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo_3 = {regroupV0_hi_6[1455:1454], regroupV0_hi_6[1447:1446]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi_3 = {regroupV0_hi_6[1471:1470], regroupV0_hi_6[1463:1462]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_7 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi_3, regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_hi_lo_9 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_7, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo_3 = {regroupV0_hi_6[1487:1486], regroupV0_hi_6[1479:1478]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi_3 = {regroupV0_hi_6[1503:1502], regroupV0_hi_6[1495:1494]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_7 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi_3, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo_3 = {regroupV0_hi_6[1519:1518], regroupV0_hi_6[1511:1510]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi_3 = {regroupV0_hi_6[1535:1534], regroupV0_hi_6[1527:1526]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_7 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi_3, regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_hi_hi_9 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_7, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_7};
  wire [31:0]        regroupV0_hi_lo_hi_lo_hi_hi_9 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_9, regroupV0_hi_lo_hi_lo_hi_hi_lo_9};
  wire [63:0]        regroupV0_hi_lo_hi_lo_hi_9 = {regroupV0_hi_lo_hi_lo_hi_hi_9, regroupV0_hi_lo_hi_lo_hi_lo_9};
  wire [127:0]       regroupV0_hi_lo_hi_lo_9 = {regroupV0_hi_lo_hi_lo_hi_9, regroupV0_hi_lo_hi_lo_lo_9};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo_3 = {regroupV0_hi_6[1551:1550], regroupV0_hi_6[1543:1542]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi_3 = {regroupV0_hi_6[1567:1566], regroupV0_hi_6[1559:1558]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_7 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi_3, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo_3 = {regroupV0_hi_6[1583:1582], regroupV0_hi_6[1575:1574]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi_3 = {regroupV0_hi_6[1599:1598], regroupV0_hi_6[1591:1590]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_7 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi_3, regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_lo_lo_9 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_7, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo_3 = {regroupV0_hi_6[1615:1614], regroupV0_hi_6[1607:1606]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi_3 = {regroupV0_hi_6[1631:1630], regroupV0_hi_6[1623:1622]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_7 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi_3, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo_3 = {regroupV0_hi_6[1647:1646], regroupV0_hi_6[1639:1638]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi_3 = {regroupV0_hi_6[1663:1662], regroupV0_hi_6[1655:1654]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_7 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi_3, regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_lo_hi_9 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_7, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_7};
  wire [31:0]        regroupV0_hi_lo_hi_hi_lo_lo_9 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_9, regroupV0_hi_lo_hi_hi_lo_lo_lo_9};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo_3 = {regroupV0_hi_6[1679:1678], regroupV0_hi_6[1671:1670]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi_3 = {regroupV0_hi_6[1695:1694], regroupV0_hi_6[1687:1686]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_7 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi_3, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo_3 = {regroupV0_hi_6[1711:1710], regroupV0_hi_6[1703:1702]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi_3 = {regroupV0_hi_6[1727:1726], regroupV0_hi_6[1719:1718]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_7 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi_3, regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_hi_lo_9 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_7, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo_3 = {regroupV0_hi_6[1743:1742], regroupV0_hi_6[1735:1734]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi_3 = {regroupV0_hi_6[1759:1758], regroupV0_hi_6[1751:1750]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_7 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi_3, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo_3 = {regroupV0_hi_6[1775:1774], regroupV0_hi_6[1767:1766]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi_3 = {regroupV0_hi_6[1791:1790], regroupV0_hi_6[1783:1782]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_7 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi_3, regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_hi_hi_9 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_7, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_7};
  wire [31:0]        regroupV0_hi_lo_hi_hi_lo_hi_9 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_9, regroupV0_hi_lo_hi_hi_lo_hi_lo_9};
  wire [63:0]        regroupV0_hi_lo_hi_hi_lo_9 = {regroupV0_hi_lo_hi_hi_lo_hi_9, regroupV0_hi_lo_hi_hi_lo_lo_9};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo_3 = {regroupV0_hi_6[1807:1806], regroupV0_hi_6[1799:1798]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi_3 = {regroupV0_hi_6[1823:1822], regroupV0_hi_6[1815:1814]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_7 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi_3, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo_3 = {regroupV0_hi_6[1839:1838], regroupV0_hi_6[1831:1830]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi_3 = {regroupV0_hi_6[1855:1854], regroupV0_hi_6[1847:1846]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_7 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi_3, regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_lo_lo_9 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_7, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo_3 = {regroupV0_hi_6[1871:1870], regroupV0_hi_6[1863:1862]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi_3 = {regroupV0_hi_6[1887:1886], regroupV0_hi_6[1879:1878]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_7 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi_3, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo_3 = {regroupV0_hi_6[1903:1902], regroupV0_hi_6[1895:1894]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi_3 = {regroupV0_hi_6[1919:1918], regroupV0_hi_6[1911:1910]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_7 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi_3, regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_lo_hi_9 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_7, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_7};
  wire [31:0]        regroupV0_hi_lo_hi_hi_hi_lo_9 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_9, regroupV0_hi_lo_hi_hi_hi_lo_lo_9};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo_3 = {regroupV0_hi_6[1935:1934], regroupV0_hi_6[1927:1926]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi_3 = {regroupV0_hi_6[1951:1950], regroupV0_hi_6[1943:1942]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_7 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi_3, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo_3 = {regroupV0_hi_6[1967:1966], regroupV0_hi_6[1959:1958]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi_3 = {regroupV0_hi_6[1983:1982], regroupV0_hi_6[1975:1974]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_7 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi_3, regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_hi_lo_9 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_7, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo_3 = {regroupV0_hi_6[1999:1998], regroupV0_hi_6[1991:1990]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi_3 = {regroupV0_hi_6[2015:2014], regroupV0_hi_6[2007:2006]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_7 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi_3, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo_3 = {regroupV0_hi_6[2031:2030], regroupV0_hi_6[2023:2022]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi_3 = {regroupV0_hi_6[2047:2046], regroupV0_hi_6[2039:2038]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_7 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi_3, regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_hi_hi_9 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_7, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_7};
  wire [31:0]        regroupV0_hi_lo_hi_hi_hi_hi_9 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_9, regroupV0_hi_lo_hi_hi_hi_hi_lo_9};
  wire [63:0]        regroupV0_hi_lo_hi_hi_hi_9 = {regroupV0_hi_lo_hi_hi_hi_hi_9, regroupV0_hi_lo_hi_hi_hi_lo_9};
  wire [127:0]       regroupV0_hi_lo_hi_hi_9 = {regroupV0_hi_lo_hi_hi_hi_9, regroupV0_hi_lo_hi_hi_lo_9};
  wire [255:0]       regroupV0_hi_lo_hi_9 = {regroupV0_hi_lo_hi_hi_9, regroupV0_hi_lo_hi_lo_9};
  wire [511:0]       regroupV0_hi_lo_9 = {regroupV0_hi_lo_hi_9, regroupV0_hi_lo_lo_9};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo_3 = {regroupV0_hi_6[2063:2062], regroupV0_hi_6[2055:2054]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi_3 = {regroupV0_hi_6[2079:2078], regroupV0_hi_6[2071:2070]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_7 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi_3, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo_3 = {regroupV0_hi_6[2095:2094], regroupV0_hi_6[2087:2086]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi_3 = {regroupV0_hi_6[2111:2110], regroupV0_hi_6[2103:2102]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_7 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi_3, regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_lo_lo_9 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_7, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo_3 = {regroupV0_hi_6[2127:2126], regroupV0_hi_6[2119:2118]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi_3 = {regroupV0_hi_6[2143:2142], regroupV0_hi_6[2135:2134]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_7 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi_3, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo_3 = {regroupV0_hi_6[2159:2158], regroupV0_hi_6[2151:2150]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi_3 = {regroupV0_hi_6[2175:2174], regroupV0_hi_6[2167:2166]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_7 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi_3, regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_lo_hi_9 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_7, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_7};
  wire [31:0]        regroupV0_hi_hi_lo_lo_lo_lo_9 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_9, regroupV0_hi_hi_lo_lo_lo_lo_lo_9};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo_3 = {regroupV0_hi_6[2191:2190], regroupV0_hi_6[2183:2182]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi_3 = {regroupV0_hi_6[2207:2206], regroupV0_hi_6[2199:2198]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_7 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi_3, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo_3 = {regroupV0_hi_6[2223:2222], regroupV0_hi_6[2215:2214]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi_3 = {regroupV0_hi_6[2239:2238], regroupV0_hi_6[2231:2230]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_7 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi_3, regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_hi_lo_9 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_7, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo_3 = {regroupV0_hi_6[2255:2254], regroupV0_hi_6[2247:2246]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi_3 = {regroupV0_hi_6[2271:2270], regroupV0_hi_6[2263:2262]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_7 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi_3, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo_3 = {regroupV0_hi_6[2287:2286], regroupV0_hi_6[2279:2278]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi_3 = {regroupV0_hi_6[2303:2302], regroupV0_hi_6[2295:2294]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_7 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi_3, regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_hi_hi_9 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_7, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_7};
  wire [31:0]        regroupV0_hi_hi_lo_lo_lo_hi_9 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_9, regroupV0_hi_hi_lo_lo_lo_hi_lo_9};
  wire [63:0]        regroupV0_hi_hi_lo_lo_lo_9 = {regroupV0_hi_hi_lo_lo_lo_hi_9, regroupV0_hi_hi_lo_lo_lo_lo_9};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo_3 = {regroupV0_hi_6[2319:2318], regroupV0_hi_6[2311:2310]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi_3 = {regroupV0_hi_6[2335:2334], regroupV0_hi_6[2327:2326]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_7 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi_3, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo_3 = {regroupV0_hi_6[2351:2350], regroupV0_hi_6[2343:2342]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi_3 = {regroupV0_hi_6[2367:2366], regroupV0_hi_6[2359:2358]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_7 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi_3, regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_lo_lo_9 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_7, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo_3 = {regroupV0_hi_6[2383:2382], regroupV0_hi_6[2375:2374]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi_3 = {regroupV0_hi_6[2399:2398], regroupV0_hi_6[2391:2390]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_7 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi_3, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo_3 = {regroupV0_hi_6[2415:2414], regroupV0_hi_6[2407:2406]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi_3 = {regroupV0_hi_6[2431:2430], regroupV0_hi_6[2423:2422]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_7 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi_3, regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_lo_hi_9 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_7, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_7};
  wire [31:0]        regroupV0_hi_hi_lo_lo_hi_lo_9 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_9, regroupV0_hi_hi_lo_lo_hi_lo_lo_9};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo_3 = {regroupV0_hi_6[2447:2446], regroupV0_hi_6[2439:2438]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi_3 = {regroupV0_hi_6[2463:2462], regroupV0_hi_6[2455:2454]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_7 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi_3, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo_3 = {regroupV0_hi_6[2479:2478], regroupV0_hi_6[2471:2470]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi_3 = {regroupV0_hi_6[2495:2494], regroupV0_hi_6[2487:2486]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_7 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi_3, regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_hi_lo_9 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_7, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo_3 = {regroupV0_hi_6[2511:2510], regroupV0_hi_6[2503:2502]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi_3 = {regroupV0_hi_6[2527:2526], regroupV0_hi_6[2519:2518]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_7 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi_3, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo_3 = {regroupV0_hi_6[2543:2542], regroupV0_hi_6[2535:2534]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi_3 = {regroupV0_hi_6[2559:2558], regroupV0_hi_6[2551:2550]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_7 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi_3, regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_hi_hi_9 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_7, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_7};
  wire [31:0]        regroupV0_hi_hi_lo_lo_hi_hi_9 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_9, regroupV0_hi_hi_lo_lo_hi_hi_lo_9};
  wire [63:0]        regroupV0_hi_hi_lo_lo_hi_9 = {regroupV0_hi_hi_lo_lo_hi_hi_9, regroupV0_hi_hi_lo_lo_hi_lo_9};
  wire [127:0]       regroupV0_hi_hi_lo_lo_9 = {regroupV0_hi_hi_lo_lo_hi_9, regroupV0_hi_hi_lo_lo_lo_9};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo_3 = {regroupV0_hi_6[2575:2574], regroupV0_hi_6[2567:2566]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi_3 = {regroupV0_hi_6[2591:2590], regroupV0_hi_6[2583:2582]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_7 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi_3, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo_3 = {regroupV0_hi_6[2607:2606], regroupV0_hi_6[2599:2598]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi_3 = {regroupV0_hi_6[2623:2622], regroupV0_hi_6[2615:2614]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_7 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi_3, regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_lo_lo_9 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_7, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo_3 = {regroupV0_hi_6[2639:2638], regroupV0_hi_6[2631:2630]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi_3 = {regroupV0_hi_6[2655:2654], regroupV0_hi_6[2647:2646]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_7 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi_3, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo_3 = {regroupV0_hi_6[2671:2670], regroupV0_hi_6[2663:2662]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi_3 = {regroupV0_hi_6[2687:2686], regroupV0_hi_6[2679:2678]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_7 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi_3, regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_lo_hi_9 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_7, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_7};
  wire [31:0]        regroupV0_hi_hi_lo_hi_lo_lo_9 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_9, regroupV0_hi_hi_lo_hi_lo_lo_lo_9};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo_3 = {regroupV0_hi_6[2703:2702], regroupV0_hi_6[2695:2694]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi_3 = {regroupV0_hi_6[2719:2718], regroupV0_hi_6[2711:2710]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_7 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi_3, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo_3 = {regroupV0_hi_6[2735:2734], regroupV0_hi_6[2727:2726]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi_3 = {regroupV0_hi_6[2751:2750], regroupV0_hi_6[2743:2742]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_7 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi_3, regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_hi_lo_9 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_7, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo_3 = {regroupV0_hi_6[2767:2766], regroupV0_hi_6[2759:2758]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi_3 = {regroupV0_hi_6[2783:2782], regroupV0_hi_6[2775:2774]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_7 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi_3, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo_3 = {regroupV0_hi_6[2799:2798], regroupV0_hi_6[2791:2790]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi_3 = {regroupV0_hi_6[2815:2814], regroupV0_hi_6[2807:2806]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_7 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi_3, regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_hi_hi_9 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_7, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_7};
  wire [31:0]        regroupV0_hi_hi_lo_hi_lo_hi_9 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_9, regroupV0_hi_hi_lo_hi_lo_hi_lo_9};
  wire [63:0]        regroupV0_hi_hi_lo_hi_lo_9 = {regroupV0_hi_hi_lo_hi_lo_hi_9, regroupV0_hi_hi_lo_hi_lo_lo_9};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo_3 = {regroupV0_hi_6[2831:2830], regroupV0_hi_6[2823:2822]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi_3 = {regroupV0_hi_6[2847:2846], regroupV0_hi_6[2839:2838]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_7 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi_3, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo_3 = {regroupV0_hi_6[2863:2862], regroupV0_hi_6[2855:2854]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi_3 = {regroupV0_hi_6[2879:2878], regroupV0_hi_6[2871:2870]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_7 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi_3, regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_lo_lo_9 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_7, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo_3 = {regroupV0_hi_6[2895:2894], regroupV0_hi_6[2887:2886]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi_3 = {regroupV0_hi_6[2911:2910], regroupV0_hi_6[2903:2902]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_7 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi_3, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo_3 = {regroupV0_hi_6[2927:2926], regroupV0_hi_6[2919:2918]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi_3 = {regroupV0_hi_6[2943:2942], regroupV0_hi_6[2935:2934]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_7 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi_3, regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_lo_hi_9 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_7, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_7};
  wire [31:0]        regroupV0_hi_hi_lo_hi_hi_lo_9 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_9, regroupV0_hi_hi_lo_hi_hi_lo_lo_9};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo_3 = {regroupV0_hi_6[2959:2958], regroupV0_hi_6[2951:2950]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi_3 = {regroupV0_hi_6[2975:2974], regroupV0_hi_6[2967:2966]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_7 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi_3, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo_3 = {regroupV0_hi_6[2991:2990], regroupV0_hi_6[2983:2982]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi_3 = {regroupV0_hi_6[3007:3006], regroupV0_hi_6[2999:2998]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_7 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi_3, regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_hi_lo_9 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_7, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo_3 = {regroupV0_hi_6[3023:3022], regroupV0_hi_6[3015:3014]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi_3 = {regroupV0_hi_6[3039:3038], regroupV0_hi_6[3031:3030]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_7 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi_3, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo_3 = {regroupV0_hi_6[3055:3054], regroupV0_hi_6[3047:3046]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi_3 = {regroupV0_hi_6[3071:3070], regroupV0_hi_6[3063:3062]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_7 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi_3, regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_hi_hi_9 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_7, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_7};
  wire [31:0]        regroupV0_hi_hi_lo_hi_hi_hi_9 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_9, regroupV0_hi_hi_lo_hi_hi_hi_lo_9};
  wire [63:0]        regroupV0_hi_hi_lo_hi_hi_9 = {regroupV0_hi_hi_lo_hi_hi_hi_9, regroupV0_hi_hi_lo_hi_hi_lo_9};
  wire [127:0]       regroupV0_hi_hi_lo_hi_9 = {regroupV0_hi_hi_lo_hi_hi_9, regroupV0_hi_hi_lo_hi_lo_9};
  wire [255:0]       regroupV0_hi_hi_lo_9 = {regroupV0_hi_hi_lo_hi_9, regroupV0_hi_hi_lo_lo_9};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo_3 = {regroupV0_hi_6[3087:3086], regroupV0_hi_6[3079:3078]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi_3 = {regroupV0_hi_6[3103:3102], regroupV0_hi_6[3095:3094]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_7 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi_3, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo_3 = {regroupV0_hi_6[3119:3118], regroupV0_hi_6[3111:3110]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi_3 = {regroupV0_hi_6[3135:3134], regroupV0_hi_6[3127:3126]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_7 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi_3, regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_lo_lo_9 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_7, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo_3 = {regroupV0_hi_6[3151:3150], regroupV0_hi_6[3143:3142]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi_3 = {regroupV0_hi_6[3167:3166], regroupV0_hi_6[3159:3158]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_7 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi_3, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo_3 = {regroupV0_hi_6[3183:3182], regroupV0_hi_6[3175:3174]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi_3 = {regroupV0_hi_6[3199:3198], regroupV0_hi_6[3191:3190]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_7 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi_3, regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_lo_hi_9 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_7, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_7};
  wire [31:0]        regroupV0_hi_hi_hi_lo_lo_lo_9 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_9, regroupV0_hi_hi_hi_lo_lo_lo_lo_9};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo_3 = {regroupV0_hi_6[3215:3214], regroupV0_hi_6[3207:3206]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi_3 = {regroupV0_hi_6[3231:3230], regroupV0_hi_6[3223:3222]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_7 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi_3, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo_3 = {regroupV0_hi_6[3247:3246], regroupV0_hi_6[3239:3238]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi_3 = {regroupV0_hi_6[3263:3262], regroupV0_hi_6[3255:3254]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_7 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi_3, regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_hi_lo_9 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_7, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo_3 = {regroupV0_hi_6[3279:3278], regroupV0_hi_6[3271:3270]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi_3 = {regroupV0_hi_6[3295:3294], regroupV0_hi_6[3287:3286]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_7 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi_3, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo_3 = {regroupV0_hi_6[3311:3310], regroupV0_hi_6[3303:3302]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi_3 = {regroupV0_hi_6[3327:3326], regroupV0_hi_6[3319:3318]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_7 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_hi_hi_9 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_7, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_7};
  wire [31:0]        regroupV0_hi_hi_hi_lo_lo_hi_9 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_9, regroupV0_hi_hi_hi_lo_lo_hi_lo_9};
  wire [63:0]        regroupV0_hi_hi_hi_lo_lo_9 = {regroupV0_hi_hi_hi_lo_lo_hi_9, regroupV0_hi_hi_hi_lo_lo_lo_9};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo_3 = {regroupV0_hi_6[3343:3342], regroupV0_hi_6[3335:3334]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi_3 = {regroupV0_hi_6[3359:3358], regroupV0_hi_6[3351:3350]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_7 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi_3, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo_3 = {regroupV0_hi_6[3375:3374], regroupV0_hi_6[3367:3366]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi_3 = {regroupV0_hi_6[3391:3390], regroupV0_hi_6[3383:3382]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_7 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi_3, regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_lo_lo_9 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_7, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo_3 = {regroupV0_hi_6[3407:3406], regroupV0_hi_6[3399:3398]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi_3 = {regroupV0_hi_6[3423:3422], regroupV0_hi_6[3415:3414]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_7 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi_3, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo_3 = {regroupV0_hi_6[3439:3438], regroupV0_hi_6[3431:3430]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi_3 = {regroupV0_hi_6[3455:3454], regroupV0_hi_6[3447:3446]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_7 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi_3, regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_lo_hi_9 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_7, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_7};
  wire [31:0]        regroupV0_hi_hi_hi_lo_hi_lo_9 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_9, regroupV0_hi_hi_hi_lo_hi_lo_lo_9};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo_3 = {regroupV0_hi_6[3471:3470], regroupV0_hi_6[3463:3462]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi_3 = {regroupV0_hi_6[3487:3486], regroupV0_hi_6[3479:3478]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_7 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi_3, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo_3 = {regroupV0_hi_6[3503:3502], regroupV0_hi_6[3495:3494]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi_3 = {regroupV0_hi_6[3519:3518], regroupV0_hi_6[3511:3510]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_7 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi_3, regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_hi_lo_9 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_7, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo_3 = {regroupV0_hi_6[3535:3534], regroupV0_hi_6[3527:3526]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi_3 = {regroupV0_hi_6[3551:3550], regroupV0_hi_6[3543:3542]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_7 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi_3, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo_3 = {regroupV0_hi_6[3567:3566], regroupV0_hi_6[3559:3558]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi_3 = {regroupV0_hi_6[3583:3582], regroupV0_hi_6[3575:3574]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_7 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_hi_hi_9 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_7, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_7};
  wire [31:0]        regroupV0_hi_hi_hi_lo_hi_hi_9 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_9, regroupV0_hi_hi_hi_lo_hi_hi_lo_9};
  wire [63:0]        regroupV0_hi_hi_hi_lo_hi_9 = {regroupV0_hi_hi_hi_lo_hi_hi_9, regroupV0_hi_hi_hi_lo_hi_lo_9};
  wire [127:0]       regroupV0_hi_hi_hi_lo_9 = {regroupV0_hi_hi_hi_lo_hi_9, regroupV0_hi_hi_hi_lo_lo_9};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo_3 = {regroupV0_hi_6[3599:3598], regroupV0_hi_6[3591:3590]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi_3 = {regroupV0_hi_6[3615:3614], regroupV0_hi_6[3607:3606]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_7 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi_3, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo_3 = {regroupV0_hi_6[3631:3630], regroupV0_hi_6[3623:3622]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi_3 = {regroupV0_hi_6[3647:3646], regroupV0_hi_6[3639:3638]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_7 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi_3, regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_lo_lo_9 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_7, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo_3 = {regroupV0_hi_6[3663:3662], regroupV0_hi_6[3655:3654]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi_3 = {regroupV0_hi_6[3679:3678], regroupV0_hi_6[3671:3670]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_7 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi_3, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo_3 = {regroupV0_hi_6[3695:3694], regroupV0_hi_6[3687:3686]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi_3 = {regroupV0_hi_6[3711:3710], regroupV0_hi_6[3703:3702]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_7 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi_3, regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_lo_hi_9 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_7, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_7};
  wire [31:0]        regroupV0_hi_hi_hi_hi_lo_lo_9 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_9, regroupV0_hi_hi_hi_hi_lo_lo_lo_9};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo_3 = {regroupV0_hi_6[3727:3726], regroupV0_hi_6[3719:3718]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi_3 = {regroupV0_hi_6[3743:3742], regroupV0_hi_6[3735:3734]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_7 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi_3, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo_3 = {regroupV0_hi_6[3759:3758], regroupV0_hi_6[3751:3750]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi_3 = {regroupV0_hi_6[3775:3774], regroupV0_hi_6[3767:3766]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_7 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi_3, regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_hi_lo_9 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_7, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo_3 = {regroupV0_hi_6[3791:3790], regroupV0_hi_6[3783:3782]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi_3 = {regroupV0_hi_6[3807:3806], regroupV0_hi_6[3799:3798]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_7 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi_3, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo_3 = {regroupV0_hi_6[3823:3822], regroupV0_hi_6[3815:3814]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi_3 = {regroupV0_hi_6[3839:3838], regroupV0_hi_6[3831:3830]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_7 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_hi_hi_9 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_7, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_7};
  wire [31:0]        regroupV0_hi_hi_hi_hi_lo_hi_9 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_9, regroupV0_hi_hi_hi_hi_lo_hi_lo_9};
  wire [63:0]        regroupV0_hi_hi_hi_hi_lo_9 = {regroupV0_hi_hi_hi_hi_lo_hi_9, regroupV0_hi_hi_hi_hi_lo_lo_9};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo_3 = {regroupV0_hi_6[3855:3854], regroupV0_hi_6[3847:3846]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi_3 = {regroupV0_hi_6[3871:3870], regroupV0_hi_6[3863:3862]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_7 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi_3, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo_3 = {regroupV0_hi_6[3887:3886], regroupV0_hi_6[3879:3878]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi_3 = {regroupV0_hi_6[3903:3902], regroupV0_hi_6[3895:3894]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_7 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi_3, regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_lo_lo_9 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_7, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo_3 = {regroupV0_hi_6[3919:3918], regroupV0_hi_6[3911:3910]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi_3 = {regroupV0_hi_6[3935:3934], regroupV0_hi_6[3927:3926]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_7 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi_3, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo_3 = {regroupV0_hi_6[3951:3950], regroupV0_hi_6[3943:3942]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi_3 = {regroupV0_hi_6[3967:3966], regroupV0_hi_6[3959:3958]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_7 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi_3, regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_lo_hi_9 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_7, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_7};
  wire [31:0]        regroupV0_hi_hi_hi_hi_hi_lo_9 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_9, regroupV0_hi_hi_hi_hi_hi_lo_lo_9};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo_3 = {regroupV0_hi_6[3983:3982], regroupV0_hi_6[3975:3974]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi_3 = {regroupV0_hi_6[3999:3998], regroupV0_hi_6[3991:3990]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_7 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi_3, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo_3 = {regroupV0_hi_6[4015:4014], regroupV0_hi_6[4007:4006]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi_3 = {regroupV0_hi_6[4031:4030], regroupV0_hi_6[4023:4022]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_7 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi_3, regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_hi_lo_9 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_7, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo_3 = {regroupV0_hi_6[4047:4046], regroupV0_hi_6[4039:4038]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi_3 = {regroupV0_hi_6[4063:4062], regroupV0_hi_6[4055:4054]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_7 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi_3, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo_3 = {regroupV0_hi_6[4079:4078], regroupV0_hi_6[4071:4070]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi_3 = {regroupV0_hi_6[4095:4094], regroupV0_hi_6[4087:4086]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_7 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_hi_hi_9 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_7, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_7};
  wire [31:0]        regroupV0_hi_hi_hi_hi_hi_hi_9 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_9, regroupV0_hi_hi_hi_hi_hi_hi_lo_9};
  wire [63:0]        regroupV0_hi_hi_hi_hi_hi_9 = {regroupV0_hi_hi_hi_hi_hi_hi_9, regroupV0_hi_hi_hi_hi_hi_lo_9};
  wire [127:0]       regroupV0_hi_hi_hi_hi_9 = {regroupV0_hi_hi_hi_hi_hi_9, regroupV0_hi_hi_hi_hi_lo_9};
  wire [255:0]       regroupV0_hi_hi_hi_9 = {regroupV0_hi_hi_hi_hi_9, regroupV0_hi_hi_hi_lo_9};
  wire [511:0]       regroupV0_hi_hi_9 = {regroupV0_hi_hi_hi_9, regroupV0_hi_hi_lo_9};
  wire [1023:0]      regroupV0_hi_10 = {regroupV0_hi_hi_9, regroupV0_hi_lo_9};
  wire [4095:0]      regroupV0_lo_11 = {regroupV0_hi_8, regroupV0_lo_8, regroupV0_hi_7, regroupV0_lo_7};
  wire [4095:0]      regroupV0_hi_11 = {regroupV0_hi_10, regroupV0_lo_10, regroupV0_hi_9, regroupV0_lo_9};
  wire [8191:0]      regroupV0_1 = {regroupV0_hi_11, regroupV0_lo_11};
  wire [127:0]       regroupV0_lo_lo_lo_lo_lo_lo_10 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_10, regroupV0_lo_lo_lo_lo_lo_lo_lo_10};
  wire [127:0]       regroupV0_lo_lo_lo_lo_lo_hi_10 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_10, regroupV0_lo_lo_lo_lo_lo_hi_lo_10};
  wire [255:0]       regroupV0_lo_lo_lo_lo_lo_10 = {regroupV0_lo_lo_lo_lo_lo_hi_10, regroupV0_lo_lo_lo_lo_lo_lo_10};
  wire [127:0]       regroupV0_lo_lo_lo_lo_hi_lo_10 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_10, regroupV0_lo_lo_lo_lo_hi_lo_lo_10};
  wire [127:0]       regroupV0_lo_lo_lo_lo_hi_hi_10 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_10, regroupV0_lo_lo_lo_lo_hi_hi_lo_10};
  wire [255:0]       regroupV0_lo_lo_lo_lo_hi_10 = {regroupV0_lo_lo_lo_lo_hi_hi_10, regroupV0_lo_lo_lo_lo_hi_lo_10};
  wire [511:0]       regroupV0_lo_lo_lo_lo_10 = {regroupV0_lo_lo_lo_lo_hi_10, regroupV0_lo_lo_lo_lo_lo_10};
  wire [127:0]       regroupV0_lo_lo_lo_hi_lo_lo_10 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_10, regroupV0_lo_lo_lo_hi_lo_lo_lo_10};
  wire [127:0]       regroupV0_lo_lo_lo_hi_lo_hi_10 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_10, regroupV0_lo_lo_lo_hi_lo_hi_lo_10};
  wire [255:0]       regroupV0_lo_lo_lo_hi_lo_10 = {regroupV0_lo_lo_lo_hi_lo_hi_10, regroupV0_lo_lo_lo_hi_lo_lo_10};
  wire [127:0]       regroupV0_lo_lo_lo_hi_hi_lo_10 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_10, regroupV0_lo_lo_lo_hi_hi_lo_lo_10};
  wire [127:0]       regroupV0_lo_lo_lo_hi_hi_hi_10 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_10, regroupV0_lo_lo_lo_hi_hi_hi_lo_10};
  wire [255:0]       regroupV0_lo_lo_lo_hi_hi_10 = {regroupV0_lo_lo_lo_hi_hi_hi_10, regroupV0_lo_lo_lo_hi_hi_lo_10};
  wire [511:0]       regroupV0_lo_lo_lo_hi_10 = {regroupV0_lo_lo_lo_hi_hi_10, regroupV0_lo_lo_lo_hi_lo_10};
  wire [1023:0]      regroupV0_lo_lo_lo_10 = {regroupV0_lo_lo_lo_hi_10, regroupV0_lo_lo_lo_lo_10};
  wire [127:0]       regroupV0_lo_lo_hi_lo_lo_lo_10 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_10, regroupV0_lo_lo_hi_lo_lo_lo_lo_10};
  wire [127:0]       regroupV0_lo_lo_hi_lo_lo_hi_10 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_10, regroupV0_lo_lo_hi_lo_lo_hi_lo_10};
  wire [255:0]       regroupV0_lo_lo_hi_lo_lo_10 = {regroupV0_lo_lo_hi_lo_lo_hi_10, regroupV0_lo_lo_hi_lo_lo_lo_10};
  wire [127:0]       regroupV0_lo_lo_hi_lo_hi_lo_10 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_10, regroupV0_lo_lo_hi_lo_hi_lo_lo_10};
  wire [127:0]       regroupV0_lo_lo_hi_lo_hi_hi_10 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_10, regroupV0_lo_lo_hi_lo_hi_hi_lo_10};
  wire [255:0]       regroupV0_lo_lo_hi_lo_hi_10 = {regroupV0_lo_lo_hi_lo_hi_hi_10, regroupV0_lo_lo_hi_lo_hi_lo_10};
  wire [511:0]       regroupV0_lo_lo_hi_lo_10 = {regroupV0_lo_lo_hi_lo_hi_10, regroupV0_lo_lo_hi_lo_lo_10};
  wire [127:0]       regroupV0_lo_lo_hi_hi_lo_lo_10 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_10, regroupV0_lo_lo_hi_hi_lo_lo_lo_10};
  wire [127:0]       regroupV0_lo_lo_hi_hi_lo_hi_10 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_10, regroupV0_lo_lo_hi_hi_lo_hi_lo_10};
  wire [255:0]       regroupV0_lo_lo_hi_hi_lo_10 = {regroupV0_lo_lo_hi_hi_lo_hi_10, regroupV0_lo_lo_hi_hi_lo_lo_10};
  wire [127:0]       regroupV0_lo_lo_hi_hi_hi_lo_10 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_10, regroupV0_lo_lo_hi_hi_hi_lo_lo_10};
  wire [127:0]       regroupV0_lo_lo_hi_hi_hi_hi_10 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_10, regroupV0_lo_lo_hi_hi_hi_hi_lo_10};
  wire [255:0]       regroupV0_lo_lo_hi_hi_hi_10 = {regroupV0_lo_lo_hi_hi_hi_hi_10, regroupV0_lo_lo_hi_hi_hi_lo_10};
  wire [511:0]       regroupV0_lo_lo_hi_hi_10 = {regroupV0_lo_lo_hi_hi_hi_10, regroupV0_lo_lo_hi_hi_lo_10};
  wire [1023:0]      regroupV0_lo_lo_hi_10 = {regroupV0_lo_lo_hi_hi_10, regroupV0_lo_lo_hi_lo_10};
  wire [2047:0]      regroupV0_lo_lo_10 = {regroupV0_lo_lo_hi_10, regroupV0_lo_lo_lo_10};
  wire [127:0]       regroupV0_lo_hi_lo_lo_lo_lo_10 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_10, regroupV0_lo_hi_lo_lo_lo_lo_lo_10};
  wire [127:0]       regroupV0_lo_hi_lo_lo_lo_hi_10 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_10, regroupV0_lo_hi_lo_lo_lo_hi_lo_10};
  wire [255:0]       regroupV0_lo_hi_lo_lo_lo_10 = {regroupV0_lo_hi_lo_lo_lo_hi_10, regroupV0_lo_hi_lo_lo_lo_lo_10};
  wire [127:0]       regroupV0_lo_hi_lo_lo_hi_lo_10 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_10, regroupV0_lo_hi_lo_lo_hi_lo_lo_10};
  wire [127:0]       regroupV0_lo_hi_lo_lo_hi_hi_10 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_10, regroupV0_lo_hi_lo_lo_hi_hi_lo_10};
  wire [255:0]       regroupV0_lo_hi_lo_lo_hi_10 = {regroupV0_lo_hi_lo_lo_hi_hi_10, regroupV0_lo_hi_lo_lo_hi_lo_10};
  wire [511:0]       regroupV0_lo_hi_lo_lo_10 = {regroupV0_lo_hi_lo_lo_hi_10, regroupV0_lo_hi_lo_lo_lo_10};
  wire [127:0]       regroupV0_lo_hi_lo_hi_lo_lo_10 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_10, regroupV0_lo_hi_lo_hi_lo_lo_lo_10};
  wire [127:0]       regroupV0_lo_hi_lo_hi_lo_hi_10 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_10, regroupV0_lo_hi_lo_hi_lo_hi_lo_10};
  wire [255:0]       regroupV0_lo_hi_lo_hi_lo_10 = {regroupV0_lo_hi_lo_hi_lo_hi_10, regroupV0_lo_hi_lo_hi_lo_lo_10};
  wire [127:0]       regroupV0_lo_hi_lo_hi_hi_lo_10 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_10, regroupV0_lo_hi_lo_hi_hi_lo_lo_10};
  wire [127:0]       regroupV0_lo_hi_lo_hi_hi_hi_10 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_10, regroupV0_lo_hi_lo_hi_hi_hi_lo_10};
  wire [255:0]       regroupV0_lo_hi_lo_hi_hi_10 = {regroupV0_lo_hi_lo_hi_hi_hi_10, regroupV0_lo_hi_lo_hi_hi_lo_10};
  wire [511:0]       regroupV0_lo_hi_lo_hi_10 = {regroupV0_lo_hi_lo_hi_hi_10, regroupV0_lo_hi_lo_hi_lo_10};
  wire [1023:0]      regroupV0_lo_hi_lo_10 = {regroupV0_lo_hi_lo_hi_10, regroupV0_lo_hi_lo_lo_10};
  wire [127:0]       regroupV0_lo_hi_hi_lo_lo_lo_10 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_10, regroupV0_lo_hi_hi_lo_lo_lo_lo_10};
  wire [127:0]       regroupV0_lo_hi_hi_lo_lo_hi_10 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_10, regroupV0_lo_hi_hi_lo_lo_hi_lo_10};
  wire [255:0]       regroupV0_lo_hi_hi_lo_lo_10 = {regroupV0_lo_hi_hi_lo_lo_hi_10, regroupV0_lo_hi_hi_lo_lo_lo_10};
  wire [127:0]       regroupV0_lo_hi_hi_lo_hi_lo_10 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_10, regroupV0_lo_hi_hi_lo_hi_lo_lo_10};
  wire [127:0]       regroupV0_lo_hi_hi_lo_hi_hi_10 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_10, regroupV0_lo_hi_hi_lo_hi_hi_lo_10};
  wire [255:0]       regroupV0_lo_hi_hi_lo_hi_10 = {regroupV0_lo_hi_hi_lo_hi_hi_10, regroupV0_lo_hi_hi_lo_hi_lo_10};
  wire [511:0]       regroupV0_lo_hi_hi_lo_10 = {regroupV0_lo_hi_hi_lo_hi_10, regroupV0_lo_hi_hi_lo_lo_10};
  wire [127:0]       regroupV0_lo_hi_hi_hi_lo_lo_10 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_10, regroupV0_lo_hi_hi_hi_lo_lo_lo_10};
  wire [127:0]       regroupV0_lo_hi_hi_hi_lo_hi_10 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_10, regroupV0_lo_hi_hi_hi_lo_hi_lo_10};
  wire [255:0]       regroupV0_lo_hi_hi_hi_lo_10 = {regroupV0_lo_hi_hi_hi_lo_hi_10, regroupV0_lo_hi_hi_hi_lo_lo_10};
  wire [127:0]       regroupV0_lo_hi_hi_hi_hi_lo_10 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_10, regroupV0_lo_hi_hi_hi_hi_lo_lo_10};
  wire [127:0]       regroupV0_lo_hi_hi_hi_hi_hi_10 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_10, regroupV0_lo_hi_hi_hi_hi_hi_lo_10};
  wire [255:0]       regroupV0_lo_hi_hi_hi_hi_10 = {regroupV0_lo_hi_hi_hi_hi_hi_10, regroupV0_lo_hi_hi_hi_hi_lo_10};
  wire [511:0]       regroupV0_lo_hi_hi_hi_10 = {regroupV0_lo_hi_hi_hi_hi_10, regroupV0_lo_hi_hi_hi_lo_10};
  wire [1023:0]      regroupV0_lo_hi_hi_10 = {regroupV0_lo_hi_hi_hi_10, regroupV0_lo_hi_hi_lo_10};
  wire [2047:0]      regroupV0_lo_hi_10 = {regroupV0_lo_hi_hi_10, regroupV0_lo_hi_lo_10};
  wire [4095:0]      regroupV0_lo_12 = {regroupV0_lo_hi_10, regroupV0_lo_lo_10};
  wire [127:0]       regroupV0_hi_lo_lo_lo_lo_lo_10 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_10, regroupV0_hi_lo_lo_lo_lo_lo_lo_10};
  wire [127:0]       regroupV0_hi_lo_lo_lo_lo_hi_10 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_10, regroupV0_hi_lo_lo_lo_lo_hi_lo_10};
  wire [255:0]       regroupV0_hi_lo_lo_lo_lo_10 = {regroupV0_hi_lo_lo_lo_lo_hi_10, regroupV0_hi_lo_lo_lo_lo_lo_10};
  wire [127:0]       regroupV0_hi_lo_lo_lo_hi_lo_10 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_10, regroupV0_hi_lo_lo_lo_hi_lo_lo_10};
  wire [127:0]       regroupV0_hi_lo_lo_lo_hi_hi_10 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_10, regroupV0_hi_lo_lo_lo_hi_hi_lo_10};
  wire [255:0]       regroupV0_hi_lo_lo_lo_hi_10 = {regroupV0_hi_lo_lo_lo_hi_hi_10, regroupV0_hi_lo_lo_lo_hi_lo_10};
  wire [511:0]       regroupV0_hi_lo_lo_lo_10 = {regroupV0_hi_lo_lo_lo_hi_10, regroupV0_hi_lo_lo_lo_lo_10};
  wire [127:0]       regroupV0_hi_lo_lo_hi_lo_lo_10 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_10, regroupV0_hi_lo_lo_hi_lo_lo_lo_10};
  wire [127:0]       regroupV0_hi_lo_lo_hi_lo_hi_10 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_10, regroupV0_hi_lo_lo_hi_lo_hi_lo_10};
  wire [255:0]       regroupV0_hi_lo_lo_hi_lo_10 = {regroupV0_hi_lo_lo_hi_lo_hi_10, regroupV0_hi_lo_lo_hi_lo_lo_10};
  wire [127:0]       regroupV0_hi_lo_lo_hi_hi_lo_10 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_10, regroupV0_hi_lo_lo_hi_hi_lo_lo_10};
  wire [127:0]       regroupV0_hi_lo_lo_hi_hi_hi_10 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_10, regroupV0_hi_lo_lo_hi_hi_hi_lo_10};
  wire [255:0]       regroupV0_hi_lo_lo_hi_hi_10 = {regroupV0_hi_lo_lo_hi_hi_hi_10, regroupV0_hi_lo_lo_hi_hi_lo_10};
  wire [511:0]       regroupV0_hi_lo_lo_hi_10 = {regroupV0_hi_lo_lo_hi_hi_10, regroupV0_hi_lo_lo_hi_lo_10};
  wire [1023:0]      regroupV0_hi_lo_lo_10 = {regroupV0_hi_lo_lo_hi_10, regroupV0_hi_lo_lo_lo_10};
  wire [127:0]       regroupV0_hi_lo_hi_lo_lo_lo_10 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_10, regroupV0_hi_lo_hi_lo_lo_lo_lo_10};
  wire [127:0]       regroupV0_hi_lo_hi_lo_lo_hi_10 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_10, regroupV0_hi_lo_hi_lo_lo_hi_lo_10};
  wire [255:0]       regroupV0_hi_lo_hi_lo_lo_10 = {regroupV0_hi_lo_hi_lo_lo_hi_10, regroupV0_hi_lo_hi_lo_lo_lo_10};
  wire [127:0]       regroupV0_hi_lo_hi_lo_hi_lo_10 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_10, regroupV0_hi_lo_hi_lo_hi_lo_lo_10};
  wire [127:0]       regroupV0_hi_lo_hi_lo_hi_hi_10 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_10, regroupV0_hi_lo_hi_lo_hi_hi_lo_10};
  wire [255:0]       regroupV0_hi_lo_hi_lo_hi_10 = {regroupV0_hi_lo_hi_lo_hi_hi_10, regroupV0_hi_lo_hi_lo_hi_lo_10};
  wire [511:0]       regroupV0_hi_lo_hi_lo_10 = {regroupV0_hi_lo_hi_lo_hi_10, regroupV0_hi_lo_hi_lo_lo_10};
  wire [127:0]       regroupV0_hi_lo_hi_hi_lo_lo_10 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_10, regroupV0_hi_lo_hi_hi_lo_lo_lo_10};
  wire [127:0]       regroupV0_hi_lo_hi_hi_lo_hi_10 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_10, regroupV0_hi_lo_hi_hi_lo_hi_lo_10};
  wire [255:0]       regroupV0_hi_lo_hi_hi_lo_10 = {regroupV0_hi_lo_hi_hi_lo_hi_10, regroupV0_hi_lo_hi_hi_lo_lo_10};
  wire [127:0]       regroupV0_hi_lo_hi_hi_hi_lo_10 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_10, regroupV0_hi_lo_hi_hi_hi_lo_lo_10};
  wire [127:0]       regroupV0_hi_lo_hi_hi_hi_hi_10 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_10, regroupV0_hi_lo_hi_hi_hi_hi_lo_10};
  wire [255:0]       regroupV0_hi_lo_hi_hi_hi_10 = {regroupV0_hi_lo_hi_hi_hi_hi_10, regroupV0_hi_lo_hi_hi_hi_lo_10};
  wire [511:0]       regroupV0_hi_lo_hi_hi_10 = {regroupV0_hi_lo_hi_hi_hi_10, regroupV0_hi_lo_hi_hi_lo_10};
  wire [1023:0]      regroupV0_hi_lo_hi_10 = {regroupV0_hi_lo_hi_hi_10, regroupV0_hi_lo_hi_lo_10};
  wire [2047:0]      regroupV0_hi_lo_10 = {regroupV0_hi_lo_hi_10, regroupV0_hi_lo_lo_10};
  wire [127:0]       regroupV0_hi_hi_lo_lo_lo_lo_10 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_10, regroupV0_hi_hi_lo_lo_lo_lo_lo_10};
  wire [127:0]       regroupV0_hi_hi_lo_lo_lo_hi_10 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_10, regroupV0_hi_hi_lo_lo_lo_hi_lo_10};
  wire [255:0]       regroupV0_hi_hi_lo_lo_lo_10 = {regroupV0_hi_hi_lo_lo_lo_hi_10, regroupV0_hi_hi_lo_lo_lo_lo_10};
  wire [127:0]       regroupV0_hi_hi_lo_lo_hi_lo_10 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_10, regroupV0_hi_hi_lo_lo_hi_lo_lo_10};
  wire [127:0]       regroupV0_hi_hi_lo_lo_hi_hi_10 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_10, regroupV0_hi_hi_lo_lo_hi_hi_lo_10};
  wire [255:0]       regroupV0_hi_hi_lo_lo_hi_10 = {regroupV0_hi_hi_lo_lo_hi_hi_10, regroupV0_hi_hi_lo_lo_hi_lo_10};
  wire [511:0]       regroupV0_hi_hi_lo_lo_10 = {regroupV0_hi_hi_lo_lo_hi_10, regroupV0_hi_hi_lo_lo_lo_10};
  wire [127:0]       regroupV0_hi_hi_lo_hi_lo_lo_10 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_10, regroupV0_hi_hi_lo_hi_lo_lo_lo_10};
  wire [127:0]       regroupV0_hi_hi_lo_hi_lo_hi_10 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_10, regroupV0_hi_hi_lo_hi_lo_hi_lo_10};
  wire [255:0]       regroupV0_hi_hi_lo_hi_lo_10 = {regroupV0_hi_hi_lo_hi_lo_hi_10, regroupV0_hi_hi_lo_hi_lo_lo_10};
  wire [127:0]       regroupV0_hi_hi_lo_hi_hi_lo_10 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_10, regroupV0_hi_hi_lo_hi_hi_lo_lo_10};
  wire [127:0]       regroupV0_hi_hi_lo_hi_hi_hi_10 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_10, regroupV0_hi_hi_lo_hi_hi_hi_lo_10};
  wire [255:0]       regroupV0_hi_hi_lo_hi_hi_10 = {regroupV0_hi_hi_lo_hi_hi_hi_10, regroupV0_hi_hi_lo_hi_hi_lo_10};
  wire [511:0]       regroupV0_hi_hi_lo_hi_10 = {regroupV0_hi_hi_lo_hi_hi_10, regroupV0_hi_hi_lo_hi_lo_10};
  wire [1023:0]      regroupV0_hi_hi_lo_10 = {regroupV0_hi_hi_lo_hi_10, regroupV0_hi_hi_lo_lo_10};
  wire [127:0]       regroupV0_hi_hi_hi_lo_lo_lo_10 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_10, regroupV0_hi_hi_hi_lo_lo_lo_lo_10};
  wire [127:0]       regroupV0_hi_hi_hi_lo_lo_hi_10 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_10, regroupV0_hi_hi_hi_lo_lo_hi_lo_10};
  wire [255:0]       regroupV0_hi_hi_hi_lo_lo_10 = {regroupV0_hi_hi_hi_lo_lo_hi_10, regroupV0_hi_hi_hi_lo_lo_lo_10};
  wire [127:0]       regroupV0_hi_hi_hi_lo_hi_lo_10 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_10, regroupV0_hi_hi_hi_lo_hi_lo_lo_10};
  wire [127:0]       regroupV0_hi_hi_hi_lo_hi_hi_10 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_10, regroupV0_hi_hi_hi_lo_hi_hi_lo_10};
  wire [255:0]       regroupV0_hi_hi_hi_lo_hi_10 = {regroupV0_hi_hi_hi_lo_hi_hi_10, regroupV0_hi_hi_hi_lo_hi_lo_10};
  wire [511:0]       regroupV0_hi_hi_hi_lo_10 = {regroupV0_hi_hi_hi_lo_hi_10, regroupV0_hi_hi_hi_lo_lo_10};
  wire [127:0]       regroupV0_hi_hi_hi_hi_lo_lo_10 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_10, regroupV0_hi_hi_hi_hi_lo_lo_lo_10};
  wire [127:0]       regroupV0_hi_hi_hi_hi_lo_hi_10 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_10, regroupV0_hi_hi_hi_hi_lo_hi_lo_10};
  wire [255:0]       regroupV0_hi_hi_hi_hi_lo_10 = {regroupV0_hi_hi_hi_hi_lo_hi_10, regroupV0_hi_hi_hi_hi_lo_lo_10};
  wire [127:0]       regroupV0_hi_hi_hi_hi_hi_lo_10 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_10, regroupV0_hi_hi_hi_hi_hi_lo_lo_10};
  wire [127:0]       regroupV0_hi_hi_hi_hi_hi_hi_10 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_10, regroupV0_hi_hi_hi_hi_hi_hi_lo_10};
  wire [255:0]       regroupV0_hi_hi_hi_hi_hi_10 = {regroupV0_hi_hi_hi_hi_hi_hi_10, regroupV0_hi_hi_hi_hi_hi_lo_10};
  wire [511:0]       regroupV0_hi_hi_hi_hi_10 = {regroupV0_hi_hi_hi_hi_hi_10, regroupV0_hi_hi_hi_hi_lo_10};
  wire [1023:0]      regroupV0_hi_hi_hi_10 = {regroupV0_hi_hi_hi_hi_10, regroupV0_hi_hi_hi_lo_10};
  wire [2047:0]      regroupV0_hi_hi_10 = {regroupV0_hi_hi_hi_10, regroupV0_hi_hi_lo_10};
  wire [4095:0]      regroupV0_hi_12 = {regroupV0_hi_hi_10, regroupV0_hi_lo_10};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo_lo = {regroupV0_lo_12[4], regroupV0_lo_12[0]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo_hi = {regroupV0_lo_12[12], regroupV0_lo_12[8]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo_4 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo_hi, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi_lo = {regroupV0_lo_12[20], regroupV0_lo_12[16]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi_hi = {regroupV0_lo_12[28], regroupV0_lo_12[24]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi_4 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi_hi, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_8 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi_4, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo_lo = {regroupV0_lo_12[36], regroupV0_lo_12[32]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo_hi = {regroupV0_lo_12[44], regroupV0_lo_12[40]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo_4 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo_hi, regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi_lo = {regroupV0_lo_12[52], regroupV0_lo_12[48]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi_hi = {regroupV0_lo_12[60], regroupV0_lo_12[56]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi_4 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi_hi, regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_8 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi_4, regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_lo_lo_11 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_8, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_8};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo_lo = {regroupV0_lo_12[68], regroupV0_lo_12[64]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo_hi = {regroupV0_lo_12[76], regroupV0_lo_12[72]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo_4 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo_hi, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi_lo = {regroupV0_lo_12[84], regroupV0_lo_12[80]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi_hi = {regroupV0_lo_12[92], regroupV0_lo_12[88]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi_4 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi_hi, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_8 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi_4, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo_lo = {regroupV0_lo_12[100], regroupV0_lo_12[96]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo_hi = {regroupV0_lo_12[108], regroupV0_lo_12[104]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo_4 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo_hi, regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi_lo = {regroupV0_lo_12[116], regroupV0_lo_12[112]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi_hi = {regroupV0_lo_12[124], regroupV0_lo_12[120]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi_4 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi_hi, regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_8 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi_4, regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_lo_hi_11 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_8, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_8};
  wire [31:0]        regroupV0_lo_lo_lo_lo_lo_lo_11 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_11, regroupV0_lo_lo_lo_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo_lo = {regroupV0_lo_12[132], regroupV0_lo_12[128]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo_hi = {regroupV0_lo_12[140], regroupV0_lo_12[136]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo_4 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo_hi, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi_lo = {regroupV0_lo_12[148], regroupV0_lo_12[144]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi_hi = {regroupV0_lo_12[156], regroupV0_lo_12[152]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi_4 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi_hi, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_8 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi_4, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo_lo = {regroupV0_lo_12[164], regroupV0_lo_12[160]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo_hi = {regroupV0_lo_12[172], regroupV0_lo_12[168]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo_4 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo_hi, regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi_lo = {regroupV0_lo_12[180], regroupV0_lo_12[176]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi_hi = {regroupV0_lo_12[188], regroupV0_lo_12[184]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi_4 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi_hi, regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_8 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi_4, regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_hi_lo_11 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_8, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_8};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo_lo = {regroupV0_lo_12[196], regroupV0_lo_12[192]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo_hi = {regroupV0_lo_12[204], regroupV0_lo_12[200]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo_4 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo_hi, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi_lo = {regroupV0_lo_12[212], regroupV0_lo_12[208]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi_hi = {regroupV0_lo_12[220], regroupV0_lo_12[216]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi_4 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi_hi, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_8 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi_4, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo_lo = {regroupV0_lo_12[228], regroupV0_lo_12[224]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo_hi = {regroupV0_lo_12[236], regroupV0_lo_12[232]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo_4 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo_hi, regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi_lo = {regroupV0_lo_12[244], regroupV0_lo_12[240]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi_hi = {regroupV0_lo_12[252], regroupV0_lo_12[248]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi_4 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi_hi, regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_8 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi_4, regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_hi_hi_11 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_8, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_8};
  wire [31:0]        regroupV0_lo_lo_lo_lo_lo_hi_11 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_11, regroupV0_lo_lo_lo_lo_lo_hi_lo_11};
  wire [63:0]        regroupV0_lo_lo_lo_lo_lo_11 = {regroupV0_lo_lo_lo_lo_lo_hi_11, regroupV0_lo_lo_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo_lo = {regroupV0_lo_12[260], regroupV0_lo_12[256]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo_hi = {regroupV0_lo_12[268], regroupV0_lo_12[264]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo_4 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo_hi, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi_lo = {regroupV0_lo_12[276], regroupV0_lo_12[272]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi_hi = {regroupV0_lo_12[284], regroupV0_lo_12[280]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi_4 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi_hi, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_8 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi_4, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo_lo = {regroupV0_lo_12[292], regroupV0_lo_12[288]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo_hi = {regroupV0_lo_12[300], regroupV0_lo_12[296]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo_4 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo_hi, regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi_lo = {regroupV0_lo_12[308], regroupV0_lo_12[304]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi_hi = {regroupV0_lo_12[316], regroupV0_lo_12[312]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi_4 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi_hi, regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_8 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi_4, regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_lo_lo_11 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_8, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_8};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo_lo = {regroupV0_lo_12[324], regroupV0_lo_12[320]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo_hi = {regroupV0_lo_12[332], regroupV0_lo_12[328]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo_4 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo_hi, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi_lo = {regroupV0_lo_12[340], regroupV0_lo_12[336]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi_hi = {regroupV0_lo_12[348], regroupV0_lo_12[344]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi_4 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi_hi, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_8 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi_4, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo_lo = {regroupV0_lo_12[356], regroupV0_lo_12[352]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo_hi = {regroupV0_lo_12[364], regroupV0_lo_12[360]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo_4 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo_hi, regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi_lo = {regroupV0_lo_12[372], regroupV0_lo_12[368]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi_hi = {regroupV0_lo_12[380], regroupV0_lo_12[376]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi_4 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi_hi, regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_8 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi_4, regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_lo_hi_11 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_8, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_8};
  wire [31:0]        regroupV0_lo_lo_lo_lo_hi_lo_11 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_11, regroupV0_lo_lo_lo_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo_lo = {regroupV0_lo_12[388], regroupV0_lo_12[384]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo_hi = {regroupV0_lo_12[396], regroupV0_lo_12[392]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo_4 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo_hi, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi_lo = {regroupV0_lo_12[404], regroupV0_lo_12[400]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi_hi = {regroupV0_lo_12[412], regroupV0_lo_12[408]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi_4 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi_hi, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_8 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi_4, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo_lo = {regroupV0_lo_12[420], regroupV0_lo_12[416]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo_hi = {regroupV0_lo_12[428], regroupV0_lo_12[424]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo_4 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo_hi, regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi_lo = {regroupV0_lo_12[436], regroupV0_lo_12[432]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi_hi = {regroupV0_lo_12[444], regroupV0_lo_12[440]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi_4 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi_hi, regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_8 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi_4, regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_hi_lo_11 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_8, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_8};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo_lo = {regroupV0_lo_12[452], regroupV0_lo_12[448]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo_hi = {regroupV0_lo_12[460], regroupV0_lo_12[456]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo_4 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo_hi, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi_lo = {regroupV0_lo_12[468], regroupV0_lo_12[464]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi_hi = {regroupV0_lo_12[476], regroupV0_lo_12[472]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi_4 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi_hi, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_8 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi_4, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo_lo = {regroupV0_lo_12[484], regroupV0_lo_12[480]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo_hi = {regroupV0_lo_12[492], regroupV0_lo_12[488]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo_4 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo_hi, regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi_lo = {regroupV0_lo_12[500], regroupV0_lo_12[496]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi_hi = {regroupV0_lo_12[508], regroupV0_lo_12[504]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi_4 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi_hi, regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_8 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi_4, regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_hi_hi_11 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_8, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_8};
  wire [31:0]        regroupV0_lo_lo_lo_lo_hi_hi_11 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_11, regroupV0_lo_lo_lo_lo_hi_hi_lo_11};
  wire [63:0]        regroupV0_lo_lo_lo_lo_hi_11 = {regroupV0_lo_lo_lo_lo_hi_hi_11, regroupV0_lo_lo_lo_lo_hi_lo_11};
  wire [127:0]       regroupV0_lo_lo_lo_lo_11 = {regroupV0_lo_lo_lo_lo_hi_11, regroupV0_lo_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo_lo = {regroupV0_lo_12[516], regroupV0_lo_12[512]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo_hi = {regroupV0_lo_12[524], regroupV0_lo_12[520]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo_4 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo_hi, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi_lo = {regroupV0_lo_12[532], regroupV0_lo_12[528]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi_hi = {regroupV0_lo_12[540], regroupV0_lo_12[536]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi_4 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi_hi, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_8 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi_4, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo_lo = {regroupV0_lo_12[548], regroupV0_lo_12[544]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo_hi = {regroupV0_lo_12[556], regroupV0_lo_12[552]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo_4 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo_hi, regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi_lo = {regroupV0_lo_12[564], regroupV0_lo_12[560]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi_hi = {regroupV0_lo_12[572], regroupV0_lo_12[568]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi_4 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi_hi, regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_8 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi_4, regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_lo_lo_11 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_8, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_8};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo_lo = {regroupV0_lo_12[580], regroupV0_lo_12[576]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo_hi = {regroupV0_lo_12[588], regroupV0_lo_12[584]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo_4 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo_hi, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi_lo = {regroupV0_lo_12[596], regroupV0_lo_12[592]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi_hi = {regroupV0_lo_12[604], regroupV0_lo_12[600]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi_4 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi_hi, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_8 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi_4, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo_lo = {regroupV0_lo_12[612], regroupV0_lo_12[608]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo_hi = {regroupV0_lo_12[620], regroupV0_lo_12[616]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo_4 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo_hi, regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi_lo = {regroupV0_lo_12[628], regroupV0_lo_12[624]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi_hi = {regroupV0_lo_12[636], regroupV0_lo_12[632]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi_4 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi_hi, regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_8 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi_4, regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_lo_hi_11 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_8, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_8};
  wire [31:0]        regroupV0_lo_lo_lo_hi_lo_lo_11 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_11, regroupV0_lo_lo_lo_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo_lo = {regroupV0_lo_12[644], regroupV0_lo_12[640]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo_hi = {regroupV0_lo_12[652], regroupV0_lo_12[648]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo_4 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo_hi, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi_lo = {regroupV0_lo_12[660], regroupV0_lo_12[656]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi_hi = {regroupV0_lo_12[668], regroupV0_lo_12[664]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi_4 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi_hi, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_8 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi_4, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo_lo = {regroupV0_lo_12[676], regroupV0_lo_12[672]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo_hi = {regroupV0_lo_12[684], regroupV0_lo_12[680]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo_4 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo_hi, regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi_lo = {regroupV0_lo_12[692], regroupV0_lo_12[688]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi_hi = {regroupV0_lo_12[700], regroupV0_lo_12[696]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi_4 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi_hi, regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_8 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi_4, regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_hi_lo_11 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_8, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_8};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo_lo = {regroupV0_lo_12[708], regroupV0_lo_12[704]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo_hi = {regroupV0_lo_12[716], regroupV0_lo_12[712]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo_4 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo_hi, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi_lo = {regroupV0_lo_12[724], regroupV0_lo_12[720]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi_hi = {regroupV0_lo_12[732], regroupV0_lo_12[728]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi_4 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi_hi, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_8 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi_4, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo_lo = {regroupV0_lo_12[740], regroupV0_lo_12[736]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo_hi = {regroupV0_lo_12[748], regroupV0_lo_12[744]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo_4 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo_hi, regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi_lo = {regroupV0_lo_12[756], regroupV0_lo_12[752]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi_hi = {regroupV0_lo_12[764], regroupV0_lo_12[760]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi_4 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi_hi, regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_8 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi_4, regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_hi_hi_11 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_8, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_8};
  wire [31:0]        regroupV0_lo_lo_lo_hi_lo_hi_11 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_11, regroupV0_lo_lo_lo_hi_lo_hi_lo_11};
  wire [63:0]        regroupV0_lo_lo_lo_hi_lo_11 = {regroupV0_lo_lo_lo_hi_lo_hi_11, regroupV0_lo_lo_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo_lo = {regroupV0_lo_12[772], regroupV0_lo_12[768]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo_hi = {regroupV0_lo_12[780], regroupV0_lo_12[776]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo_4 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo_hi, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi_lo = {regroupV0_lo_12[788], regroupV0_lo_12[784]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi_hi = {regroupV0_lo_12[796], regroupV0_lo_12[792]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi_4 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi_hi, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_8 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi_4, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo_lo = {regroupV0_lo_12[804], regroupV0_lo_12[800]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo_hi = {regroupV0_lo_12[812], regroupV0_lo_12[808]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo_4 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo_hi, regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi_lo = {regroupV0_lo_12[820], regroupV0_lo_12[816]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi_hi = {regroupV0_lo_12[828], regroupV0_lo_12[824]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi_4 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi_hi, regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_8 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi_4, regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_lo_lo_11 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_8, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_8};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo_lo = {regroupV0_lo_12[836], regroupV0_lo_12[832]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo_hi = {regroupV0_lo_12[844], regroupV0_lo_12[840]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo_4 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo_hi, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi_lo = {regroupV0_lo_12[852], regroupV0_lo_12[848]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi_hi = {regroupV0_lo_12[860], regroupV0_lo_12[856]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi_4 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi_hi, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_8 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi_4, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo_lo = {regroupV0_lo_12[868], regroupV0_lo_12[864]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo_hi = {regroupV0_lo_12[876], regroupV0_lo_12[872]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo_4 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo_hi, regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi_lo = {regroupV0_lo_12[884], regroupV0_lo_12[880]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi_hi = {regroupV0_lo_12[892], regroupV0_lo_12[888]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi_4 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi_hi, regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_8 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi_4, regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_lo_hi_11 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_8, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_8};
  wire [31:0]        regroupV0_lo_lo_lo_hi_hi_lo_11 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_11, regroupV0_lo_lo_lo_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo_lo = {regroupV0_lo_12[900], regroupV0_lo_12[896]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo_hi = {regroupV0_lo_12[908], regroupV0_lo_12[904]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo_4 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo_hi, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi_lo = {regroupV0_lo_12[916], regroupV0_lo_12[912]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi_hi = {regroupV0_lo_12[924], regroupV0_lo_12[920]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi_4 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi_hi, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_8 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi_4, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo_lo = {regroupV0_lo_12[932], regroupV0_lo_12[928]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo_hi = {regroupV0_lo_12[940], regroupV0_lo_12[936]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo_4 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo_hi, regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi_lo = {regroupV0_lo_12[948], regroupV0_lo_12[944]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi_hi = {regroupV0_lo_12[956], regroupV0_lo_12[952]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi_4 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi_hi, regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_8 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi_4, regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_hi_lo_11 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_8, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_8};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo_lo = {regroupV0_lo_12[964], regroupV0_lo_12[960]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo_hi = {regroupV0_lo_12[972], regroupV0_lo_12[968]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo_4 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo_hi, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi_lo = {regroupV0_lo_12[980], regroupV0_lo_12[976]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi_hi = {regroupV0_lo_12[988], regroupV0_lo_12[984]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi_4 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi_hi, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_8 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi_4, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo_lo = {regroupV0_lo_12[996], regroupV0_lo_12[992]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo_hi = {regroupV0_lo_12[1004], regroupV0_lo_12[1000]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo_4 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo_hi, regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi_lo = {regroupV0_lo_12[1012], regroupV0_lo_12[1008]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi_hi = {regroupV0_lo_12[1020], regroupV0_lo_12[1016]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi_4 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi_hi, regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_8 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi_4, regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_hi_hi_11 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_8, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_8};
  wire [31:0]        regroupV0_lo_lo_lo_hi_hi_hi_11 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_11, regroupV0_lo_lo_lo_hi_hi_hi_lo_11};
  wire [63:0]        regroupV0_lo_lo_lo_hi_hi_11 = {regroupV0_lo_lo_lo_hi_hi_hi_11, regroupV0_lo_lo_lo_hi_hi_lo_11};
  wire [127:0]       regroupV0_lo_lo_lo_hi_11 = {regroupV0_lo_lo_lo_hi_hi_11, regroupV0_lo_lo_lo_hi_lo_11};
  wire [255:0]       regroupV0_lo_lo_lo_11 = {regroupV0_lo_lo_lo_hi_11, regroupV0_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo_lo = {regroupV0_lo_12[1028], regroupV0_lo_12[1024]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo_hi = {regroupV0_lo_12[1036], regroupV0_lo_12[1032]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo_4 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo_hi, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi_lo = {regroupV0_lo_12[1044], regroupV0_lo_12[1040]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi_hi = {regroupV0_lo_12[1052], regroupV0_lo_12[1048]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi_4 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi_hi, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_8 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi_4, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo_lo = {regroupV0_lo_12[1060], regroupV0_lo_12[1056]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo_hi = {regroupV0_lo_12[1068], regroupV0_lo_12[1064]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo_4 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo_hi, regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi_lo = {regroupV0_lo_12[1076], regroupV0_lo_12[1072]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi_hi = {regroupV0_lo_12[1084], regroupV0_lo_12[1080]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi_4 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi_hi, regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_8 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi_4, regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_lo_lo_11 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_8, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_8};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo_lo = {regroupV0_lo_12[1092], regroupV0_lo_12[1088]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo_hi = {regroupV0_lo_12[1100], regroupV0_lo_12[1096]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo_4 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo_hi, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi_lo = {regroupV0_lo_12[1108], regroupV0_lo_12[1104]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi_hi = {regroupV0_lo_12[1116], regroupV0_lo_12[1112]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi_4 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi_hi, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_8 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi_4, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo_lo = {regroupV0_lo_12[1124], regroupV0_lo_12[1120]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo_hi = {regroupV0_lo_12[1132], regroupV0_lo_12[1128]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo_4 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo_hi, regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi_lo = {regroupV0_lo_12[1140], regroupV0_lo_12[1136]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi_hi = {regroupV0_lo_12[1148], regroupV0_lo_12[1144]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi_4 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi_hi, regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_8 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi_4, regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_lo_hi_11 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_8, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_8};
  wire [31:0]        regroupV0_lo_lo_hi_lo_lo_lo_11 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_11, regroupV0_lo_lo_hi_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo_lo = {regroupV0_lo_12[1156], regroupV0_lo_12[1152]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo_hi = {regroupV0_lo_12[1164], regroupV0_lo_12[1160]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo_4 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo_hi, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi_lo = {regroupV0_lo_12[1172], regroupV0_lo_12[1168]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi_hi = {regroupV0_lo_12[1180], regroupV0_lo_12[1176]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi_4 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi_hi, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_8 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi_4, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo_lo = {regroupV0_lo_12[1188], regroupV0_lo_12[1184]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo_hi = {regroupV0_lo_12[1196], regroupV0_lo_12[1192]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo_4 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo_hi, regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi_lo = {regroupV0_lo_12[1204], regroupV0_lo_12[1200]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi_hi = {regroupV0_lo_12[1212], regroupV0_lo_12[1208]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi_4 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi_hi, regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_8 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi_4, regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_hi_lo_11 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_8, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_8};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo_lo = {regroupV0_lo_12[1220], regroupV0_lo_12[1216]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo_hi = {regroupV0_lo_12[1228], regroupV0_lo_12[1224]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo_4 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo_hi, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi_lo = {regroupV0_lo_12[1236], regroupV0_lo_12[1232]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi_hi = {regroupV0_lo_12[1244], regroupV0_lo_12[1240]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi_4 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi_hi, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_8 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi_4, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo_lo = {regroupV0_lo_12[1252], regroupV0_lo_12[1248]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo_hi = {regroupV0_lo_12[1260], regroupV0_lo_12[1256]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo_4 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo_hi, regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi_lo = {regroupV0_lo_12[1268], regroupV0_lo_12[1264]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi_hi = {regroupV0_lo_12[1276], regroupV0_lo_12[1272]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi_4 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi_hi, regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_8 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi_4, regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_hi_hi_11 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_8, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_8};
  wire [31:0]        regroupV0_lo_lo_hi_lo_lo_hi_11 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_11, regroupV0_lo_lo_hi_lo_lo_hi_lo_11};
  wire [63:0]        regroupV0_lo_lo_hi_lo_lo_11 = {regroupV0_lo_lo_hi_lo_lo_hi_11, regroupV0_lo_lo_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo_lo = {regroupV0_lo_12[1284], regroupV0_lo_12[1280]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo_hi = {regroupV0_lo_12[1292], regroupV0_lo_12[1288]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo_4 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo_hi, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi_lo = {regroupV0_lo_12[1300], regroupV0_lo_12[1296]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi_hi = {regroupV0_lo_12[1308], regroupV0_lo_12[1304]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi_4 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi_hi, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_8 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi_4, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo_lo = {regroupV0_lo_12[1316], regroupV0_lo_12[1312]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo_hi = {regroupV0_lo_12[1324], regroupV0_lo_12[1320]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo_4 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo_hi, regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi_lo = {regroupV0_lo_12[1332], regroupV0_lo_12[1328]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi_hi = {regroupV0_lo_12[1340], regroupV0_lo_12[1336]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi_4 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi_hi, regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_8 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi_4, regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_lo_lo_11 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_8, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_8};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo_lo = {regroupV0_lo_12[1348], regroupV0_lo_12[1344]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo_hi = {regroupV0_lo_12[1356], regroupV0_lo_12[1352]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo_4 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo_hi, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi_lo = {regroupV0_lo_12[1364], regroupV0_lo_12[1360]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi_hi = {regroupV0_lo_12[1372], regroupV0_lo_12[1368]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi_4 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi_hi, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_8 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi_4, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo_lo = {regroupV0_lo_12[1380], regroupV0_lo_12[1376]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo_hi = {regroupV0_lo_12[1388], regroupV0_lo_12[1384]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo_4 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo_hi, regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi_lo = {regroupV0_lo_12[1396], regroupV0_lo_12[1392]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi_hi = {regroupV0_lo_12[1404], regroupV0_lo_12[1400]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi_4 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi_hi, regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_8 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi_4, regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_lo_hi_11 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_8, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_8};
  wire [31:0]        regroupV0_lo_lo_hi_lo_hi_lo_11 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_11, regroupV0_lo_lo_hi_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo_lo = {regroupV0_lo_12[1412], regroupV0_lo_12[1408]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo_hi = {regroupV0_lo_12[1420], regroupV0_lo_12[1416]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo_4 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo_hi, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi_lo = {regroupV0_lo_12[1428], regroupV0_lo_12[1424]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi_hi = {regroupV0_lo_12[1436], regroupV0_lo_12[1432]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi_4 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi_hi, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_8 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi_4, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo_lo = {regroupV0_lo_12[1444], regroupV0_lo_12[1440]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo_hi = {regroupV0_lo_12[1452], regroupV0_lo_12[1448]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo_4 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo_hi, regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi_lo = {regroupV0_lo_12[1460], regroupV0_lo_12[1456]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi_hi = {regroupV0_lo_12[1468], regroupV0_lo_12[1464]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi_4 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi_hi, regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_8 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi_4, regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_hi_lo_11 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_8, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_8};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo_lo = {regroupV0_lo_12[1476], regroupV0_lo_12[1472]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo_hi = {regroupV0_lo_12[1484], regroupV0_lo_12[1480]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo_4 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo_hi, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi_lo = {regroupV0_lo_12[1492], regroupV0_lo_12[1488]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi_hi = {regroupV0_lo_12[1500], regroupV0_lo_12[1496]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi_4 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi_hi, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_8 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi_4, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo_lo = {regroupV0_lo_12[1508], regroupV0_lo_12[1504]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo_hi = {regroupV0_lo_12[1516], regroupV0_lo_12[1512]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo_4 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo_hi, regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi_lo = {regroupV0_lo_12[1524], regroupV0_lo_12[1520]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi_hi = {regroupV0_lo_12[1532], regroupV0_lo_12[1528]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi_4 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi_hi, regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_8 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi_4, regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_hi_hi_11 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_8, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_8};
  wire [31:0]        regroupV0_lo_lo_hi_lo_hi_hi_11 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_11, regroupV0_lo_lo_hi_lo_hi_hi_lo_11};
  wire [63:0]        regroupV0_lo_lo_hi_lo_hi_11 = {regroupV0_lo_lo_hi_lo_hi_hi_11, regroupV0_lo_lo_hi_lo_hi_lo_11};
  wire [127:0]       regroupV0_lo_lo_hi_lo_11 = {regroupV0_lo_lo_hi_lo_hi_11, regroupV0_lo_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo_lo = {regroupV0_lo_12[1540], regroupV0_lo_12[1536]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo_hi = {regroupV0_lo_12[1548], regroupV0_lo_12[1544]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo_4 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo_hi, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi_lo = {regroupV0_lo_12[1556], regroupV0_lo_12[1552]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi_hi = {regroupV0_lo_12[1564], regroupV0_lo_12[1560]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi_4 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi_hi, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_8 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi_4, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo_lo = {regroupV0_lo_12[1572], regroupV0_lo_12[1568]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo_hi = {regroupV0_lo_12[1580], regroupV0_lo_12[1576]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo_4 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo_hi, regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi_lo = {regroupV0_lo_12[1588], regroupV0_lo_12[1584]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi_hi = {regroupV0_lo_12[1596], regroupV0_lo_12[1592]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi_4 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi_hi, regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_8 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi_4, regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_lo_lo_11 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_8, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_8};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo_lo = {regroupV0_lo_12[1604], regroupV0_lo_12[1600]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo_hi = {regroupV0_lo_12[1612], regroupV0_lo_12[1608]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo_4 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo_hi, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi_lo = {regroupV0_lo_12[1620], regroupV0_lo_12[1616]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi_hi = {regroupV0_lo_12[1628], regroupV0_lo_12[1624]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi_4 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi_hi, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_8 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi_4, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo_lo = {regroupV0_lo_12[1636], regroupV0_lo_12[1632]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo_hi = {regroupV0_lo_12[1644], regroupV0_lo_12[1640]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo_4 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo_hi, regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi_lo = {regroupV0_lo_12[1652], regroupV0_lo_12[1648]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi_hi = {regroupV0_lo_12[1660], regroupV0_lo_12[1656]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi_4 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi_hi, regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_8 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi_4, regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_lo_hi_11 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_8, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_8};
  wire [31:0]        regroupV0_lo_lo_hi_hi_lo_lo_11 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_11, regroupV0_lo_lo_hi_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo_lo = {regroupV0_lo_12[1668], regroupV0_lo_12[1664]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo_hi = {regroupV0_lo_12[1676], regroupV0_lo_12[1672]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo_4 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo_hi, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi_lo = {regroupV0_lo_12[1684], regroupV0_lo_12[1680]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi_hi = {regroupV0_lo_12[1692], regroupV0_lo_12[1688]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi_4 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi_hi, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_8 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi_4, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo_lo = {regroupV0_lo_12[1700], regroupV0_lo_12[1696]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo_hi = {regroupV0_lo_12[1708], regroupV0_lo_12[1704]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo_4 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo_hi, regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi_lo = {regroupV0_lo_12[1716], regroupV0_lo_12[1712]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi_hi = {regroupV0_lo_12[1724], regroupV0_lo_12[1720]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi_4 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi_hi, regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_8 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi_4, regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_hi_lo_11 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_8, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_8};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo_lo = {regroupV0_lo_12[1732], regroupV0_lo_12[1728]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo_hi = {regroupV0_lo_12[1740], regroupV0_lo_12[1736]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo_4 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo_hi, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi_lo = {regroupV0_lo_12[1748], regroupV0_lo_12[1744]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi_hi = {regroupV0_lo_12[1756], regroupV0_lo_12[1752]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi_4 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi_hi, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_8 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi_4, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo_lo = {regroupV0_lo_12[1764], regroupV0_lo_12[1760]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo_hi = {regroupV0_lo_12[1772], regroupV0_lo_12[1768]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo_4 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo_hi, regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi_lo = {regroupV0_lo_12[1780], regroupV0_lo_12[1776]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi_hi = {regroupV0_lo_12[1788], regroupV0_lo_12[1784]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi_4 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi_hi, regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_8 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi_4, regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_hi_hi_11 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_8, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_8};
  wire [31:0]        regroupV0_lo_lo_hi_hi_lo_hi_11 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_11, regroupV0_lo_lo_hi_hi_lo_hi_lo_11};
  wire [63:0]        regroupV0_lo_lo_hi_hi_lo_11 = {regroupV0_lo_lo_hi_hi_lo_hi_11, regroupV0_lo_lo_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo_lo = {regroupV0_lo_12[1796], regroupV0_lo_12[1792]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo_hi = {regroupV0_lo_12[1804], regroupV0_lo_12[1800]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo_4 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo_hi, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi_lo = {regroupV0_lo_12[1812], regroupV0_lo_12[1808]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi_hi = {regroupV0_lo_12[1820], regroupV0_lo_12[1816]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi_4 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi_hi, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_8 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi_4, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo_lo = {regroupV0_lo_12[1828], regroupV0_lo_12[1824]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo_hi = {regroupV0_lo_12[1836], regroupV0_lo_12[1832]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo_4 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo_hi, regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi_lo = {regroupV0_lo_12[1844], regroupV0_lo_12[1840]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi_hi = {regroupV0_lo_12[1852], regroupV0_lo_12[1848]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi_4 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi_hi, regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_8 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi_4, regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_lo_lo_11 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_8, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_8};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo_lo = {regroupV0_lo_12[1860], regroupV0_lo_12[1856]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo_hi = {regroupV0_lo_12[1868], regroupV0_lo_12[1864]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo_4 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo_hi, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi_lo = {regroupV0_lo_12[1876], regroupV0_lo_12[1872]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi_hi = {regroupV0_lo_12[1884], regroupV0_lo_12[1880]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi_4 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi_hi, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_8 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi_4, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo_lo = {regroupV0_lo_12[1892], regroupV0_lo_12[1888]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo_hi = {regroupV0_lo_12[1900], regroupV0_lo_12[1896]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo_4 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo_hi, regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi_lo = {regroupV0_lo_12[1908], regroupV0_lo_12[1904]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi_hi = {regroupV0_lo_12[1916], regroupV0_lo_12[1912]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi_4 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi_hi, regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_8 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi_4, regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_lo_hi_11 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_8, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_8};
  wire [31:0]        regroupV0_lo_lo_hi_hi_hi_lo_11 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_11, regroupV0_lo_lo_hi_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo_lo = {regroupV0_lo_12[1924], regroupV0_lo_12[1920]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo_hi = {regroupV0_lo_12[1932], regroupV0_lo_12[1928]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo_4 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo_hi, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi_lo = {regroupV0_lo_12[1940], regroupV0_lo_12[1936]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi_hi = {regroupV0_lo_12[1948], regroupV0_lo_12[1944]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi_4 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi_hi, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_8 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi_4, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo_lo = {regroupV0_lo_12[1956], regroupV0_lo_12[1952]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo_hi = {regroupV0_lo_12[1964], regroupV0_lo_12[1960]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo_4 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo_hi, regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi_lo = {regroupV0_lo_12[1972], regroupV0_lo_12[1968]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi_hi = {regroupV0_lo_12[1980], regroupV0_lo_12[1976]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi_4 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi_hi, regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_8 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi_4, regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_hi_lo_11 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_8, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_8};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo_lo = {regroupV0_lo_12[1988], regroupV0_lo_12[1984]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo_hi = {regroupV0_lo_12[1996], regroupV0_lo_12[1992]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo_4 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo_hi, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi_lo = {regroupV0_lo_12[2004], regroupV0_lo_12[2000]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi_hi = {regroupV0_lo_12[2012], regroupV0_lo_12[2008]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi_4 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi_hi, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_8 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi_4, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo_lo = {regroupV0_lo_12[2020], regroupV0_lo_12[2016]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo_hi = {regroupV0_lo_12[2028], regroupV0_lo_12[2024]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo_4 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo_hi, regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi_lo = {regroupV0_lo_12[2036], regroupV0_lo_12[2032]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi_hi = {regroupV0_lo_12[2044], regroupV0_lo_12[2040]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi_4 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi_hi, regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_8 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi_4, regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_hi_hi_11 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_8, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_8};
  wire [31:0]        regroupV0_lo_lo_hi_hi_hi_hi_11 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_11, regroupV0_lo_lo_hi_hi_hi_hi_lo_11};
  wire [63:0]        regroupV0_lo_lo_hi_hi_hi_11 = {regroupV0_lo_lo_hi_hi_hi_hi_11, regroupV0_lo_lo_hi_hi_hi_lo_11};
  wire [127:0]       regroupV0_lo_lo_hi_hi_11 = {regroupV0_lo_lo_hi_hi_hi_11, regroupV0_lo_lo_hi_hi_lo_11};
  wire [255:0]       regroupV0_lo_lo_hi_11 = {regroupV0_lo_lo_hi_hi_11, regroupV0_lo_lo_hi_lo_11};
  wire [511:0]       regroupV0_lo_lo_11 = {regroupV0_lo_lo_hi_11, regroupV0_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo_lo = {regroupV0_lo_12[2052], regroupV0_lo_12[2048]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo_hi = {regroupV0_lo_12[2060], regroupV0_lo_12[2056]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo_4 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo_hi, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi_lo = {regroupV0_lo_12[2068], regroupV0_lo_12[2064]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi_hi = {regroupV0_lo_12[2076], regroupV0_lo_12[2072]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi_4 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi_hi, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_8 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi_4, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo_lo = {regroupV0_lo_12[2084], regroupV0_lo_12[2080]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo_hi = {regroupV0_lo_12[2092], regroupV0_lo_12[2088]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo_4 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo_hi, regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi_lo = {regroupV0_lo_12[2100], regroupV0_lo_12[2096]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi_hi = {regroupV0_lo_12[2108], regroupV0_lo_12[2104]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi_4 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi_hi, regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_8 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi_4, regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_lo_lo_11 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_8, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_8};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo_lo = {regroupV0_lo_12[2116], regroupV0_lo_12[2112]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo_hi = {regroupV0_lo_12[2124], regroupV0_lo_12[2120]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo_4 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo_hi, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi_lo = {regroupV0_lo_12[2132], regroupV0_lo_12[2128]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi_hi = {regroupV0_lo_12[2140], regroupV0_lo_12[2136]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi_4 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi_hi, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_8 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi_4, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo_lo = {regroupV0_lo_12[2148], regroupV0_lo_12[2144]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo_hi = {regroupV0_lo_12[2156], regroupV0_lo_12[2152]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo_4 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo_hi, regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi_lo = {regroupV0_lo_12[2164], regroupV0_lo_12[2160]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi_hi = {regroupV0_lo_12[2172], regroupV0_lo_12[2168]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi_4 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi_hi, regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_8 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi_4, regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_lo_hi_11 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_8, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_8};
  wire [31:0]        regroupV0_lo_hi_lo_lo_lo_lo_11 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_11, regroupV0_lo_hi_lo_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo_lo = {regroupV0_lo_12[2180], regroupV0_lo_12[2176]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo_hi = {regroupV0_lo_12[2188], regroupV0_lo_12[2184]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo_4 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo_hi, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi_lo = {regroupV0_lo_12[2196], regroupV0_lo_12[2192]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi_hi = {regroupV0_lo_12[2204], regroupV0_lo_12[2200]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi_4 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi_hi, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_8 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi_4, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo_lo = {regroupV0_lo_12[2212], regroupV0_lo_12[2208]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo_hi = {regroupV0_lo_12[2220], regroupV0_lo_12[2216]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo_4 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo_hi, regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi_lo = {regroupV0_lo_12[2228], regroupV0_lo_12[2224]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi_hi = {regroupV0_lo_12[2236], regroupV0_lo_12[2232]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi_4 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi_hi, regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_8 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi_4, regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_hi_lo_11 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_8, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_8};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo_lo = {regroupV0_lo_12[2244], regroupV0_lo_12[2240]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo_hi = {regroupV0_lo_12[2252], regroupV0_lo_12[2248]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo_4 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo_hi, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi_lo = {regroupV0_lo_12[2260], regroupV0_lo_12[2256]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi_hi = {regroupV0_lo_12[2268], regroupV0_lo_12[2264]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi_4 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi_hi, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_8 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi_4, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo_lo = {regroupV0_lo_12[2276], regroupV0_lo_12[2272]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo_hi = {regroupV0_lo_12[2284], regroupV0_lo_12[2280]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo_4 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo_hi, regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi_lo = {regroupV0_lo_12[2292], regroupV0_lo_12[2288]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi_hi = {regroupV0_lo_12[2300], regroupV0_lo_12[2296]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi_4 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi_hi, regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_8 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi_4, regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_hi_hi_11 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_8, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_8};
  wire [31:0]        regroupV0_lo_hi_lo_lo_lo_hi_11 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_11, regroupV0_lo_hi_lo_lo_lo_hi_lo_11};
  wire [63:0]        regroupV0_lo_hi_lo_lo_lo_11 = {regroupV0_lo_hi_lo_lo_lo_hi_11, regroupV0_lo_hi_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo_lo = {regroupV0_lo_12[2308], regroupV0_lo_12[2304]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo_hi = {regroupV0_lo_12[2316], regroupV0_lo_12[2312]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo_4 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo_hi, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi_lo = {regroupV0_lo_12[2324], regroupV0_lo_12[2320]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi_hi = {regroupV0_lo_12[2332], regroupV0_lo_12[2328]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi_4 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi_hi, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_8 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi_4, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo_lo = {regroupV0_lo_12[2340], regroupV0_lo_12[2336]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo_hi = {regroupV0_lo_12[2348], regroupV0_lo_12[2344]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo_4 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo_hi, regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi_lo = {regroupV0_lo_12[2356], regroupV0_lo_12[2352]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi_hi = {regroupV0_lo_12[2364], regroupV0_lo_12[2360]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi_4 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi_hi, regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_8 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi_4, regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_lo_lo_11 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_8, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_8};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo_lo = {regroupV0_lo_12[2372], regroupV0_lo_12[2368]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo_hi = {regroupV0_lo_12[2380], regroupV0_lo_12[2376]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo_4 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo_hi, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi_lo = {regroupV0_lo_12[2388], regroupV0_lo_12[2384]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi_hi = {regroupV0_lo_12[2396], regroupV0_lo_12[2392]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi_4 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi_hi, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_8 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi_4, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo_lo = {regroupV0_lo_12[2404], regroupV0_lo_12[2400]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo_hi = {regroupV0_lo_12[2412], regroupV0_lo_12[2408]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo_4 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo_hi, regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi_lo = {regroupV0_lo_12[2420], regroupV0_lo_12[2416]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi_hi = {regroupV0_lo_12[2428], regroupV0_lo_12[2424]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi_4 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi_hi, regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_8 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi_4, regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_lo_hi_11 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_8, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_8};
  wire [31:0]        regroupV0_lo_hi_lo_lo_hi_lo_11 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_11, regroupV0_lo_hi_lo_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo_lo = {regroupV0_lo_12[2436], regroupV0_lo_12[2432]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo_hi = {regroupV0_lo_12[2444], regroupV0_lo_12[2440]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo_4 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo_hi, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi_lo = {regroupV0_lo_12[2452], regroupV0_lo_12[2448]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi_hi = {regroupV0_lo_12[2460], regroupV0_lo_12[2456]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi_4 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi_hi, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_8 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi_4, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo_lo = {regroupV0_lo_12[2468], regroupV0_lo_12[2464]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo_hi = {regroupV0_lo_12[2476], regroupV0_lo_12[2472]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo_4 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo_hi, regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi_lo = {regroupV0_lo_12[2484], regroupV0_lo_12[2480]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi_hi = {regroupV0_lo_12[2492], regroupV0_lo_12[2488]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi_4 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi_hi, regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_8 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi_4, regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_hi_lo_11 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_8, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_8};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo_lo = {regroupV0_lo_12[2500], regroupV0_lo_12[2496]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo_hi = {regroupV0_lo_12[2508], regroupV0_lo_12[2504]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo_4 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo_hi, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi_lo = {regroupV0_lo_12[2516], regroupV0_lo_12[2512]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi_hi = {regroupV0_lo_12[2524], regroupV0_lo_12[2520]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi_4 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi_hi, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_8 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi_4, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo_lo = {regroupV0_lo_12[2532], regroupV0_lo_12[2528]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo_hi = {regroupV0_lo_12[2540], regroupV0_lo_12[2536]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo_4 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo_hi, regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi_lo = {regroupV0_lo_12[2548], regroupV0_lo_12[2544]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi_hi = {regroupV0_lo_12[2556], regroupV0_lo_12[2552]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi_4 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi_hi, regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_8 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi_4, regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_hi_hi_11 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_8, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_8};
  wire [31:0]        regroupV0_lo_hi_lo_lo_hi_hi_11 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_11, regroupV0_lo_hi_lo_lo_hi_hi_lo_11};
  wire [63:0]        regroupV0_lo_hi_lo_lo_hi_11 = {regroupV0_lo_hi_lo_lo_hi_hi_11, regroupV0_lo_hi_lo_lo_hi_lo_11};
  wire [127:0]       regroupV0_lo_hi_lo_lo_11 = {regroupV0_lo_hi_lo_lo_hi_11, regroupV0_lo_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo_lo = {regroupV0_lo_12[2564], regroupV0_lo_12[2560]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo_hi = {regroupV0_lo_12[2572], regroupV0_lo_12[2568]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo_4 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo_hi, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi_lo = {regroupV0_lo_12[2580], regroupV0_lo_12[2576]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi_hi = {regroupV0_lo_12[2588], regroupV0_lo_12[2584]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi_4 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi_hi, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_8 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi_4, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo_lo = {regroupV0_lo_12[2596], regroupV0_lo_12[2592]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo_hi = {regroupV0_lo_12[2604], regroupV0_lo_12[2600]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo_4 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo_hi, regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi_lo = {regroupV0_lo_12[2612], regroupV0_lo_12[2608]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi_hi = {regroupV0_lo_12[2620], regroupV0_lo_12[2616]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi_4 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi_hi, regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_8 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi_4, regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_lo_lo_11 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_8, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_8};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo_lo = {regroupV0_lo_12[2628], regroupV0_lo_12[2624]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo_hi = {regroupV0_lo_12[2636], regroupV0_lo_12[2632]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo_4 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo_hi, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi_lo = {regroupV0_lo_12[2644], regroupV0_lo_12[2640]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi_hi = {regroupV0_lo_12[2652], regroupV0_lo_12[2648]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi_4 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi_hi, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_8 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi_4, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo_lo = {regroupV0_lo_12[2660], regroupV0_lo_12[2656]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo_hi = {regroupV0_lo_12[2668], regroupV0_lo_12[2664]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo_4 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo_hi, regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi_lo = {regroupV0_lo_12[2676], regroupV0_lo_12[2672]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi_hi = {regroupV0_lo_12[2684], regroupV0_lo_12[2680]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi_4 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi_hi, regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_8 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi_4, regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_lo_hi_11 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_8, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_8};
  wire [31:0]        regroupV0_lo_hi_lo_hi_lo_lo_11 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_11, regroupV0_lo_hi_lo_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo_lo = {regroupV0_lo_12[2692], regroupV0_lo_12[2688]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo_hi = {regroupV0_lo_12[2700], regroupV0_lo_12[2696]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo_4 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo_hi, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi_lo = {regroupV0_lo_12[2708], regroupV0_lo_12[2704]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi_hi = {regroupV0_lo_12[2716], regroupV0_lo_12[2712]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi_4 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi_hi, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_8 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi_4, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo_lo = {regroupV0_lo_12[2724], regroupV0_lo_12[2720]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo_hi = {regroupV0_lo_12[2732], regroupV0_lo_12[2728]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo_4 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo_hi, regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi_lo = {regroupV0_lo_12[2740], regroupV0_lo_12[2736]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi_hi = {regroupV0_lo_12[2748], regroupV0_lo_12[2744]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi_4 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi_hi, regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_8 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi_4, regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_hi_lo_11 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_8, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_8};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo_lo = {regroupV0_lo_12[2756], regroupV0_lo_12[2752]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo_hi = {regroupV0_lo_12[2764], regroupV0_lo_12[2760]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo_4 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo_hi, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi_lo = {regroupV0_lo_12[2772], regroupV0_lo_12[2768]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi_hi = {regroupV0_lo_12[2780], regroupV0_lo_12[2776]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi_4 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi_hi, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_8 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi_4, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo_lo = {regroupV0_lo_12[2788], regroupV0_lo_12[2784]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo_hi = {regroupV0_lo_12[2796], regroupV0_lo_12[2792]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo_4 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo_hi, regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi_lo = {regroupV0_lo_12[2804], regroupV0_lo_12[2800]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi_hi = {regroupV0_lo_12[2812], regroupV0_lo_12[2808]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi_4 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi_hi, regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_8 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi_4, regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_hi_hi_11 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_8, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_8};
  wire [31:0]        regroupV0_lo_hi_lo_hi_lo_hi_11 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_11, regroupV0_lo_hi_lo_hi_lo_hi_lo_11};
  wire [63:0]        regroupV0_lo_hi_lo_hi_lo_11 = {regroupV0_lo_hi_lo_hi_lo_hi_11, regroupV0_lo_hi_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo_lo = {regroupV0_lo_12[2820], regroupV0_lo_12[2816]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo_hi = {regroupV0_lo_12[2828], regroupV0_lo_12[2824]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo_4 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo_hi, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi_lo = {regroupV0_lo_12[2836], regroupV0_lo_12[2832]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi_hi = {regroupV0_lo_12[2844], regroupV0_lo_12[2840]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi_4 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi_hi, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_8 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi_4, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo_lo = {regroupV0_lo_12[2852], regroupV0_lo_12[2848]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo_hi = {regroupV0_lo_12[2860], regroupV0_lo_12[2856]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo_4 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo_hi, regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi_lo = {regroupV0_lo_12[2868], regroupV0_lo_12[2864]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi_hi = {regroupV0_lo_12[2876], regroupV0_lo_12[2872]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi_4 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi_hi, regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_8 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi_4, regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_lo_lo_11 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_8, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_8};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo_lo = {regroupV0_lo_12[2884], regroupV0_lo_12[2880]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo_hi = {regroupV0_lo_12[2892], regroupV0_lo_12[2888]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo_4 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo_hi, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi_lo = {regroupV0_lo_12[2900], regroupV0_lo_12[2896]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi_hi = {regroupV0_lo_12[2908], regroupV0_lo_12[2904]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi_4 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi_hi, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_8 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi_4, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo_lo = {regroupV0_lo_12[2916], regroupV0_lo_12[2912]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo_hi = {regroupV0_lo_12[2924], regroupV0_lo_12[2920]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo_4 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo_hi, regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi_lo = {regroupV0_lo_12[2932], regroupV0_lo_12[2928]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi_hi = {regroupV0_lo_12[2940], regroupV0_lo_12[2936]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi_4 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi_hi, regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_8 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi_4, regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_lo_hi_11 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_8, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_8};
  wire [31:0]        regroupV0_lo_hi_lo_hi_hi_lo_11 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_11, regroupV0_lo_hi_lo_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo_lo = {regroupV0_lo_12[2948], regroupV0_lo_12[2944]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo_hi = {regroupV0_lo_12[2956], regroupV0_lo_12[2952]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo_4 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo_hi, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi_lo = {regroupV0_lo_12[2964], regroupV0_lo_12[2960]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi_hi = {regroupV0_lo_12[2972], regroupV0_lo_12[2968]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi_4 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi_hi, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_8 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi_4, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo_lo = {regroupV0_lo_12[2980], regroupV0_lo_12[2976]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo_hi = {regroupV0_lo_12[2988], regroupV0_lo_12[2984]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo_4 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo_hi, regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi_lo = {regroupV0_lo_12[2996], regroupV0_lo_12[2992]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi_hi = {regroupV0_lo_12[3004], regroupV0_lo_12[3000]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi_4 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi_hi, regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_8 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi_4, regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_hi_lo_11 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_8, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_8};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo_lo = {regroupV0_lo_12[3012], regroupV0_lo_12[3008]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo_hi = {regroupV0_lo_12[3020], regroupV0_lo_12[3016]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo_4 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo_hi, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi_lo = {regroupV0_lo_12[3028], regroupV0_lo_12[3024]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi_hi = {regroupV0_lo_12[3036], regroupV0_lo_12[3032]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi_4 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi_hi, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_8 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi_4, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo_lo = {regroupV0_lo_12[3044], regroupV0_lo_12[3040]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo_hi = {regroupV0_lo_12[3052], regroupV0_lo_12[3048]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo_4 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo_hi, regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi_lo = {regroupV0_lo_12[3060], regroupV0_lo_12[3056]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi_hi = {regroupV0_lo_12[3068], regroupV0_lo_12[3064]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi_4 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi_hi, regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_8 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi_4, regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_hi_hi_11 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_8, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_8};
  wire [31:0]        regroupV0_lo_hi_lo_hi_hi_hi_11 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_11, regroupV0_lo_hi_lo_hi_hi_hi_lo_11};
  wire [63:0]        regroupV0_lo_hi_lo_hi_hi_11 = {regroupV0_lo_hi_lo_hi_hi_hi_11, regroupV0_lo_hi_lo_hi_hi_lo_11};
  wire [127:0]       regroupV0_lo_hi_lo_hi_11 = {regroupV0_lo_hi_lo_hi_hi_11, regroupV0_lo_hi_lo_hi_lo_11};
  wire [255:0]       regroupV0_lo_hi_lo_11 = {regroupV0_lo_hi_lo_hi_11, regroupV0_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo_lo = {regroupV0_lo_12[3076], regroupV0_lo_12[3072]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo_hi = {regroupV0_lo_12[3084], regroupV0_lo_12[3080]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo_4 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo_hi, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi_lo = {regroupV0_lo_12[3092], regroupV0_lo_12[3088]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi_hi = {regroupV0_lo_12[3100], regroupV0_lo_12[3096]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi_4 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi_hi, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_8 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi_4, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo_lo = {regroupV0_lo_12[3108], regroupV0_lo_12[3104]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo_hi = {regroupV0_lo_12[3116], regroupV0_lo_12[3112]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo_4 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo_hi, regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi_lo = {regroupV0_lo_12[3124], regroupV0_lo_12[3120]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi_hi = {regroupV0_lo_12[3132], regroupV0_lo_12[3128]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi_4 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi_hi, regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_8 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi_4, regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_lo_lo_11 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_8, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_8};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo_lo = {regroupV0_lo_12[3140], regroupV0_lo_12[3136]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo_hi = {regroupV0_lo_12[3148], regroupV0_lo_12[3144]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo_4 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo_hi, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi_lo = {regroupV0_lo_12[3156], regroupV0_lo_12[3152]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi_hi = {regroupV0_lo_12[3164], regroupV0_lo_12[3160]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi_4 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi_hi, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_8 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi_4, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo_lo = {regroupV0_lo_12[3172], regroupV0_lo_12[3168]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo_hi = {regroupV0_lo_12[3180], regroupV0_lo_12[3176]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo_4 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo_hi, regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi_lo = {regroupV0_lo_12[3188], regroupV0_lo_12[3184]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi_hi = {regroupV0_lo_12[3196], regroupV0_lo_12[3192]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi_4 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi_hi, regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_8 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi_4, regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_lo_hi_11 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_8, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_8};
  wire [31:0]        regroupV0_lo_hi_hi_lo_lo_lo_11 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_11, regroupV0_lo_hi_hi_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo_lo = {regroupV0_lo_12[3204], regroupV0_lo_12[3200]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo_hi = {regroupV0_lo_12[3212], regroupV0_lo_12[3208]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo_4 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo_hi, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi_lo = {regroupV0_lo_12[3220], regroupV0_lo_12[3216]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi_hi = {regroupV0_lo_12[3228], regroupV0_lo_12[3224]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi_4 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi_hi, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_8 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi_4, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo_lo = {regroupV0_lo_12[3236], regroupV0_lo_12[3232]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo_hi = {regroupV0_lo_12[3244], regroupV0_lo_12[3240]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo_4 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo_hi, regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi_lo = {regroupV0_lo_12[3252], regroupV0_lo_12[3248]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi_hi = {regroupV0_lo_12[3260], regroupV0_lo_12[3256]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi_4 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi_hi, regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_8 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi_4, regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_hi_lo_11 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_8, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_8};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo_lo = {regroupV0_lo_12[3268], regroupV0_lo_12[3264]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo_hi = {regroupV0_lo_12[3276], regroupV0_lo_12[3272]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo_4 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo_hi, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi_lo = {regroupV0_lo_12[3284], regroupV0_lo_12[3280]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi_hi = {regroupV0_lo_12[3292], regroupV0_lo_12[3288]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi_4 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi_hi, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_8 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi_4, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo_lo = {regroupV0_lo_12[3300], regroupV0_lo_12[3296]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo_hi = {regroupV0_lo_12[3308], regroupV0_lo_12[3304]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo_4 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo_hi, regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi_lo = {regroupV0_lo_12[3316], regroupV0_lo_12[3312]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi_hi = {regroupV0_lo_12[3324], regroupV0_lo_12[3320]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi_4 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi_hi, regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_8 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi_4, regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_hi_hi_11 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_8, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_8};
  wire [31:0]        regroupV0_lo_hi_hi_lo_lo_hi_11 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_11, regroupV0_lo_hi_hi_lo_lo_hi_lo_11};
  wire [63:0]        regroupV0_lo_hi_hi_lo_lo_11 = {regroupV0_lo_hi_hi_lo_lo_hi_11, regroupV0_lo_hi_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo_lo = {regroupV0_lo_12[3332], regroupV0_lo_12[3328]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo_hi = {regroupV0_lo_12[3340], regroupV0_lo_12[3336]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo_4 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo_hi, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi_lo = {regroupV0_lo_12[3348], regroupV0_lo_12[3344]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi_hi = {regroupV0_lo_12[3356], regroupV0_lo_12[3352]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi_4 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi_hi, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_8 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi_4, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo_lo = {regroupV0_lo_12[3364], regroupV0_lo_12[3360]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo_hi = {regroupV0_lo_12[3372], regroupV0_lo_12[3368]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo_4 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo_hi, regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi_lo = {regroupV0_lo_12[3380], regroupV0_lo_12[3376]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi_hi = {regroupV0_lo_12[3388], regroupV0_lo_12[3384]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi_4 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi_hi, regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_8 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi_4, regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_lo_lo_11 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_8, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_8};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo_lo = {regroupV0_lo_12[3396], regroupV0_lo_12[3392]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo_hi = {regroupV0_lo_12[3404], regroupV0_lo_12[3400]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo_4 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo_hi, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi_lo = {regroupV0_lo_12[3412], regroupV0_lo_12[3408]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi_hi = {regroupV0_lo_12[3420], regroupV0_lo_12[3416]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi_4 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi_hi, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_8 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi_4, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo_lo = {regroupV0_lo_12[3428], regroupV0_lo_12[3424]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo_hi = {regroupV0_lo_12[3436], regroupV0_lo_12[3432]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo_4 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo_hi, regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi_lo = {regroupV0_lo_12[3444], regroupV0_lo_12[3440]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi_hi = {regroupV0_lo_12[3452], regroupV0_lo_12[3448]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi_4 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi_hi, regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_8 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi_4, regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_lo_hi_11 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_8, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_8};
  wire [31:0]        regroupV0_lo_hi_hi_lo_hi_lo_11 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_11, regroupV0_lo_hi_hi_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo_lo = {regroupV0_lo_12[3460], regroupV0_lo_12[3456]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo_hi = {regroupV0_lo_12[3468], regroupV0_lo_12[3464]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo_4 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo_hi, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi_lo = {regroupV0_lo_12[3476], regroupV0_lo_12[3472]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi_hi = {regroupV0_lo_12[3484], regroupV0_lo_12[3480]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi_4 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi_hi, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_8 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi_4, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo_lo = {regroupV0_lo_12[3492], regroupV0_lo_12[3488]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo_hi = {regroupV0_lo_12[3500], regroupV0_lo_12[3496]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo_4 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo_hi, regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi_lo = {regroupV0_lo_12[3508], regroupV0_lo_12[3504]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi_hi = {regroupV0_lo_12[3516], regroupV0_lo_12[3512]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi_4 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi_hi, regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_8 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi_4, regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_hi_lo_11 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_8, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_8};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo_lo = {regroupV0_lo_12[3524], regroupV0_lo_12[3520]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo_hi = {regroupV0_lo_12[3532], regroupV0_lo_12[3528]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo_4 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo_hi, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi_lo = {regroupV0_lo_12[3540], regroupV0_lo_12[3536]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi_hi = {regroupV0_lo_12[3548], regroupV0_lo_12[3544]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi_4 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi_hi, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_8 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi_4, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo_lo = {regroupV0_lo_12[3556], regroupV0_lo_12[3552]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo_hi = {regroupV0_lo_12[3564], regroupV0_lo_12[3560]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo_4 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo_hi, regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi_lo = {regroupV0_lo_12[3572], regroupV0_lo_12[3568]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi_hi = {regroupV0_lo_12[3580], regroupV0_lo_12[3576]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi_4 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi_hi, regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_8 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi_4, regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_hi_hi_11 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_8, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_8};
  wire [31:0]        regroupV0_lo_hi_hi_lo_hi_hi_11 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_11, regroupV0_lo_hi_hi_lo_hi_hi_lo_11};
  wire [63:0]        regroupV0_lo_hi_hi_lo_hi_11 = {regroupV0_lo_hi_hi_lo_hi_hi_11, regroupV0_lo_hi_hi_lo_hi_lo_11};
  wire [127:0]       regroupV0_lo_hi_hi_lo_11 = {regroupV0_lo_hi_hi_lo_hi_11, regroupV0_lo_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo_lo = {regroupV0_lo_12[3588], regroupV0_lo_12[3584]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo_hi = {regroupV0_lo_12[3596], regroupV0_lo_12[3592]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo_4 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo_hi, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi_lo = {regroupV0_lo_12[3604], regroupV0_lo_12[3600]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi_hi = {regroupV0_lo_12[3612], regroupV0_lo_12[3608]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi_4 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi_hi, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_8 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi_4, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo_lo = {regroupV0_lo_12[3620], regroupV0_lo_12[3616]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo_hi = {regroupV0_lo_12[3628], regroupV0_lo_12[3624]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo_4 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo_hi, regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi_lo = {regroupV0_lo_12[3636], regroupV0_lo_12[3632]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi_hi = {regroupV0_lo_12[3644], regroupV0_lo_12[3640]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi_4 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi_hi, regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_8 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi_4, regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_lo_lo_11 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_8, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_8};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo_lo = {regroupV0_lo_12[3652], regroupV0_lo_12[3648]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo_hi = {regroupV0_lo_12[3660], regroupV0_lo_12[3656]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo_4 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo_hi, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi_lo = {regroupV0_lo_12[3668], regroupV0_lo_12[3664]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi_hi = {regroupV0_lo_12[3676], regroupV0_lo_12[3672]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi_4 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi_hi, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_8 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi_4, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo_lo = {regroupV0_lo_12[3684], regroupV0_lo_12[3680]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo_hi = {regroupV0_lo_12[3692], regroupV0_lo_12[3688]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo_4 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo_hi, regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi_lo = {regroupV0_lo_12[3700], regroupV0_lo_12[3696]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi_hi = {regroupV0_lo_12[3708], regroupV0_lo_12[3704]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi_4 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi_hi, regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_8 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi_4, regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_lo_hi_11 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_8, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_8};
  wire [31:0]        regroupV0_lo_hi_hi_hi_lo_lo_11 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_11, regroupV0_lo_hi_hi_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo_lo = {regroupV0_lo_12[3716], regroupV0_lo_12[3712]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo_hi = {regroupV0_lo_12[3724], regroupV0_lo_12[3720]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo_4 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo_hi, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi_lo = {regroupV0_lo_12[3732], regroupV0_lo_12[3728]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi_hi = {regroupV0_lo_12[3740], regroupV0_lo_12[3736]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi_4 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi_hi, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_8 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi_4, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo_lo = {regroupV0_lo_12[3748], regroupV0_lo_12[3744]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo_hi = {regroupV0_lo_12[3756], regroupV0_lo_12[3752]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo_4 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo_hi, regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi_lo = {regroupV0_lo_12[3764], regroupV0_lo_12[3760]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi_hi = {regroupV0_lo_12[3772], regroupV0_lo_12[3768]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi_4 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi_hi, regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_8 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi_4, regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_hi_lo_11 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_8, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_8};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo_lo = {regroupV0_lo_12[3780], regroupV0_lo_12[3776]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo_hi = {regroupV0_lo_12[3788], regroupV0_lo_12[3784]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo_4 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo_hi, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi_lo = {regroupV0_lo_12[3796], regroupV0_lo_12[3792]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi_hi = {regroupV0_lo_12[3804], regroupV0_lo_12[3800]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi_4 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi_hi, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_8 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi_4, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo_lo = {regroupV0_lo_12[3812], regroupV0_lo_12[3808]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo_hi = {regroupV0_lo_12[3820], regroupV0_lo_12[3816]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo_4 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo_hi, regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi_lo = {regroupV0_lo_12[3828], regroupV0_lo_12[3824]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi_hi = {regroupV0_lo_12[3836], regroupV0_lo_12[3832]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi_4 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi_hi, regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_8 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi_4, regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_hi_hi_11 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_8, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_8};
  wire [31:0]        regroupV0_lo_hi_hi_hi_lo_hi_11 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_11, regroupV0_lo_hi_hi_hi_lo_hi_lo_11};
  wire [63:0]        regroupV0_lo_hi_hi_hi_lo_11 = {regroupV0_lo_hi_hi_hi_lo_hi_11, regroupV0_lo_hi_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo_lo = {regroupV0_lo_12[3844], regroupV0_lo_12[3840]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo_hi = {regroupV0_lo_12[3852], regroupV0_lo_12[3848]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo_4 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo_hi, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi_lo = {regroupV0_lo_12[3860], regroupV0_lo_12[3856]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi_hi = {regroupV0_lo_12[3868], regroupV0_lo_12[3864]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi_4 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi_hi, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_8 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi_4, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo_lo = {regroupV0_lo_12[3876], regroupV0_lo_12[3872]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo_hi = {regroupV0_lo_12[3884], regroupV0_lo_12[3880]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo_4 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo_hi, regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi_lo = {regroupV0_lo_12[3892], regroupV0_lo_12[3888]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi_hi = {regroupV0_lo_12[3900], regroupV0_lo_12[3896]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi_4 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi_hi, regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_8 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi_4, regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_lo_lo_11 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_8, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_8};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo_lo = {regroupV0_lo_12[3908], regroupV0_lo_12[3904]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo_hi = {regroupV0_lo_12[3916], regroupV0_lo_12[3912]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo_4 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo_hi, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi_lo = {regroupV0_lo_12[3924], regroupV0_lo_12[3920]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi_hi = {regroupV0_lo_12[3932], regroupV0_lo_12[3928]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi_4 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi_hi, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_8 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi_4, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo_lo = {regroupV0_lo_12[3940], regroupV0_lo_12[3936]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo_hi = {regroupV0_lo_12[3948], regroupV0_lo_12[3944]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo_4 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo_hi, regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi_lo = {regroupV0_lo_12[3956], regroupV0_lo_12[3952]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi_hi = {regroupV0_lo_12[3964], regroupV0_lo_12[3960]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi_4 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi_hi, regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_8 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi_4, regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_lo_hi_11 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_8, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_8};
  wire [31:0]        regroupV0_lo_hi_hi_hi_hi_lo_11 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_11, regroupV0_lo_hi_hi_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo_lo = {regroupV0_lo_12[3972], regroupV0_lo_12[3968]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo_hi = {regroupV0_lo_12[3980], regroupV0_lo_12[3976]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo_4 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo_hi, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi_lo = {regroupV0_lo_12[3988], regroupV0_lo_12[3984]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi_hi = {regroupV0_lo_12[3996], regroupV0_lo_12[3992]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi_4 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi_hi, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_8 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi_4, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo_lo = {regroupV0_lo_12[4004], regroupV0_lo_12[4000]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo_hi = {regroupV0_lo_12[4012], regroupV0_lo_12[4008]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo_4 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo_hi, regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi_lo = {regroupV0_lo_12[4020], regroupV0_lo_12[4016]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi_hi = {regroupV0_lo_12[4028], regroupV0_lo_12[4024]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi_4 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi_hi, regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_8 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi_4, regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_hi_lo_11 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_8, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_8};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo_lo = {regroupV0_lo_12[4036], regroupV0_lo_12[4032]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo_hi = {regroupV0_lo_12[4044], regroupV0_lo_12[4040]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo_4 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo_hi, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi_lo = {regroupV0_lo_12[4052], regroupV0_lo_12[4048]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi_hi = {regroupV0_lo_12[4060], regroupV0_lo_12[4056]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi_4 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi_hi, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_8 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi_4, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo_lo = {regroupV0_lo_12[4068], regroupV0_lo_12[4064]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo_hi = {regroupV0_lo_12[4076], regroupV0_lo_12[4072]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo_4 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo_hi, regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi_lo = {regroupV0_lo_12[4084], regroupV0_lo_12[4080]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi_hi = {regroupV0_lo_12[4092], regroupV0_lo_12[4088]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi_4 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi_hi, regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_8 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi_4, regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_hi_hi_11 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_8, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_8};
  wire [31:0]        regroupV0_lo_hi_hi_hi_hi_hi_11 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_11, regroupV0_lo_hi_hi_hi_hi_hi_lo_11};
  wire [63:0]        regroupV0_lo_hi_hi_hi_hi_11 = {regroupV0_lo_hi_hi_hi_hi_hi_11, regroupV0_lo_hi_hi_hi_hi_lo_11};
  wire [127:0]       regroupV0_lo_hi_hi_hi_11 = {regroupV0_lo_hi_hi_hi_hi_11, regroupV0_lo_hi_hi_hi_lo_11};
  wire [255:0]       regroupV0_lo_hi_hi_11 = {regroupV0_lo_hi_hi_hi_11, regroupV0_lo_hi_hi_lo_11};
  wire [511:0]       regroupV0_lo_hi_11 = {regroupV0_lo_hi_hi_11, regroupV0_lo_hi_lo_11};
  wire [1023:0]      regroupV0_lo_13 = {regroupV0_lo_hi_11, regroupV0_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo_lo = {regroupV0_hi_12[4], regroupV0_hi_12[0]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo_hi = {regroupV0_hi_12[12], regroupV0_hi_12[8]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo_4 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo_hi, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi_lo = {regroupV0_hi_12[20], regroupV0_hi_12[16]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi_hi = {regroupV0_hi_12[28], regroupV0_hi_12[24]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi_4 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi_hi, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_8 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi_4, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo_lo = {regroupV0_hi_12[36], regroupV0_hi_12[32]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo_hi = {regroupV0_hi_12[44], regroupV0_hi_12[40]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo_4 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo_hi, regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi_lo = {regroupV0_hi_12[52], regroupV0_hi_12[48]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi_hi = {regroupV0_hi_12[60], regroupV0_hi_12[56]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi_4 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi_hi, regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_8 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi_4, regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_lo_lo_11 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_8, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_8};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo_lo = {regroupV0_hi_12[68], regroupV0_hi_12[64]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo_hi = {regroupV0_hi_12[76], regroupV0_hi_12[72]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo_4 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo_hi, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi_lo = {regroupV0_hi_12[84], regroupV0_hi_12[80]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi_hi = {regroupV0_hi_12[92], regroupV0_hi_12[88]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi_4 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi_hi, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_8 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi_4, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo_lo = {regroupV0_hi_12[100], regroupV0_hi_12[96]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo_hi = {regroupV0_hi_12[108], regroupV0_hi_12[104]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo_4 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo_hi, regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi_lo = {regroupV0_hi_12[116], regroupV0_hi_12[112]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi_hi = {regroupV0_hi_12[124], regroupV0_hi_12[120]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi_4 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi_hi, regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_8 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi_4, regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_lo_hi_11 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_8, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_8};
  wire [31:0]        regroupV0_hi_lo_lo_lo_lo_lo_11 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_11, regroupV0_hi_lo_lo_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo_lo = {regroupV0_hi_12[132], regroupV0_hi_12[128]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo_hi = {regroupV0_hi_12[140], regroupV0_hi_12[136]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo_4 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo_hi, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi_lo = {regroupV0_hi_12[148], regroupV0_hi_12[144]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi_hi = {regroupV0_hi_12[156], regroupV0_hi_12[152]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi_4 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi_hi, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_8 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi_4, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo_lo = {regroupV0_hi_12[164], regroupV0_hi_12[160]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo_hi = {regroupV0_hi_12[172], regroupV0_hi_12[168]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo_4 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo_hi, regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi_lo = {regroupV0_hi_12[180], regroupV0_hi_12[176]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi_hi = {regroupV0_hi_12[188], regroupV0_hi_12[184]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi_4 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi_hi, regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_8 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi_4, regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_hi_lo_11 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_8, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_8};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo_lo = {regroupV0_hi_12[196], regroupV0_hi_12[192]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo_hi = {regroupV0_hi_12[204], regroupV0_hi_12[200]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo_4 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo_hi, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi_lo = {regroupV0_hi_12[212], regroupV0_hi_12[208]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi_hi = {regroupV0_hi_12[220], regroupV0_hi_12[216]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi_4 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi_hi, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_8 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi_4, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo_lo = {regroupV0_hi_12[228], regroupV0_hi_12[224]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo_hi = {regroupV0_hi_12[236], regroupV0_hi_12[232]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo_4 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo_hi, regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi_lo = {regroupV0_hi_12[244], regroupV0_hi_12[240]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi_hi = {regroupV0_hi_12[252], regroupV0_hi_12[248]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi_4 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi_hi, regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_8 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi_4, regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_hi_hi_11 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_8, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_8};
  wire [31:0]        regroupV0_hi_lo_lo_lo_lo_hi_11 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_11, regroupV0_hi_lo_lo_lo_lo_hi_lo_11};
  wire [63:0]        regroupV0_hi_lo_lo_lo_lo_11 = {regroupV0_hi_lo_lo_lo_lo_hi_11, regroupV0_hi_lo_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo_lo = {regroupV0_hi_12[260], regroupV0_hi_12[256]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo_hi = {regroupV0_hi_12[268], regroupV0_hi_12[264]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo_4 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo_hi, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi_lo = {regroupV0_hi_12[276], regroupV0_hi_12[272]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi_hi = {regroupV0_hi_12[284], regroupV0_hi_12[280]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi_4 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi_hi, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_8 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi_4, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo_lo = {regroupV0_hi_12[292], regroupV0_hi_12[288]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo_hi = {regroupV0_hi_12[300], regroupV0_hi_12[296]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo_4 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo_hi, regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi_lo = {regroupV0_hi_12[308], regroupV0_hi_12[304]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi_hi = {regroupV0_hi_12[316], regroupV0_hi_12[312]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi_4 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi_hi, regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_8 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi_4, regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_lo_lo_11 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_8, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_8};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo_lo = {regroupV0_hi_12[324], regroupV0_hi_12[320]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo_hi = {regroupV0_hi_12[332], regroupV0_hi_12[328]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo_4 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo_hi, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi_lo = {regroupV0_hi_12[340], regroupV0_hi_12[336]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi_hi = {regroupV0_hi_12[348], regroupV0_hi_12[344]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi_4 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi_hi, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_8 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi_4, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo_lo = {regroupV0_hi_12[356], regroupV0_hi_12[352]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo_hi = {regroupV0_hi_12[364], regroupV0_hi_12[360]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo_4 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo_hi, regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi_lo = {regroupV0_hi_12[372], regroupV0_hi_12[368]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi_hi = {regroupV0_hi_12[380], regroupV0_hi_12[376]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi_4 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi_hi, regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_8 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi_4, regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_lo_hi_11 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_8, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_8};
  wire [31:0]        regroupV0_hi_lo_lo_lo_hi_lo_11 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_11, regroupV0_hi_lo_lo_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo_lo = {regroupV0_hi_12[388], regroupV0_hi_12[384]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo_hi = {regroupV0_hi_12[396], regroupV0_hi_12[392]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo_4 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo_hi, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi_lo = {regroupV0_hi_12[404], regroupV0_hi_12[400]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi_hi = {regroupV0_hi_12[412], regroupV0_hi_12[408]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi_4 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi_hi, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_8 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi_4, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo_lo = {regroupV0_hi_12[420], regroupV0_hi_12[416]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo_hi = {regroupV0_hi_12[428], regroupV0_hi_12[424]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo_4 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo_hi, regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi_lo = {regroupV0_hi_12[436], regroupV0_hi_12[432]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi_hi = {regroupV0_hi_12[444], regroupV0_hi_12[440]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi_4 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi_hi, regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_8 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi_4, regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_hi_lo_11 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_8, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_8};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo_lo = {regroupV0_hi_12[452], regroupV0_hi_12[448]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo_hi = {regroupV0_hi_12[460], regroupV0_hi_12[456]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo_4 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo_hi, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi_lo = {regroupV0_hi_12[468], regroupV0_hi_12[464]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi_hi = {regroupV0_hi_12[476], regroupV0_hi_12[472]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi_4 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi_hi, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_8 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi_4, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo_lo = {regroupV0_hi_12[484], regroupV0_hi_12[480]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo_hi = {regroupV0_hi_12[492], regroupV0_hi_12[488]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo_4 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo_hi, regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi_lo = {regroupV0_hi_12[500], regroupV0_hi_12[496]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi_hi = {regroupV0_hi_12[508], regroupV0_hi_12[504]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi_4 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi_hi, regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_8 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi_4, regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_hi_hi_11 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_8, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_8};
  wire [31:0]        regroupV0_hi_lo_lo_lo_hi_hi_11 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_11, regroupV0_hi_lo_lo_lo_hi_hi_lo_11};
  wire [63:0]        regroupV0_hi_lo_lo_lo_hi_11 = {regroupV0_hi_lo_lo_lo_hi_hi_11, regroupV0_hi_lo_lo_lo_hi_lo_11};
  wire [127:0]       regroupV0_hi_lo_lo_lo_11 = {regroupV0_hi_lo_lo_lo_hi_11, regroupV0_hi_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo_lo = {regroupV0_hi_12[516], regroupV0_hi_12[512]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo_hi = {regroupV0_hi_12[524], regroupV0_hi_12[520]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo_4 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo_hi, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi_lo = {regroupV0_hi_12[532], regroupV0_hi_12[528]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi_hi = {regroupV0_hi_12[540], regroupV0_hi_12[536]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi_4 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi_hi, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_8 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi_4, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo_lo = {regroupV0_hi_12[548], regroupV0_hi_12[544]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo_hi = {regroupV0_hi_12[556], regroupV0_hi_12[552]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo_4 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo_hi, regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi_lo = {regroupV0_hi_12[564], regroupV0_hi_12[560]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi_hi = {regroupV0_hi_12[572], regroupV0_hi_12[568]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi_4 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi_hi, regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_8 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi_4, regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_lo_lo_11 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_8, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_8};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo_lo = {regroupV0_hi_12[580], regroupV0_hi_12[576]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo_hi = {regroupV0_hi_12[588], regroupV0_hi_12[584]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo_4 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo_hi, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi_lo = {regroupV0_hi_12[596], regroupV0_hi_12[592]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi_hi = {regroupV0_hi_12[604], regroupV0_hi_12[600]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi_4 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi_hi, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_8 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi_4, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo_lo = {regroupV0_hi_12[612], regroupV0_hi_12[608]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo_hi = {regroupV0_hi_12[620], regroupV0_hi_12[616]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo_4 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo_hi, regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi_lo = {regroupV0_hi_12[628], regroupV0_hi_12[624]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi_hi = {regroupV0_hi_12[636], regroupV0_hi_12[632]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi_4 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi_hi, regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_8 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi_4, regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_lo_hi_11 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_8, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_8};
  wire [31:0]        regroupV0_hi_lo_lo_hi_lo_lo_11 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_11, regroupV0_hi_lo_lo_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo_lo = {regroupV0_hi_12[644], regroupV0_hi_12[640]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo_hi = {regroupV0_hi_12[652], regroupV0_hi_12[648]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo_4 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo_hi, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi_lo = {regroupV0_hi_12[660], regroupV0_hi_12[656]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi_hi = {regroupV0_hi_12[668], regroupV0_hi_12[664]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi_4 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi_hi, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_8 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi_4, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo_lo = {regroupV0_hi_12[676], regroupV0_hi_12[672]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo_hi = {regroupV0_hi_12[684], regroupV0_hi_12[680]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo_4 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo_hi, regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi_lo = {regroupV0_hi_12[692], regroupV0_hi_12[688]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi_hi = {regroupV0_hi_12[700], regroupV0_hi_12[696]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi_4 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi_hi, regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_8 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi_4, regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_hi_lo_11 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_8, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_8};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo_lo = {regroupV0_hi_12[708], regroupV0_hi_12[704]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo_hi = {regroupV0_hi_12[716], regroupV0_hi_12[712]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo_4 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo_hi, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi_lo = {regroupV0_hi_12[724], regroupV0_hi_12[720]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi_hi = {regroupV0_hi_12[732], regroupV0_hi_12[728]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi_4 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi_hi, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_8 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi_4, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo_lo = {regroupV0_hi_12[740], regroupV0_hi_12[736]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo_hi = {regroupV0_hi_12[748], regroupV0_hi_12[744]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo_4 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo_hi, regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi_lo = {regroupV0_hi_12[756], regroupV0_hi_12[752]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi_hi = {regroupV0_hi_12[764], regroupV0_hi_12[760]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi_4 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi_hi, regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_8 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi_4, regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_hi_hi_11 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_8, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_8};
  wire [31:0]        regroupV0_hi_lo_lo_hi_lo_hi_11 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_11, regroupV0_hi_lo_lo_hi_lo_hi_lo_11};
  wire [63:0]        regroupV0_hi_lo_lo_hi_lo_11 = {regroupV0_hi_lo_lo_hi_lo_hi_11, regroupV0_hi_lo_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo_lo = {regroupV0_hi_12[772], regroupV0_hi_12[768]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo_hi = {regroupV0_hi_12[780], regroupV0_hi_12[776]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo_4 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo_hi, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi_lo = {regroupV0_hi_12[788], regroupV0_hi_12[784]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi_hi = {regroupV0_hi_12[796], regroupV0_hi_12[792]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi_4 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi_hi, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_8 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi_4, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo_lo = {regroupV0_hi_12[804], regroupV0_hi_12[800]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo_hi = {regroupV0_hi_12[812], regroupV0_hi_12[808]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo_4 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo_hi, regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi_lo = {regroupV0_hi_12[820], regroupV0_hi_12[816]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi_hi = {regroupV0_hi_12[828], regroupV0_hi_12[824]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi_4 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi_hi, regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_8 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi_4, regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_lo_lo_11 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_8, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_8};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo_lo = {regroupV0_hi_12[836], regroupV0_hi_12[832]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo_hi = {regroupV0_hi_12[844], regroupV0_hi_12[840]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo_4 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo_hi, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi_lo = {regroupV0_hi_12[852], regroupV0_hi_12[848]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi_hi = {regroupV0_hi_12[860], regroupV0_hi_12[856]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi_4 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi_hi, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_8 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi_4, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo_lo = {regroupV0_hi_12[868], regroupV0_hi_12[864]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo_hi = {regroupV0_hi_12[876], regroupV0_hi_12[872]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo_4 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo_hi, regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi_lo = {regroupV0_hi_12[884], regroupV0_hi_12[880]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi_hi = {regroupV0_hi_12[892], regroupV0_hi_12[888]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi_4 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi_hi, regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_8 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi_4, regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_lo_hi_11 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_8, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_8};
  wire [31:0]        regroupV0_hi_lo_lo_hi_hi_lo_11 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_11, regroupV0_hi_lo_lo_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo_lo = {regroupV0_hi_12[900], regroupV0_hi_12[896]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo_hi = {regroupV0_hi_12[908], regroupV0_hi_12[904]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo_4 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo_hi, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi_lo = {regroupV0_hi_12[916], regroupV0_hi_12[912]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi_hi = {regroupV0_hi_12[924], regroupV0_hi_12[920]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi_4 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi_hi, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_8 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi_4, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo_lo = {regroupV0_hi_12[932], regroupV0_hi_12[928]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo_hi = {regroupV0_hi_12[940], regroupV0_hi_12[936]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo_4 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo_hi, regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi_lo = {regroupV0_hi_12[948], regroupV0_hi_12[944]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi_hi = {regroupV0_hi_12[956], regroupV0_hi_12[952]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi_4 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi_hi, regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_8 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi_4, regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_hi_lo_11 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_8, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_8};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo_lo = {regroupV0_hi_12[964], regroupV0_hi_12[960]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo_hi = {regroupV0_hi_12[972], regroupV0_hi_12[968]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo_4 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo_hi, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi_lo = {regroupV0_hi_12[980], regroupV0_hi_12[976]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi_hi = {regroupV0_hi_12[988], regroupV0_hi_12[984]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi_4 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi_hi, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_8 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi_4, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo_lo = {regroupV0_hi_12[996], regroupV0_hi_12[992]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo_hi = {regroupV0_hi_12[1004], regroupV0_hi_12[1000]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo_4 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo_hi, regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi_lo = {regroupV0_hi_12[1012], regroupV0_hi_12[1008]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi_hi = {regroupV0_hi_12[1020], regroupV0_hi_12[1016]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi_4 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi_hi, regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_8 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi_4, regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_hi_hi_11 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_8, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_8};
  wire [31:0]        regroupV0_hi_lo_lo_hi_hi_hi_11 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_11, regroupV0_hi_lo_lo_hi_hi_hi_lo_11};
  wire [63:0]        regroupV0_hi_lo_lo_hi_hi_11 = {regroupV0_hi_lo_lo_hi_hi_hi_11, regroupV0_hi_lo_lo_hi_hi_lo_11};
  wire [127:0]       regroupV0_hi_lo_lo_hi_11 = {regroupV0_hi_lo_lo_hi_hi_11, regroupV0_hi_lo_lo_hi_lo_11};
  wire [255:0]       regroupV0_hi_lo_lo_11 = {regroupV0_hi_lo_lo_hi_11, regroupV0_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo_lo = {regroupV0_hi_12[1028], regroupV0_hi_12[1024]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo_hi = {regroupV0_hi_12[1036], regroupV0_hi_12[1032]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo_4 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo_hi, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi_lo = {regroupV0_hi_12[1044], regroupV0_hi_12[1040]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi_hi = {regroupV0_hi_12[1052], regroupV0_hi_12[1048]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi_4 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi_hi, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_8 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi_4, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo_lo = {regroupV0_hi_12[1060], regroupV0_hi_12[1056]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo_hi = {regroupV0_hi_12[1068], regroupV0_hi_12[1064]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo_4 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo_hi, regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi_lo = {regroupV0_hi_12[1076], regroupV0_hi_12[1072]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi_hi = {regroupV0_hi_12[1084], regroupV0_hi_12[1080]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi_4 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi_hi, regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_8 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi_4, regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_lo_lo_11 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_8, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_8};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo_lo = {regroupV0_hi_12[1092], regroupV0_hi_12[1088]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo_hi = {regroupV0_hi_12[1100], regroupV0_hi_12[1096]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo_4 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo_hi, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi_lo = {regroupV0_hi_12[1108], regroupV0_hi_12[1104]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi_hi = {regroupV0_hi_12[1116], regroupV0_hi_12[1112]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi_4 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi_hi, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_8 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi_4, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo_lo = {regroupV0_hi_12[1124], regroupV0_hi_12[1120]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo_hi = {regroupV0_hi_12[1132], regroupV0_hi_12[1128]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo_4 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo_hi, regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi_lo = {regroupV0_hi_12[1140], regroupV0_hi_12[1136]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi_hi = {regroupV0_hi_12[1148], regroupV0_hi_12[1144]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi_4 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi_hi, regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_8 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi_4, regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_lo_hi_11 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_8, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_8};
  wire [31:0]        regroupV0_hi_lo_hi_lo_lo_lo_11 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_11, regroupV0_hi_lo_hi_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo_lo = {regroupV0_hi_12[1156], regroupV0_hi_12[1152]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo_hi = {regroupV0_hi_12[1164], regroupV0_hi_12[1160]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo_4 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo_hi, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi_lo = {regroupV0_hi_12[1172], regroupV0_hi_12[1168]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi_hi = {regroupV0_hi_12[1180], regroupV0_hi_12[1176]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi_4 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi_hi, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_8 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi_4, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo_lo = {regroupV0_hi_12[1188], regroupV0_hi_12[1184]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo_hi = {regroupV0_hi_12[1196], regroupV0_hi_12[1192]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo_4 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo_hi, regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi_lo = {regroupV0_hi_12[1204], regroupV0_hi_12[1200]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi_hi = {regroupV0_hi_12[1212], regroupV0_hi_12[1208]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi_4 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi_hi, regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_8 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi_4, regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_hi_lo_11 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_8, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_8};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo_lo = {regroupV0_hi_12[1220], regroupV0_hi_12[1216]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo_hi = {regroupV0_hi_12[1228], regroupV0_hi_12[1224]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo_4 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo_hi, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi_lo = {regroupV0_hi_12[1236], regroupV0_hi_12[1232]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi_hi = {regroupV0_hi_12[1244], regroupV0_hi_12[1240]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi_4 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi_hi, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_8 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi_4, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo_lo = {regroupV0_hi_12[1252], regroupV0_hi_12[1248]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo_hi = {regroupV0_hi_12[1260], regroupV0_hi_12[1256]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo_4 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo_hi, regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi_lo = {regroupV0_hi_12[1268], regroupV0_hi_12[1264]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi_hi = {regroupV0_hi_12[1276], regroupV0_hi_12[1272]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi_4 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi_hi, regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_8 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi_4, regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_hi_hi_11 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_8, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_8};
  wire [31:0]        regroupV0_hi_lo_hi_lo_lo_hi_11 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_11, regroupV0_hi_lo_hi_lo_lo_hi_lo_11};
  wire [63:0]        regroupV0_hi_lo_hi_lo_lo_11 = {regroupV0_hi_lo_hi_lo_lo_hi_11, regroupV0_hi_lo_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo_lo = {regroupV0_hi_12[1284], regroupV0_hi_12[1280]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo_hi = {regroupV0_hi_12[1292], regroupV0_hi_12[1288]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo_4 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo_hi, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi_lo = {regroupV0_hi_12[1300], regroupV0_hi_12[1296]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi_hi = {regroupV0_hi_12[1308], regroupV0_hi_12[1304]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi_4 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi_hi, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_8 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi_4, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo_lo = {regroupV0_hi_12[1316], regroupV0_hi_12[1312]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo_hi = {regroupV0_hi_12[1324], regroupV0_hi_12[1320]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo_4 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo_hi, regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi_lo = {regroupV0_hi_12[1332], regroupV0_hi_12[1328]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi_hi = {regroupV0_hi_12[1340], regroupV0_hi_12[1336]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi_4 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi_hi, regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_8 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi_4, regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_lo_lo_11 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_8, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_8};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo_lo = {regroupV0_hi_12[1348], regroupV0_hi_12[1344]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo_hi = {regroupV0_hi_12[1356], regroupV0_hi_12[1352]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo_4 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo_hi, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi_lo = {regroupV0_hi_12[1364], regroupV0_hi_12[1360]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi_hi = {regroupV0_hi_12[1372], regroupV0_hi_12[1368]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi_4 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi_hi, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_8 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi_4, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo_lo = {regroupV0_hi_12[1380], regroupV0_hi_12[1376]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo_hi = {regroupV0_hi_12[1388], regroupV0_hi_12[1384]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo_4 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo_hi, regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi_lo = {regroupV0_hi_12[1396], regroupV0_hi_12[1392]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi_hi = {regroupV0_hi_12[1404], regroupV0_hi_12[1400]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi_4 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi_hi, regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_8 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi_4, regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_lo_hi_11 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_8, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_8};
  wire [31:0]        regroupV0_hi_lo_hi_lo_hi_lo_11 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_11, regroupV0_hi_lo_hi_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo_lo = {regroupV0_hi_12[1412], regroupV0_hi_12[1408]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo_hi = {regroupV0_hi_12[1420], regroupV0_hi_12[1416]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo_4 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo_hi, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi_lo = {regroupV0_hi_12[1428], regroupV0_hi_12[1424]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi_hi = {regroupV0_hi_12[1436], regroupV0_hi_12[1432]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi_4 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi_hi, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_8 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi_4, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo_lo = {regroupV0_hi_12[1444], regroupV0_hi_12[1440]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo_hi = {regroupV0_hi_12[1452], regroupV0_hi_12[1448]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo_4 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo_hi, regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi_lo = {regroupV0_hi_12[1460], regroupV0_hi_12[1456]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi_hi = {regroupV0_hi_12[1468], regroupV0_hi_12[1464]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi_4 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi_hi, regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_8 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi_4, regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_hi_lo_11 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_8, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_8};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo_lo = {regroupV0_hi_12[1476], regroupV0_hi_12[1472]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo_hi = {regroupV0_hi_12[1484], regroupV0_hi_12[1480]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo_4 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo_hi, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi_lo = {regroupV0_hi_12[1492], regroupV0_hi_12[1488]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi_hi = {regroupV0_hi_12[1500], regroupV0_hi_12[1496]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi_4 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi_hi, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_8 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi_4, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo_lo = {regroupV0_hi_12[1508], regroupV0_hi_12[1504]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo_hi = {regroupV0_hi_12[1516], regroupV0_hi_12[1512]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo_4 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo_hi, regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi_lo = {regroupV0_hi_12[1524], regroupV0_hi_12[1520]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi_hi = {regroupV0_hi_12[1532], regroupV0_hi_12[1528]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi_4 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi_hi, regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_8 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi_4, regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_hi_hi_11 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_8, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_8};
  wire [31:0]        regroupV0_hi_lo_hi_lo_hi_hi_11 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_11, regroupV0_hi_lo_hi_lo_hi_hi_lo_11};
  wire [63:0]        regroupV0_hi_lo_hi_lo_hi_11 = {regroupV0_hi_lo_hi_lo_hi_hi_11, regroupV0_hi_lo_hi_lo_hi_lo_11};
  wire [127:0]       regroupV0_hi_lo_hi_lo_11 = {regroupV0_hi_lo_hi_lo_hi_11, regroupV0_hi_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo_lo = {regroupV0_hi_12[1540], regroupV0_hi_12[1536]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo_hi = {regroupV0_hi_12[1548], regroupV0_hi_12[1544]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo_4 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo_hi, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi_lo = {regroupV0_hi_12[1556], regroupV0_hi_12[1552]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi_hi = {regroupV0_hi_12[1564], regroupV0_hi_12[1560]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi_4 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi_hi, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_8 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi_4, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo_lo = {regroupV0_hi_12[1572], regroupV0_hi_12[1568]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo_hi = {regroupV0_hi_12[1580], regroupV0_hi_12[1576]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo_4 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo_hi, regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi_lo = {regroupV0_hi_12[1588], regroupV0_hi_12[1584]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi_hi = {regroupV0_hi_12[1596], regroupV0_hi_12[1592]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi_4 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi_hi, regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_8 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi_4, regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_lo_lo_11 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_8, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_8};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo_lo = {regroupV0_hi_12[1604], regroupV0_hi_12[1600]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo_hi = {regroupV0_hi_12[1612], regroupV0_hi_12[1608]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo_4 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo_hi, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi_lo = {regroupV0_hi_12[1620], regroupV0_hi_12[1616]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi_hi = {regroupV0_hi_12[1628], regroupV0_hi_12[1624]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi_4 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi_hi, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_8 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi_4, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo_lo = {regroupV0_hi_12[1636], regroupV0_hi_12[1632]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo_hi = {regroupV0_hi_12[1644], regroupV0_hi_12[1640]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo_4 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo_hi, regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi_lo = {regroupV0_hi_12[1652], regroupV0_hi_12[1648]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi_hi = {regroupV0_hi_12[1660], regroupV0_hi_12[1656]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi_4 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi_hi, regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_8 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi_4, regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_lo_hi_11 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_8, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_8};
  wire [31:0]        regroupV0_hi_lo_hi_hi_lo_lo_11 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_11, regroupV0_hi_lo_hi_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo_lo = {regroupV0_hi_12[1668], regroupV0_hi_12[1664]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo_hi = {regroupV0_hi_12[1676], regroupV0_hi_12[1672]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo_4 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo_hi, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi_lo = {regroupV0_hi_12[1684], regroupV0_hi_12[1680]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi_hi = {regroupV0_hi_12[1692], regroupV0_hi_12[1688]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi_4 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi_hi, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_8 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi_4, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo_lo = {regroupV0_hi_12[1700], regroupV0_hi_12[1696]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo_hi = {regroupV0_hi_12[1708], regroupV0_hi_12[1704]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo_4 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo_hi, regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi_lo = {regroupV0_hi_12[1716], regroupV0_hi_12[1712]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi_hi = {regroupV0_hi_12[1724], regroupV0_hi_12[1720]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi_4 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi_hi, regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_8 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi_4, regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_hi_lo_11 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_8, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_8};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo_lo = {regroupV0_hi_12[1732], regroupV0_hi_12[1728]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo_hi = {regroupV0_hi_12[1740], regroupV0_hi_12[1736]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo_4 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo_hi, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi_lo = {regroupV0_hi_12[1748], regroupV0_hi_12[1744]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi_hi = {regroupV0_hi_12[1756], regroupV0_hi_12[1752]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi_4 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi_hi, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_8 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi_4, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo_lo = {regroupV0_hi_12[1764], regroupV0_hi_12[1760]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo_hi = {regroupV0_hi_12[1772], regroupV0_hi_12[1768]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo_4 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo_hi, regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi_lo = {regroupV0_hi_12[1780], regroupV0_hi_12[1776]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi_hi = {regroupV0_hi_12[1788], regroupV0_hi_12[1784]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi_4 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi_hi, regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_8 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi_4, regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_hi_hi_11 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_8, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_8};
  wire [31:0]        regroupV0_hi_lo_hi_hi_lo_hi_11 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_11, regroupV0_hi_lo_hi_hi_lo_hi_lo_11};
  wire [63:0]        regroupV0_hi_lo_hi_hi_lo_11 = {regroupV0_hi_lo_hi_hi_lo_hi_11, regroupV0_hi_lo_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo_lo = {regroupV0_hi_12[1796], regroupV0_hi_12[1792]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo_hi = {regroupV0_hi_12[1804], regroupV0_hi_12[1800]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo_4 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo_hi, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi_lo = {regroupV0_hi_12[1812], regroupV0_hi_12[1808]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi_hi = {regroupV0_hi_12[1820], regroupV0_hi_12[1816]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi_4 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi_hi, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_8 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi_4, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo_lo = {regroupV0_hi_12[1828], regroupV0_hi_12[1824]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo_hi = {regroupV0_hi_12[1836], regroupV0_hi_12[1832]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo_4 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo_hi, regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi_lo = {regroupV0_hi_12[1844], regroupV0_hi_12[1840]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi_hi = {regroupV0_hi_12[1852], regroupV0_hi_12[1848]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi_4 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi_hi, regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_8 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi_4, regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_lo_lo_11 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_8, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_8};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo_lo = {regroupV0_hi_12[1860], regroupV0_hi_12[1856]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo_hi = {regroupV0_hi_12[1868], regroupV0_hi_12[1864]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo_4 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo_hi, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi_lo = {regroupV0_hi_12[1876], regroupV0_hi_12[1872]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi_hi = {regroupV0_hi_12[1884], regroupV0_hi_12[1880]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi_4 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi_hi, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_8 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi_4, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo_lo = {regroupV0_hi_12[1892], regroupV0_hi_12[1888]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo_hi = {regroupV0_hi_12[1900], regroupV0_hi_12[1896]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo_4 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo_hi, regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi_lo = {regroupV0_hi_12[1908], regroupV0_hi_12[1904]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi_hi = {regroupV0_hi_12[1916], regroupV0_hi_12[1912]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi_4 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi_hi, regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_8 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi_4, regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_lo_hi_11 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_8, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_8};
  wire [31:0]        regroupV0_hi_lo_hi_hi_hi_lo_11 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_11, regroupV0_hi_lo_hi_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo_lo = {regroupV0_hi_12[1924], regroupV0_hi_12[1920]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo_hi = {regroupV0_hi_12[1932], regroupV0_hi_12[1928]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo_4 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo_hi, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi_lo = {regroupV0_hi_12[1940], regroupV0_hi_12[1936]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi_hi = {regroupV0_hi_12[1948], regroupV0_hi_12[1944]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi_4 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi_hi, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_8 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi_4, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo_lo = {regroupV0_hi_12[1956], regroupV0_hi_12[1952]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo_hi = {regroupV0_hi_12[1964], regroupV0_hi_12[1960]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo_4 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo_hi, regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi_lo = {regroupV0_hi_12[1972], regroupV0_hi_12[1968]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi_hi = {regroupV0_hi_12[1980], regroupV0_hi_12[1976]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi_4 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi_hi, regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_8 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi_4, regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_hi_lo_11 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_8, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_8};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo_lo = {regroupV0_hi_12[1988], regroupV0_hi_12[1984]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo_hi = {regroupV0_hi_12[1996], regroupV0_hi_12[1992]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo_4 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo_hi, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi_lo = {regroupV0_hi_12[2004], regroupV0_hi_12[2000]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi_hi = {regroupV0_hi_12[2012], regroupV0_hi_12[2008]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi_4 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi_hi, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_8 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi_4, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo_lo = {regroupV0_hi_12[2020], regroupV0_hi_12[2016]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo_hi = {regroupV0_hi_12[2028], regroupV0_hi_12[2024]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo_4 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo_hi, regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi_lo = {regroupV0_hi_12[2036], regroupV0_hi_12[2032]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi_hi = {regroupV0_hi_12[2044], regroupV0_hi_12[2040]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi_4 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi_hi, regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_8 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi_4, regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_hi_hi_11 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_8, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_8};
  wire [31:0]        regroupV0_hi_lo_hi_hi_hi_hi_11 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_11, regroupV0_hi_lo_hi_hi_hi_hi_lo_11};
  wire [63:0]        regroupV0_hi_lo_hi_hi_hi_11 = {regroupV0_hi_lo_hi_hi_hi_hi_11, regroupV0_hi_lo_hi_hi_hi_lo_11};
  wire [127:0]       regroupV0_hi_lo_hi_hi_11 = {regroupV0_hi_lo_hi_hi_hi_11, regroupV0_hi_lo_hi_hi_lo_11};
  wire [255:0]       regroupV0_hi_lo_hi_11 = {regroupV0_hi_lo_hi_hi_11, regroupV0_hi_lo_hi_lo_11};
  wire [511:0]       regroupV0_hi_lo_11 = {regroupV0_hi_lo_hi_11, regroupV0_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo_lo = {regroupV0_hi_12[2052], regroupV0_hi_12[2048]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo_hi = {regroupV0_hi_12[2060], regroupV0_hi_12[2056]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo_4 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo_hi, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi_lo = {regroupV0_hi_12[2068], regroupV0_hi_12[2064]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi_hi = {regroupV0_hi_12[2076], regroupV0_hi_12[2072]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi_4 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi_hi, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_8 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi_4, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo_lo = {regroupV0_hi_12[2084], regroupV0_hi_12[2080]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo_hi = {regroupV0_hi_12[2092], regroupV0_hi_12[2088]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo_4 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo_hi, regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi_lo = {regroupV0_hi_12[2100], regroupV0_hi_12[2096]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi_hi = {regroupV0_hi_12[2108], regroupV0_hi_12[2104]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi_4 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi_hi, regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_8 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi_4, regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_lo_lo_11 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_8, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_8};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo_lo = {regroupV0_hi_12[2116], regroupV0_hi_12[2112]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo_hi = {regroupV0_hi_12[2124], regroupV0_hi_12[2120]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo_4 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo_hi, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi_lo = {regroupV0_hi_12[2132], regroupV0_hi_12[2128]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi_hi = {regroupV0_hi_12[2140], regroupV0_hi_12[2136]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi_4 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi_hi, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_8 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi_4, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo_lo = {regroupV0_hi_12[2148], regroupV0_hi_12[2144]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo_hi = {regroupV0_hi_12[2156], regroupV0_hi_12[2152]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo_4 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo_hi, regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi_lo = {regroupV0_hi_12[2164], regroupV0_hi_12[2160]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi_hi = {regroupV0_hi_12[2172], regroupV0_hi_12[2168]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi_4 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi_hi, regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_8 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi_4, regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_lo_hi_11 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_8, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_8};
  wire [31:0]        regroupV0_hi_hi_lo_lo_lo_lo_11 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_11, regroupV0_hi_hi_lo_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo_lo = {regroupV0_hi_12[2180], regroupV0_hi_12[2176]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo_hi = {regroupV0_hi_12[2188], regroupV0_hi_12[2184]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo_4 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo_hi, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi_lo = {regroupV0_hi_12[2196], regroupV0_hi_12[2192]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi_hi = {regroupV0_hi_12[2204], regroupV0_hi_12[2200]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi_4 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi_hi, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_8 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi_4, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo_lo = {regroupV0_hi_12[2212], regroupV0_hi_12[2208]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo_hi = {regroupV0_hi_12[2220], regroupV0_hi_12[2216]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo_4 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo_hi, regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi_lo = {regroupV0_hi_12[2228], regroupV0_hi_12[2224]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi_hi = {regroupV0_hi_12[2236], regroupV0_hi_12[2232]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi_4 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi_hi, regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_8 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi_4, regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_hi_lo_11 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_8, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_8};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo_lo = {regroupV0_hi_12[2244], regroupV0_hi_12[2240]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo_hi = {regroupV0_hi_12[2252], regroupV0_hi_12[2248]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo_4 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo_hi, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi_lo = {regroupV0_hi_12[2260], regroupV0_hi_12[2256]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi_hi = {regroupV0_hi_12[2268], regroupV0_hi_12[2264]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi_4 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi_hi, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_8 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi_4, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo_lo = {regroupV0_hi_12[2276], regroupV0_hi_12[2272]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo_hi = {regroupV0_hi_12[2284], regroupV0_hi_12[2280]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo_4 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo_hi, regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi_lo = {regroupV0_hi_12[2292], regroupV0_hi_12[2288]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi_hi = {regroupV0_hi_12[2300], regroupV0_hi_12[2296]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi_4 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi_hi, regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_8 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi_4, regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_hi_hi_11 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_8, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_8};
  wire [31:0]        regroupV0_hi_hi_lo_lo_lo_hi_11 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_11, regroupV0_hi_hi_lo_lo_lo_hi_lo_11};
  wire [63:0]        regroupV0_hi_hi_lo_lo_lo_11 = {regroupV0_hi_hi_lo_lo_lo_hi_11, regroupV0_hi_hi_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo_lo = {regroupV0_hi_12[2308], regroupV0_hi_12[2304]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo_hi = {regroupV0_hi_12[2316], regroupV0_hi_12[2312]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo_4 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo_hi, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi_lo = {regroupV0_hi_12[2324], regroupV0_hi_12[2320]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi_hi = {regroupV0_hi_12[2332], regroupV0_hi_12[2328]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi_4 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi_hi, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_8 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi_4, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo_lo = {regroupV0_hi_12[2340], regroupV0_hi_12[2336]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo_hi = {regroupV0_hi_12[2348], regroupV0_hi_12[2344]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo_4 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo_hi, regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi_lo = {regroupV0_hi_12[2356], regroupV0_hi_12[2352]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi_hi = {regroupV0_hi_12[2364], regroupV0_hi_12[2360]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi_4 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi_hi, regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_8 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi_4, regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_lo_lo_11 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_8, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_8};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo_lo = {regroupV0_hi_12[2372], regroupV0_hi_12[2368]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo_hi = {regroupV0_hi_12[2380], regroupV0_hi_12[2376]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo_4 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo_hi, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi_lo = {regroupV0_hi_12[2388], regroupV0_hi_12[2384]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi_hi = {regroupV0_hi_12[2396], regroupV0_hi_12[2392]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi_4 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi_hi, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_8 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi_4, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo_lo = {regroupV0_hi_12[2404], regroupV0_hi_12[2400]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo_hi = {regroupV0_hi_12[2412], regroupV0_hi_12[2408]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo_4 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo_hi, regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi_lo = {regroupV0_hi_12[2420], regroupV0_hi_12[2416]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi_hi = {regroupV0_hi_12[2428], regroupV0_hi_12[2424]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi_4 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi_hi, regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_8 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi_4, regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_lo_hi_11 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_8, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_8};
  wire [31:0]        regroupV0_hi_hi_lo_lo_hi_lo_11 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_11, regroupV0_hi_hi_lo_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo_lo = {regroupV0_hi_12[2436], regroupV0_hi_12[2432]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo_hi = {regroupV0_hi_12[2444], regroupV0_hi_12[2440]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo_4 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo_hi, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi_lo = {regroupV0_hi_12[2452], regroupV0_hi_12[2448]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi_hi = {regroupV0_hi_12[2460], regroupV0_hi_12[2456]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi_4 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi_hi, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_8 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi_4, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo_lo = {regroupV0_hi_12[2468], regroupV0_hi_12[2464]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo_hi = {regroupV0_hi_12[2476], regroupV0_hi_12[2472]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo_4 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo_hi, regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi_lo = {regroupV0_hi_12[2484], regroupV0_hi_12[2480]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi_hi = {regroupV0_hi_12[2492], regroupV0_hi_12[2488]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi_4 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi_hi, regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_8 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi_4, regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_hi_lo_11 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_8, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_8};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo_lo = {regroupV0_hi_12[2500], regroupV0_hi_12[2496]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo_hi = {regroupV0_hi_12[2508], regroupV0_hi_12[2504]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo_4 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo_hi, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi_lo = {regroupV0_hi_12[2516], regroupV0_hi_12[2512]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi_hi = {regroupV0_hi_12[2524], regroupV0_hi_12[2520]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi_4 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi_hi, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_8 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi_4, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo_lo = {regroupV0_hi_12[2532], regroupV0_hi_12[2528]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo_hi = {regroupV0_hi_12[2540], regroupV0_hi_12[2536]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo_4 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo_hi, regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi_lo = {regroupV0_hi_12[2548], regroupV0_hi_12[2544]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi_hi = {regroupV0_hi_12[2556], regroupV0_hi_12[2552]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi_4 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi_hi, regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_8 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi_4, regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_hi_hi_11 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_8, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_8};
  wire [31:0]        regroupV0_hi_hi_lo_lo_hi_hi_11 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_11, regroupV0_hi_hi_lo_lo_hi_hi_lo_11};
  wire [63:0]        regroupV0_hi_hi_lo_lo_hi_11 = {regroupV0_hi_hi_lo_lo_hi_hi_11, regroupV0_hi_hi_lo_lo_hi_lo_11};
  wire [127:0]       regroupV0_hi_hi_lo_lo_11 = {regroupV0_hi_hi_lo_lo_hi_11, regroupV0_hi_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo_lo = {regroupV0_hi_12[2564], regroupV0_hi_12[2560]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo_hi = {regroupV0_hi_12[2572], regroupV0_hi_12[2568]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo_4 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo_hi, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi_lo = {regroupV0_hi_12[2580], regroupV0_hi_12[2576]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi_hi = {regroupV0_hi_12[2588], regroupV0_hi_12[2584]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi_4 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi_hi, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_8 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi_4, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo_lo = {regroupV0_hi_12[2596], regroupV0_hi_12[2592]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo_hi = {regroupV0_hi_12[2604], regroupV0_hi_12[2600]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo_4 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo_hi, regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi_lo = {regroupV0_hi_12[2612], regroupV0_hi_12[2608]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi_hi = {regroupV0_hi_12[2620], regroupV0_hi_12[2616]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi_4 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi_hi, regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_8 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi_4, regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_lo_lo_11 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_8, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_8};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo_lo = {regroupV0_hi_12[2628], regroupV0_hi_12[2624]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo_hi = {regroupV0_hi_12[2636], regroupV0_hi_12[2632]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo_4 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo_hi, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi_lo = {regroupV0_hi_12[2644], regroupV0_hi_12[2640]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi_hi = {regroupV0_hi_12[2652], regroupV0_hi_12[2648]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi_4 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi_hi, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_8 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi_4, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo_lo = {regroupV0_hi_12[2660], regroupV0_hi_12[2656]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo_hi = {regroupV0_hi_12[2668], regroupV0_hi_12[2664]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo_4 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo_hi, regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi_lo = {regroupV0_hi_12[2676], regroupV0_hi_12[2672]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi_hi = {regroupV0_hi_12[2684], regroupV0_hi_12[2680]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi_4 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi_hi, regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_8 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi_4, regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_lo_hi_11 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_8, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_8};
  wire [31:0]        regroupV0_hi_hi_lo_hi_lo_lo_11 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_11, regroupV0_hi_hi_lo_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo_lo = {regroupV0_hi_12[2692], regroupV0_hi_12[2688]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo_hi = {regroupV0_hi_12[2700], regroupV0_hi_12[2696]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo_4 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo_hi, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi_lo = {regroupV0_hi_12[2708], regroupV0_hi_12[2704]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi_hi = {regroupV0_hi_12[2716], regroupV0_hi_12[2712]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi_4 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi_hi, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_8 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi_4, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo_lo = {regroupV0_hi_12[2724], regroupV0_hi_12[2720]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo_hi = {regroupV0_hi_12[2732], regroupV0_hi_12[2728]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo_4 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo_hi, regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi_lo = {regroupV0_hi_12[2740], regroupV0_hi_12[2736]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi_hi = {regroupV0_hi_12[2748], regroupV0_hi_12[2744]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi_4 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi_hi, regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_8 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi_4, regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_hi_lo_11 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_8, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_8};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo_lo = {regroupV0_hi_12[2756], regroupV0_hi_12[2752]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo_hi = {regroupV0_hi_12[2764], regroupV0_hi_12[2760]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo_4 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo_hi, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi_lo = {regroupV0_hi_12[2772], regroupV0_hi_12[2768]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi_hi = {regroupV0_hi_12[2780], regroupV0_hi_12[2776]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi_4 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi_hi, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_8 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi_4, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo_lo = {regroupV0_hi_12[2788], regroupV0_hi_12[2784]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo_hi = {regroupV0_hi_12[2796], regroupV0_hi_12[2792]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo_4 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo_hi, regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi_lo = {regroupV0_hi_12[2804], regroupV0_hi_12[2800]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi_hi = {regroupV0_hi_12[2812], regroupV0_hi_12[2808]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi_4 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi_hi, regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_8 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi_4, regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_hi_hi_11 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_8, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_8};
  wire [31:0]        regroupV0_hi_hi_lo_hi_lo_hi_11 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_11, regroupV0_hi_hi_lo_hi_lo_hi_lo_11};
  wire [63:0]        regroupV0_hi_hi_lo_hi_lo_11 = {regroupV0_hi_hi_lo_hi_lo_hi_11, regroupV0_hi_hi_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo_lo = {regroupV0_hi_12[2820], regroupV0_hi_12[2816]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo_hi = {regroupV0_hi_12[2828], regroupV0_hi_12[2824]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo_4 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo_hi, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi_lo = {regroupV0_hi_12[2836], regroupV0_hi_12[2832]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi_hi = {regroupV0_hi_12[2844], regroupV0_hi_12[2840]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi_4 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi_hi, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_8 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi_4, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo_lo = {regroupV0_hi_12[2852], regroupV0_hi_12[2848]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo_hi = {regroupV0_hi_12[2860], regroupV0_hi_12[2856]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo_4 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo_hi, regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi_lo = {regroupV0_hi_12[2868], regroupV0_hi_12[2864]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi_hi = {regroupV0_hi_12[2876], regroupV0_hi_12[2872]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi_4 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi_hi, regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_8 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi_4, regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_lo_lo_11 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_8, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_8};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo_lo = {regroupV0_hi_12[2884], regroupV0_hi_12[2880]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo_hi = {regroupV0_hi_12[2892], regroupV0_hi_12[2888]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo_4 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo_hi, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi_lo = {regroupV0_hi_12[2900], regroupV0_hi_12[2896]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi_hi = {regroupV0_hi_12[2908], regroupV0_hi_12[2904]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi_4 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi_hi, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_8 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi_4, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo_lo = {regroupV0_hi_12[2916], regroupV0_hi_12[2912]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo_hi = {regroupV0_hi_12[2924], regroupV0_hi_12[2920]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo_4 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo_hi, regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi_lo = {regroupV0_hi_12[2932], regroupV0_hi_12[2928]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi_hi = {regroupV0_hi_12[2940], regroupV0_hi_12[2936]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi_4 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi_hi, regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_8 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi_4, regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_lo_hi_11 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_8, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_8};
  wire [31:0]        regroupV0_hi_hi_lo_hi_hi_lo_11 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_11, regroupV0_hi_hi_lo_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo_lo = {regroupV0_hi_12[2948], regroupV0_hi_12[2944]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo_hi = {regroupV0_hi_12[2956], regroupV0_hi_12[2952]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo_4 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo_hi, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi_lo = {regroupV0_hi_12[2964], regroupV0_hi_12[2960]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi_hi = {regroupV0_hi_12[2972], regroupV0_hi_12[2968]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi_4 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi_hi, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_8 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi_4, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo_lo = {regroupV0_hi_12[2980], regroupV0_hi_12[2976]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo_hi = {regroupV0_hi_12[2988], regroupV0_hi_12[2984]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo_4 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo_hi, regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi_lo = {regroupV0_hi_12[2996], regroupV0_hi_12[2992]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi_hi = {regroupV0_hi_12[3004], regroupV0_hi_12[3000]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi_4 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi_hi, regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_8 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi_4, regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_hi_lo_11 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_8, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_8};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo_lo = {regroupV0_hi_12[3012], regroupV0_hi_12[3008]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo_hi = {regroupV0_hi_12[3020], regroupV0_hi_12[3016]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo_4 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo_hi, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi_lo = {regroupV0_hi_12[3028], regroupV0_hi_12[3024]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi_hi = {regroupV0_hi_12[3036], regroupV0_hi_12[3032]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi_4 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi_hi, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_8 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi_4, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo_lo = {regroupV0_hi_12[3044], regroupV0_hi_12[3040]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo_hi = {regroupV0_hi_12[3052], regroupV0_hi_12[3048]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo_4 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo_hi, regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi_lo = {regroupV0_hi_12[3060], regroupV0_hi_12[3056]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi_hi = {regroupV0_hi_12[3068], regroupV0_hi_12[3064]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi_4 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi_hi, regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_8 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi_4, regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_hi_hi_11 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_8, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_8};
  wire [31:0]        regroupV0_hi_hi_lo_hi_hi_hi_11 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_11, regroupV0_hi_hi_lo_hi_hi_hi_lo_11};
  wire [63:0]        regroupV0_hi_hi_lo_hi_hi_11 = {regroupV0_hi_hi_lo_hi_hi_hi_11, regroupV0_hi_hi_lo_hi_hi_lo_11};
  wire [127:0]       regroupV0_hi_hi_lo_hi_11 = {regroupV0_hi_hi_lo_hi_hi_11, regroupV0_hi_hi_lo_hi_lo_11};
  wire [255:0]       regroupV0_hi_hi_lo_11 = {regroupV0_hi_hi_lo_hi_11, regroupV0_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo_lo = {regroupV0_hi_12[3076], regroupV0_hi_12[3072]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo_hi = {regroupV0_hi_12[3084], regroupV0_hi_12[3080]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo_4 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo_hi, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi_lo = {regroupV0_hi_12[3092], regroupV0_hi_12[3088]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi_hi = {regroupV0_hi_12[3100], regroupV0_hi_12[3096]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi_4 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi_hi, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_8 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi_4, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo_lo = {regroupV0_hi_12[3108], regroupV0_hi_12[3104]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo_hi = {regroupV0_hi_12[3116], regroupV0_hi_12[3112]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo_4 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo_hi, regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi_lo = {regroupV0_hi_12[3124], regroupV0_hi_12[3120]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi_hi = {regroupV0_hi_12[3132], regroupV0_hi_12[3128]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi_4 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi_hi, regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_8 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi_4, regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_lo_lo_11 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_8, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_8};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo_lo = {regroupV0_hi_12[3140], regroupV0_hi_12[3136]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo_hi = {regroupV0_hi_12[3148], regroupV0_hi_12[3144]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo_4 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo_hi, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi_lo = {regroupV0_hi_12[3156], regroupV0_hi_12[3152]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi_hi = {regroupV0_hi_12[3164], regroupV0_hi_12[3160]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi_4 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi_hi, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_8 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi_4, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo_lo = {regroupV0_hi_12[3172], regroupV0_hi_12[3168]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo_hi = {regroupV0_hi_12[3180], regroupV0_hi_12[3176]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo_4 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo_hi, regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi_lo = {regroupV0_hi_12[3188], regroupV0_hi_12[3184]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi_hi = {regroupV0_hi_12[3196], regroupV0_hi_12[3192]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi_4 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi_hi, regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_8 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi_4, regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_lo_hi_11 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_8, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_8};
  wire [31:0]        regroupV0_hi_hi_hi_lo_lo_lo_11 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_11, regroupV0_hi_hi_hi_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo_lo = {regroupV0_hi_12[3204], regroupV0_hi_12[3200]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo_hi = {regroupV0_hi_12[3212], regroupV0_hi_12[3208]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo_4 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo_hi, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi_lo = {regroupV0_hi_12[3220], regroupV0_hi_12[3216]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi_hi = {regroupV0_hi_12[3228], regroupV0_hi_12[3224]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi_4 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi_hi, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_8 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi_4, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo_lo = {regroupV0_hi_12[3236], regroupV0_hi_12[3232]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo_hi = {regroupV0_hi_12[3244], regroupV0_hi_12[3240]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo_4 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo_hi, regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi_lo = {regroupV0_hi_12[3252], regroupV0_hi_12[3248]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi_hi = {regroupV0_hi_12[3260], regroupV0_hi_12[3256]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi_4 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi_hi, regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_8 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi_4, regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_hi_lo_11 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_8, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_8};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo_lo = {regroupV0_hi_12[3268], regroupV0_hi_12[3264]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo_hi = {regroupV0_hi_12[3276], regroupV0_hi_12[3272]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo_4 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo_hi, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi_lo = {regroupV0_hi_12[3284], regroupV0_hi_12[3280]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi_hi = {regroupV0_hi_12[3292], regroupV0_hi_12[3288]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi_4 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi_hi, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_8 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi_4, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo_lo = {regroupV0_hi_12[3300], regroupV0_hi_12[3296]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo_hi = {regroupV0_hi_12[3308], regroupV0_hi_12[3304]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo_4 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo_hi, regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi_lo = {regroupV0_hi_12[3316], regroupV0_hi_12[3312]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi_hi = {regroupV0_hi_12[3324], regroupV0_hi_12[3320]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi_4 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi_hi, regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_8 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi_4, regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_hi_hi_11 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_8, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_8};
  wire [31:0]        regroupV0_hi_hi_hi_lo_lo_hi_11 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_11, regroupV0_hi_hi_hi_lo_lo_hi_lo_11};
  wire [63:0]        regroupV0_hi_hi_hi_lo_lo_11 = {regroupV0_hi_hi_hi_lo_lo_hi_11, regroupV0_hi_hi_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo_lo = {regroupV0_hi_12[3332], regroupV0_hi_12[3328]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo_hi = {regroupV0_hi_12[3340], regroupV0_hi_12[3336]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo_4 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo_hi, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi_lo = {regroupV0_hi_12[3348], regroupV0_hi_12[3344]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi_hi = {regroupV0_hi_12[3356], regroupV0_hi_12[3352]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi_4 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi_hi, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_8 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi_4, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo_lo = {regroupV0_hi_12[3364], regroupV0_hi_12[3360]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo_hi = {regroupV0_hi_12[3372], regroupV0_hi_12[3368]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo_4 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo_hi, regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi_lo = {regroupV0_hi_12[3380], regroupV0_hi_12[3376]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi_hi = {regroupV0_hi_12[3388], regroupV0_hi_12[3384]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi_4 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi_hi, regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_8 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi_4, regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_lo_lo_11 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_8, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_8};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo_lo = {regroupV0_hi_12[3396], regroupV0_hi_12[3392]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo_hi = {regroupV0_hi_12[3404], regroupV0_hi_12[3400]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo_4 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo_hi, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi_lo = {regroupV0_hi_12[3412], regroupV0_hi_12[3408]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi_hi = {regroupV0_hi_12[3420], regroupV0_hi_12[3416]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi_4 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi_hi, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_8 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi_4, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo_lo = {regroupV0_hi_12[3428], regroupV0_hi_12[3424]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo_hi = {regroupV0_hi_12[3436], regroupV0_hi_12[3432]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo_4 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo_hi, regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi_lo = {regroupV0_hi_12[3444], regroupV0_hi_12[3440]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi_hi = {regroupV0_hi_12[3452], regroupV0_hi_12[3448]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi_4 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi_hi, regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_8 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi_4, regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_lo_hi_11 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_8, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_8};
  wire [31:0]        regroupV0_hi_hi_hi_lo_hi_lo_11 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_11, regroupV0_hi_hi_hi_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo_lo = {regroupV0_hi_12[3460], regroupV0_hi_12[3456]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo_hi = {regroupV0_hi_12[3468], regroupV0_hi_12[3464]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo_4 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo_hi, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi_lo = {regroupV0_hi_12[3476], regroupV0_hi_12[3472]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi_hi = {regroupV0_hi_12[3484], regroupV0_hi_12[3480]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi_4 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi_hi, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_8 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi_4, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo_lo = {regroupV0_hi_12[3492], regroupV0_hi_12[3488]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo_hi = {regroupV0_hi_12[3500], regroupV0_hi_12[3496]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo_4 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo_hi, regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi_lo = {regroupV0_hi_12[3508], regroupV0_hi_12[3504]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi_hi = {regroupV0_hi_12[3516], regroupV0_hi_12[3512]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi_4 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi_hi, regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_8 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi_4, regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_hi_lo_11 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_8, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_8};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo_lo = {regroupV0_hi_12[3524], regroupV0_hi_12[3520]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo_hi = {regroupV0_hi_12[3532], regroupV0_hi_12[3528]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo_4 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo_hi, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi_lo = {regroupV0_hi_12[3540], regroupV0_hi_12[3536]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi_hi = {regroupV0_hi_12[3548], regroupV0_hi_12[3544]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi_4 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi_hi, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_8 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi_4, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo_lo = {regroupV0_hi_12[3556], regroupV0_hi_12[3552]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo_hi = {regroupV0_hi_12[3564], regroupV0_hi_12[3560]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo_4 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo_hi, regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi_lo = {regroupV0_hi_12[3572], regroupV0_hi_12[3568]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi_hi = {regroupV0_hi_12[3580], regroupV0_hi_12[3576]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi_4 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi_hi, regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_8 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi_4, regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_hi_hi_11 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_8, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_8};
  wire [31:0]        regroupV0_hi_hi_hi_lo_hi_hi_11 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_11, regroupV0_hi_hi_hi_lo_hi_hi_lo_11};
  wire [63:0]        regroupV0_hi_hi_hi_lo_hi_11 = {regroupV0_hi_hi_hi_lo_hi_hi_11, regroupV0_hi_hi_hi_lo_hi_lo_11};
  wire [127:0]       regroupV0_hi_hi_hi_lo_11 = {regroupV0_hi_hi_hi_lo_hi_11, regroupV0_hi_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo_lo = {regroupV0_hi_12[3588], regroupV0_hi_12[3584]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo_hi = {regroupV0_hi_12[3596], regroupV0_hi_12[3592]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo_4 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo_hi, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi_lo = {regroupV0_hi_12[3604], regroupV0_hi_12[3600]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi_hi = {regroupV0_hi_12[3612], regroupV0_hi_12[3608]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi_4 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi_hi, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_8 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi_4, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo_lo = {regroupV0_hi_12[3620], regroupV0_hi_12[3616]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo_hi = {regroupV0_hi_12[3628], regroupV0_hi_12[3624]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo_4 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo_hi, regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi_lo = {regroupV0_hi_12[3636], regroupV0_hi_12[3632]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi_hi = {regroupV0_hi_12[3644], regroupV0_hi_12[3640]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi_4 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi_hi, regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_8 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi_4, regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_lo_lo_11 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_8, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_8};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo_lo = {regroupV0_hi_12[3652], regroupV0_hi_12[3648]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo_hi = {regroupV0_hi_12[3660], regroupV0_hi_12[3656]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo_4 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo_hi, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi_lo = {regroupV0_hi_12[3668], regroupV0_hi_12[3664]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi_hi = {regroupV0_hi_12[3676], regroupV0_hi_12[3672]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi_4 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi_hi, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_8 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi_4, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo_lo = {regroupV0_hi_12[3684], regroupV0_hi_12[3680]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo_hi = {regroupV0_hi_12[3692], regroupV0_hi_12[3688]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo_4 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo_hi, regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi_lo = {regroupV0_hi_12[3700], regroupV0_hi_12[3696]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi_hi = {regroupV0_hi_12[3708], regroupV0_hi_12[3704]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi_4 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi_hi, regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_8 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi_4, regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_lo_hi_11 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_8, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_8};
  wire [31:0]        regroupV0_hi_hi_hi_hi_lo_lo_11 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_11, regroupV0_hi_hi_hi_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo_lo = {regroupV0_hi_12[3716], regroupV0_hi_12[3712]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo_hi = {regroupV0_hi_12[3724], regroupV0_hi_12[3720]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo_4 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo_hi, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi_lo = {regroupV0_hi_12[3732], regroupV0_hi_12[3728]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi_hi = {regroupV0_hi_12[3740], regroupV0_hi_12[3736]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi_4 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi_hi, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_8 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi_4, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo_lo = {regroupV0_hi_12[3748], regroupV0_hi_12[3744]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo_hi = {regroupV0_hi_12[3756], regroupV0_hi_12[3752]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo_4 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo_hi, regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi_lo = {regroupV0_hi_12[3764], regroupV0_hi_12[3760]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi_hi = {regroupV0_hi_12[3772], regroupV0_hi_12[3768]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi_4 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi_hi, regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_8 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi_4, regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_hi_lo_11 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_8, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_8};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo_lo = {regroupV0_hi_12[3780], regroupV0_hi_12[3776]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo_hi = {regroupV0_hi_12[3788], regroupV0_hi_12[3784]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo_4 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo_hi, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi_lo = {regroupV0_hi_12[3796], regroupV0_hi_12[3792]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi_hi = {regroupV0_hi_12[3804], regroupV0_hi_12[3800]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi_4 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi_hi, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_8 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi_4, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo_lo = {regroupV0_hi_12[3812], regroupV0_hi_12[3808]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo_hi = {regroupV0_hi_12[3820], regroupV0_hi_12[3816]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo_4 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo_hi, regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi_lo = {regroupV0_hi_12[3828], regroupV0_hi_12[3824]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi_hi = {regroupV0_hi_12[3836], regroupV0_hi_12[3832]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi_4 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi_hi, regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_8 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi_4, regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_hi_hi_11 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_8, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_8};
  wire [31:0]        regroupV0_hi_hi_hi_hi_lo_hi_11 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_11, regroupV0_hi_hi_hi_hi_lo_hi_lo_11};
  wire [63:0]        regroupV0_hi_hi_hi_hi_lo_11 = {regroupV0_hi_hi_hi_hi_lo_hi_11, regroupV0_hi_hi_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo_lo = {regroupV0_hi_12[3844], regroupV0_hi_12[3840]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo_hi = {regroupV0_hi_12[3852], regroupV0_hi_12[3848]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo_4 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo_hi, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi_lo = {regroupV0_hi_12[3860], regroupV0_hi_12[3856]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi_hi = {regroupV0_hi_12[3868], regroupV0_hi_12[3864]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi_4 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi_hi, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_8 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi_4, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo_lo = {regroupV0_hi_12[3876], regroupV0_hi_12[3872]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo_hi = {regroupV0_hi_12[3884], regroupV0_hi_12[3880]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo_4 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo_hi, regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi_lo = {regroupV0_hi_12[3892], regroupV0_hi_12[3888]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi_hi = {regroupV0_hi_12[3900], regroupV0_hi_12[3896]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi_4 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi_hi, regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_8 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi_4, regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_lo_lo_11 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_8, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_8};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo_lo = {regroupV0_hi_12[3908], regroupV0_hi_12[3904]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo_hi = {regroupV0_hi_12[3916], regroupV0_hi_12[3912]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo_4 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo_hi, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi_lo = {regroupV0_hi_12[3924], regroupV0_hi_12[3920]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi_hi = {regroupV0_hi_12[3932], regroupV0_hi_12[3928]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi_4 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi_hi, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_8 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi_4, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo_lo = {regroupV0_hi_12[3940], regroupV0_hi_12[3936]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo_hi = {regroupV0_hi_12[3948], regroupV0_hi_12[3944]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo_4 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo_hi, regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi_lo = {regroupV0_hi_12[3956], regroupV0_hi_12[3952]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi_hi = {regroupV0_hi_12[3964], regroupV0_hi_12[3960]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi_4 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi_hi, regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_8 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi_4, regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_lo_hi_11 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_8, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_8};
  wire [31:0]        regroupV0_hi_hi_hi_hi_hi_lo_11 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_11, regroupV0_hi_hi_hi_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo_lo = {regroupV0_hi_12[3972], regroupV0_hi_12[3968]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo_hi = {regroupV0_hi_12[3980], regroupV0_hi_12[3976]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo_4 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo_hi, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi_lo = {regroupV0_hi_12[3988], regroupV0_hi_12[3984]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi_hi = {regroupV0_hi_12[3996], regroupV0_hi_12[3992]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi_4 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi_hi, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_8 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi_4, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo_lo = {regroupV0_hi_12[4004], regroupV0_hi_12[4000]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo_hi = {regroupV0_hi_12[4012], regroupV0_hi_12[4008]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo_4 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo_hi, regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi_lo = {regroupV0_hi_12[4020], regroupV0_hi_12[4016]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi_hi = {regroupV0_hi_12[4028], regroupV0_hi_12[4024]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi_4 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi_hi, regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_8 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi_4, regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_hi_lo_11 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_8, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_8};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo_lo = {regroupV0_hi_12[4036], regroupV0_hi_12[4032]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo_hi = {regroupV0_hi_12[4044], regroupV0_hi_12[4040]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo_4 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo_hi, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi_lo = {regroupV0_hi_12[4052], regroupV0_hi_12[4048]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi_hi = {regroupV0_hi_12[4060], regroupV0_hi_12[4056]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi_4 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi_hi, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_8 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi_4, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo_lo = {regroupV0_hi_12[4068], regroupV0_hi_12[4064]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo_hi = {regroupV0_hi_12[4076], regroupV0_hi_12[4072]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo_4 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo_hi, regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi_lo = {regroupV0_hi_12[4084], regroupV0_hi_12[4080]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi_hi = {regroupV0_hi_12[4092], regroupV0_hi_12[4088]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi_4 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi_hi, regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_8 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi_4, regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_hi_hi_11 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_8, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_8};
  wire [31:0]        regroupV0_hi_hi_hi_hi_hi_hi_11 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_11, regroupV0_hi_hi_hi_hi_hi_hi_lo_11};
  wire [63:0]        regroupV0_hi_hi_hi_hi_hi_11 = {regroupV0_hi_hi_hi_hi_hi_hi_11, regroupV0_hi_hi_hi_hi_hi_lo_11};
  wire [127:0]       regroupV0_hi_hi_hi_hi_11 = {regroupV0_hi_hi_hi_hi_hi_11, regroupV0_hi_hi_hi_hi_lo_11};
  wire [255:0]       regroupV0_hi_hi_hi_11 = {regroupV0_hi_hi_hi_hi_11, regroupV0_hi_hi_hi_lo_11};
  wire [511:0]       regroupV0_hi_hi_11 = {regroupV0_hi_hi_hi_11, regroupV0_hi_hi_lo_11};
  wire [1023:0]      regroupV0_hi_13 = {regroupV0_hi_hi_11, regroupV0_hi_lo_11};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo_lo_1 = {regroupV0_lo_12[5], regroupV0_lo_12[1]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo_hi_1 = {regroupV0_lo_12[13], regroupV0_lo_12[9]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo_5 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi_lo_1 = {regroupV0_lo_12[21], regroupV0_lo_12[17]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi_hi_1 = {regroupV0_lo_12[29], regroupV0_lo_12[25]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi_5 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi_hi_1, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_9 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi_5, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo_lo_1 = {regroupV0_lo_12[37], regroupV0_lo_12[33]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo_hi_1 = {regroupV0_lo_12[45], regroupV0_lo_12[41]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo_5 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo_hi_1, regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi_lo_1 = {regroupV0_lo_12[53], regroupV0_lo_12[49]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi_hi_1 = {regroupV0_lo_12[61], regroupV0_lo_12[57]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi_5 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi_hi_1, regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_9 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi_5, regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_lo_lo_12 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_9, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_9};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo_lo_1 = {regroupV0_lo_12[69], regroupV0_lo_12[65]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo_hi_1 = {regroupV0_lo_12[77], regroupV0_lo_12[73]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo_5 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi_lo_1 = {regroupV0_lo_12[85], regroupV0_lo_12[81]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi_hi_1 = {regroupV0_lo_12[93], regroupV0_lo_12[89]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi_5 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi_hi_1, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_9 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi_5, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo_lo_1 = {regroupV0_lo_12[101], regroupV0_lo_12[97]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo_hi_1 = {regroupV0_lo_12[109], regroupV0_lo_12[105]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo_5 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo_hi_1, regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi_lo_1 = {regroupV0_lo_12[117], regroupV0_lo_12[113]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi_hi_1 = {regroupV0_lo_12[125], regroupV0_lo_12[121]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi_5 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi_hi_1, regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_9 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi_5, regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_lo_hi_12 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_9, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_9};
  wire [31:0]        regroupV0_lo_lo_lo_lo_lo_lo_12 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_12, regroupV0_lo_lo_lo_lo_lo_lo_lo_12};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo_lo_1 = {regroupV0_lo_12[133], regroupV0_lo_12[129]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo_hi_1 = {regroupV0_lo_12[141], regroupV0_lo_12[137]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo_5 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi_lo_1 = {regroupV0_lo_12[149], regroupV0_lo_12[145]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi_hi_1 = {regroupV0_lo_12[157], regroupV0_lo_12[153]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi_5 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi_hi_1, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_9 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi_5, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo_lo_1 = {regroupV0_lo_12[165], regroupV0_lo_12[161]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo_hi_1 = {regroupV0_lo_12[173], regroupV0_lo_12[169]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo_5 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo_hi_1, regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi_lo_1 = {regroupV0_lo_12[181], regroupV0_lo_12[177]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi_hi_1 = {regroupV0_lo_12[189], regroupV0_lo_12[185]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi_5 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi_hi_1, regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_9 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi_5, regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_hi_lo_12 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_9, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_9};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo_lo_1 = {regroupV0_lo_12[197], regroupV0_lo_12[193]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo_hi_1 = {regroupV0_lo_12[205], regroupV0_lo_12[201]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo_5 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi_lo_1 = {regroupV0_lo_12[213], regroupV0_lo_12[209]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi_hi_1 = {regroupV0_lo_12[221], regroupV0_lo_12[217]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi_5 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi_hi_1, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_9 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi_5, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo_lo_1 = {regroupV0_lo_12[229], regroupV0_lo_12[225]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo_hi_1 = {regroupV0_lo_12[237], regroupV0_lo_12[233]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo_5 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo_hi_1, regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi_lo_1 = {regroupV0_lo_12[245], regroupV0_lo_12[241]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi_hi_1 = {regroupV0_lo_12[253], regroupV0_lo_12[249]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi_5 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi_hi_1, regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_9 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi_5, regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_hi_hi_12 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_9, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_9};
  wire [31:0]        regroupV0_lo_lo_lo_lo_lo_hi_12 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_12, regroupV0_lo_lo_lo_lo_lo_hi_lo_12};
  wire [63:0]        regroupV0_lo_lo_lo_lo_lo_12 = {regroupV0_lo_lo_lo_lo_lo_hi_12, regroupV0_lo_lo_lo_lo_lo_lo_12};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo_lo_1 = {regroupV0_lo_12[261], regroupV0_lo_12[257]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo_hi_1 = {regroupV0_lo_12[269], regroupV0_lo_12[265]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo_5 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi_lo_1 = {regroupV0_lo_12[277], regroupV0_lo_12[273]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi_hi_1 = {regroupV0_lo_12[285], regroupV0_lo_12[281]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi_5 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi_hi_1, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_9 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi_5, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo_lo_1 = {regroupV0_lo_12[293], regroupV0_lo_12[289]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo_hi_1 = {regroupV0_lo_12[301], regroupV0_lo_12[297]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo_5 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo_hi_1, regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi_lo_1 = {regroupV0_lo_12[309], regroupV0_lo_12[305]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi_hi_1 = {regroupV0_lo_12[317], regroupV0_lo_12[313]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi_5 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi_hi_1, regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_9 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi_5, regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_lo_lo_12 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_9, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_9};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo_lo_1 = {regroupV0_lo_12[325], regroupV0_lo_12[321]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo_hi_1 = {regroupV0_lo_12[333], regroupV0_lo_12[329]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo_5 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi_lo_1 = {regroupV0_lo_12[341], regroupV0_lo_12[337]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi_hi_1 = {regroupV0_lo_12[349], regroupV0_lo_12[345]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi_5 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi_hi_1, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_9 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi_5, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo_lo_1 = {regroupV0_lo_12[357], regroupV0_lo_12[353]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo_hi_1 = {regroupV0_lo_12[365], regroupV0_lo_12[361]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo_5 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo_hi_1, regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi_lo_1 = {regroupV0_lo_12[373], regroupV0_lo_12[369]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi_hi_1 = {regroupV0_lo_12[381], regroupV0_lo_12[377]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi_5 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi_hi_1, regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_9 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi_5, regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_lo_hi_12 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_9, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_9};
  wire [31:0]        regroupV0_lo_lo_lo_lo_hi_lo_12 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_12, regroupV0_lo_lo_lo_lo_hi_lo_lo_12};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo_lo_1 = {regroupV0_lo_12[389], regroupV0_lo_12[385]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo_hi_1 = {regroupV0_lo_12[397], regroupV0_lo_12[393]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo_5 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi_lo_1 = {regroupV0_lo_12[405], regroupV0_lo_12[401]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi_hi_1 = {regroupV0_lo_12[413], regroupV0_lo_12[409]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi_5 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi_hi_1, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_9 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi_5, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo_lo_1 = {regroupV0_lo_12[421], regroupV0_lo_12[417]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo_hi_1 = {regroupV0_lo_12[429], regroupV0_lo_12[425]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo_5 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo_hi_1, regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi_lo_1 = {regroupV0_lo_12[437], regroupV0_lo_12[433]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi_hi_1 = {regroupV0_lo_12[445], regroupV0_lo_12[441]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi_5 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi_hi_1, regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_9 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi_5, regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_hi_lo_12 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_9, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_9};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo_lo_1 = {regroupV0_lo_12[453], regroupV0_lo_12[449]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo_hi_1 = {regroupV0_lo_12[461], regroupV0_lo_12[457]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo_5 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi_lo_1 = {regroupV0_lo_12[469], regroupV0_lo_12[465]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi_hi_1 = {regroupV0_lo_12[477], regroupV0_lo_12[473]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi_5 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi_hi_1, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_9 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi_5, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo_lo_1 = {regroupV0_lo_12[485], regroupV0_lo_12[481]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo_hi_1 = {regroupV0_lo_12[493], regroupV0_lo_12[489]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo_5 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo_hi_1, regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi_lo_1 = {regroupV0_lo_12[501], regroupV0_lo_12[497]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi_hi_1 = {regroupV0_lo_12[509], regroupV0_lo_12[505]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi_5 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi_hi_1, regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_9 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi_5, regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_hi_hi_12 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_9, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_9};
  wire [31:0]        regroupV0_lo_lo_lo_lo_hi_hi_12 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_12, regroupV0_lo_lo_lo_lo_hi_hi_lo_12};
  wire [63:0]        regroupV0_lo_lo_lo_lo_hi_12 = {regroupV0_lo_lo_lo_lo_hi_hi_12, regroupV0_lo_lo_lo_lo_hi_lo_12};
  wire [127:0]       regroupV0_lo_lo_lo_lo_12 = {regroupV0_lo_lo_lo_lo_hi_12, regroupV0_lo_lo_lo_lo_lo_12};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo_lo_1 = {regroupV0_lo_12[517], regroupV0_lo_12[513]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo_hi_1 = {regroupV0_lo_12[525], regroupV0_lo_12[521]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo_5 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi_lo_1 = {regroupV0_lo_12[533], regroupV0_lo_12[529]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi_hi_1 = {regroupV0_lo_12[541], regroupV0_lo_12[537]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi_5 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi_hi_1, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_9 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi_5, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo_lo_1 = {regroupV0_lo_12[549], regroupV0_lo_12[545]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo_hi_1 = {regroupV0_lo_12[557], regroupV0_lo_12[553]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo_5 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo_hi_1, regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi_lo_1 = {regroupV0_lo_12[565], regroupV0_lo_12[561]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi_hi_1 = {regroupV0_lo_12[573], regroupV0_lo_12[569]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi_5 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi_hi_1, regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_9 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi_5, regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_lo_lo_12 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_9, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_9};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo_lo_1 = {regroupV0_lo_12[581], regroupV0_lo_12[577]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo_hi_1 = {regroupV0_lo_12[589], regroupV0_lo_12[585]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo_5 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo_hi_1, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi_lo_1 = {regroupV0_lo_12[597], regroupV0_lo_12[593]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi_hi_1 = {regroupV0_lo_12[605], regroupV0_lo_12[601]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi_5 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi_hi_1, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_9 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi_5, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo_lo_1 = {regroupV0_lo_12[613], regroupV0_lo_12[609]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo_hi_1 = {regroupV0_lo_12[621], regroupV0_lo_12[617]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo_5 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo_hi_1, regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi_lo_1 = {regroupV0_lo_12[629], regroupV0_lo_12[625]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi_hi_1 = {regroupV0_lo_12[637], regroupV0_lo_12[633]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi_5 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi_hi_1, regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_9 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi_5, regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_lo_hi_12 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_9, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_9};
  wire [31:0]        regroupV0_lo_lo_lo_hi_lo_lo_12 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_12, regroupV0_lo_lo_lo_hi_lo_lo_lo_12};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo_lo_1 = {regroupV0_lo_12[645], regroupV0_lo_12[641]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo_hi_1 = {regroupV0_lo_12[653], regroupV0_lo_12[649]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo_5 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi_lo_1 = {regroupV0_lo_12[661], regroupV0_lo_12[657]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi_hi_1 = {regroupV0_lo_12[669], regroupV0_lo_12[665]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi_5 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi_hi_1, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_9 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi_5, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo_lo_1 = {regroupV0_lo_12[677], regroupV0_lo_12[673]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo_hi_1 = {regroupV0_lo_12[685], regroupV0_lo_12[681]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo_5 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo_hi_1, regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi_lo_1 = {regroupV0_lo_12[693], regroupV0_lo_12[689]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi_hi_1 = {regroupV0_lo_12[701], regroupV0_lo_12[697]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi_5 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi_hi_1, regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_9 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi_5, regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_hi_lo_12 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_9, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_9};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo_lo_1 = {regroupV0_lo_12[709], regroupV0_lo_12[705]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo_hi_1 = {regroupV0_lo_12[717], regroupV0_lo_12[713]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo_5 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo_hi_1, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi_lo_1 = {regroupV0_lo_12[725], regroupV0_lo_12[721]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi_hi_1 = {regroupV0_lo_12[733], regroupV0_lo_12[729]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi_5 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi_hi_1, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_9 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi_5, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo_lo_1 = {regroupV0_lo_12[741], regroupV0_lo_12[737]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo_hi_1 = {regroupV0_lo_12[749], regroupV0_lo_12[745]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo_5 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo_hi_1, regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi_lo_1 = {regroupV0_lo_12[757], regroupV0_lo_12[753]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi_hi_1 = {regroupV0_lo_12[765], regroupV0_lo_12[761]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi_5 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi_hi_1, regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_9 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi_5, regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_hi_hi_12 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_9, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_9};
  wire [31:0]        regroupV0_lo_lo_lo_hi_lo_hi_12 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_12, regroupV0_lo_lo_lo_hi_lo_hi_lo_12};
  wire [63:0]        regroupV0_lo_lo_lo_hi_lo_12 = {regroupV0_lo_lo_lo_hi_lo_hi_12, regroupV0_lo_lo_lo_hi_lo_lo_12};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo_lo_1 = {regroupV0_lo_12[773], regroupV0_lo_12[769]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo_hi_1 = {regroupV0_lo_12[781], regroupV0_lo_12[777]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo_5 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi_lo_1 = {regroupV0_lo_12[789], regroupV0_lo_12[785]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi_hi_1 = {regroupV0_lo_12[797], regroupV0_lo_12[793]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi_5 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi_hi_1, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_9 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi_5, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo_lo_1 = {regroupV0_lo_12[805], regroupV0_lo_12[801]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo_hi_1 = {regroupV0_lo_12[813], regroupV0_lo_12[809]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo_5 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo_hi_1, regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi_lo_1 = {regroupV0_lo_12[821], regroupV0_lo_12[817]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi_hi_1 = {regroupV0_lo_12[829], regroupV0_lo_12[825]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi_5 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi_hi_1, regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_9 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi_5, regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_lo_lo_12 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_9, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_9};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo_lo_1 = {regroupV0_lo_12[837], regroupV0_lo_12[833]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo_hi_1 = {regroupV0_lo_12[845], regroupV0_lo_12[841]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo_5 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo_hi_1, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi_lo_1 = {regroupV0_lo_12[853], regroupV0_lo_12[849]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi_hi_1 = {regroupV0_lo_12[861], regroupV0_lo_12[857]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi_5 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi_hi_1, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_9 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi_5, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo_lo_1 = {regroupV0_lo_12[869], regroupV0_lo_12[865]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo_hi_1 = {regroupV0_lo_12[877], regroupV0_lo_12[873]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo_5 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo_hi_1, regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi_lo_1 = {regroupV0_lo_12[885], regroupV0_lo_12[881]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi_hi_1 = {regroupV0_lo_12[893], regroupV0_lo_12[889]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi_5 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi_hi_1, regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_9 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi_5, regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_lo_hi_12 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_9, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_9};
  wire [31:0]        regroupV0_lo_lo_lo_hi_hi_lo_12 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_12, regroupV0_lo_lo_lo_hi_hi_lo_lo_12};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo_lo_1 = {regroupV0_lo_12[901], regroupV0_lo_12[897]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo_hi_1 = {regroupV0_lo_12[909], regroupV0_lo_12[905]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo_5 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi_lo_1 = {regroupV0_lo_12[917], regroupV0_lo_12[913]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi_hi_1 = {regroupV0_lo_12[925], regroupV0_lo_12[921]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi_5 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi_hi_1, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_9 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi_5, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo_lo_1 = {regroupV0_lo_12[933], regroupV0_lo_12[929]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo_hi_1 = {regroupV0_lo_12[941], regroupV0_lo_12[937]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo_5 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo_hi_1, regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi_lo_1 = {regroupV0_lo_12[949], regroupV0_lo_12[945]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi_hi_1 = {regroupV0_lo_12[957], regroupV0_lo_12[953]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi_5 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi_hi_1, regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_9 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi_5, regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_hi_lo_12 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_9, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_9};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo_lo_1 = {regroupV0_lo_12[965], regroupV0_lo_12[961]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo_hi_1 = {regroupV0_lo_12[973], regroupV0_lo_12[969]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo_5 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo_hi_1, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi_lo_1 = {regroupV0_lo_12[981], regroupV0_lo_12[977]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi_hi_1 = {regroupV0_lo_12[989], regroupV0_lo_12[985]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi_5 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi_hi_1, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_9 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi_5, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo_lo_1 = {regroupV0_lo_12[997], regroupV0_lo_12[993]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo_hi_1 = {regroupV0_lo_12[1005], regroupV0_lo_12[1001]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo_5 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo_hi_1, regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi_lo_1 = {regroupV0_lo_12[1013], regroupV0_lo_12[1009]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi_hi_1 = {regroupV0_lo_12[1021], regroupV0_lo_12[1017]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi_5 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi_hi_1, regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_9 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi_5, regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_hi_hi_12 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_9, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_9};
  wire [31:0]        regroupV0_lo_lo_lo_hi_hi_hi_12 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_12, regroupV0_lo_lo_lo_hi_hi_hi_lo_12};
  wire [63:0]        regroupV0_lo_lo_lo_hi_hi_12 = {regroupV0_lo_lo_lo_hi_hi_hi_12, regroupV0_lo_lo_lo_hi_hi_lo_12};
  wire [127:0]       regroupV0_lo_lo_lo_hi_12 = {regroupV0_lo_lo_lo_hi_hi_12, regroupV0_lo_lo_lo_hi_lo_12};
  wire [255:0]       regroupV0_lo_lo_lo_12 = {regroupV0_lo_lo_lo_hi_12, regroupV0_lo_lo_lo_lo_12};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo_lo_1 = {regroupV0_lo_12[1029], regroupV0_lo_12[1025]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo_hi_1 = {regroupV0_lo_12[1037], regroupV0_lo_12[1033]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo_5 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo_hi_1, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi_lo_1 = {regroupV0_lo_12[1045], regroupV0_lo_12[1041]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi_hi_1 = {regroupV0_lo_12[1053], regroupV0_lo_12[1049]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi_5 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi_hi_1, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_9 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi_5, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo_lo_1 = {regroupV0_lo_12[1061], regroupV0_lo_12[1057]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo_hi_1 = {regroupV0_lo_12[1069], regroupV0_lo_12[1065]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo_5 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo_hi_1, regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi_lo_1 = {regroupV0_lo_12[1077], regroupV0_lo_12[1073]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi_hi_1 = {regroupV0_lo_12[1085], regroupV0_lo_12[1081]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi_5 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi_hi_1, regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_9 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi_5, regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_lo_lo_12 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_9, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_9};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo_lo_1 = {regroupV0_lo_12[1093], regroupV0_lo_12[1089]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo_hi_1 = {regroupV0_lo_12[1101], regroupV0_lo_12[1097]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo_5 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo_hi_1, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi_lo_1 = {regroupV0_lo_12[1109], regroupV0_lo_12[1105]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi_hi_1 = {regroupV0_lo_12[1117], regroupV0_lo_12[1113]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi_5 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi_hi_1, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_9 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi_5, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo_lo_1 = {regroupV0_lo_12[1125], regroupV0_lo_12[1121]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo_hi_1 = {regroupV0_lo_12[1133], regroupV0_lo_12[1129]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo_5 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo_hi_1, regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi_lo_1 = {regroupV0_lo_12[1141], regroupV0_lo_12[1137]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi_hi_1 = {regroupV0_lo_12[1149], regroupV0_lo_12[1145]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi_5 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi_hi_1, regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_9 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi_5, regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_lo_hi_12 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_9, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_9};
  wire [31:0]        regroupV0_lo_lo_hi_lo_lo_lo_12 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_12, regroupV0_lo_lo_hi_lo_lo_lo_lo_12};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo_lo_1 = {regroupV0_lo_12[1157], regroupV0_lo_12[1153]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo_hi_1 = {regroupV0_lo_12[1165], regroupV0_lo_12[1161]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo_5 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo_hi_1, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi_lo_1 = {regroupV0_lo_12[1173], regroupV0_lo_12[1169]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi_hi_1 = {regroupV0_lo_12[1181], regroupV0_lo_12[1177]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi_5 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi_hi_1, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_9 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi_5, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo_lo_1 = {regroupV0_lo_12[1189], regroupV0_lo_12[1185]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo_hi_1 = {regroupV0_lo_12[1197], regroupV0_lo_12[1193]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo_5 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo_hi_1, regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi_lo_1 = {regroupV0_lo_12[1205], regroupV0_lo_12[1201]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi_hi_1 = {regroupV0_lo_12[1213], regroupV0_lo_12[1209]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi_5 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi_hi_1, regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_9 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi_5, regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_hi_lo_12 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_9, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_9};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo_lo_1 = {regroupV0_lo_12[1221], regroupV0_lo_12[1217]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo_hi_1 = {regroupV0_lo_12[1229], regroupV0_lo_12[1225]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo_5 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo_hi_1, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi_lo_1 = {regroupV0_lo_12[1237], regroupV0_lo_12[1233]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi_hi_1 = {regroupV0_lo_12[1245], regroupV0_lo_12[1241]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi_5 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi_hi_1, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_9 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi_5, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo_lo_1 = {regroupV0_lo_12[1253], regroupV0_lo_12[1249]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo_hi_1 = {regroupV0_lo_12[1261], regroupV0_lo_12[1257]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo_5 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo_hi_1, regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi_lo_1 = {regroupV0_lo_12[1269], regroupV0_lo_12[1265]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi_hi_1 = {regroupV0_lo_12[1277], regroupV0_lo_12[1273]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi_5 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi_hi_1, regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_9 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi_5, regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_hi_hi_12 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_9, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_9};
  wire [31:0]        regroupV0_lo_lo_hi_lo_lo_hi_12 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_12, regroupV0_lo_lo_hi_lo_lo_hi_lo_12};
  wire [63:0]        regroupV0_lo_lo_hi_lo_lo_12 = {regroupV0_lo_lo_hi_lo_lo_hi_12, regroupV0_lo_lo_hi_lo_lo_lo_12};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo_lo_1 = {regroupV0_lo_12[1285], regroupV0_lo_12[1281]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo_hi_1 = {regroupV0_lo_12[1293], regroupV0_lo_12[1289]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo_5 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo_hi_1, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi_lo_1 = {regroupV0_lo_12[1301], regroupV0_lo_12[1297]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi_hi_1 = {regroupV0_lo_12[1309], regroupV0_lo_12[1305]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi_5 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi_hi_1, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_9 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi_5, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo_lo_1 = {regroupV0_lo_12[1317], regroupV0_lo_12[1313]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo_hi_1 = {regroupV0_lo_12[1325], regroupV0_lo_12[1321]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo_5 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo_hi_1, regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi_lo_1 = {regroupV0_lo_12[1333], regroupV0_lo_12[1329]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi_hi_1 = {regroupV0_lo_12[1341], regroupV0_lo_12[1337]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi_5 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi_hi_1, regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_9 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi_5, regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_lo_lo_12 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_9, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_9};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo_lo_1 = {regroupV0_lo_12[1349], regroupV0_lo_12[1345]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo_hi_1 = {regroupV0_lo_12[1357], regroupV0_lo_12[1353]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo_5 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo_hi_1, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi_lo_1 = {regroupV0_lo_12[1365], regroupV0_lo_12[1361]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi_hi_1 = {regroupV0_lo_12[1373], regroupV0_lo_12[1369]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi_5 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi_hi_1, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_9 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi_5, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo_lo_1 = {regroupV0_lo_12[1381], regroupV0_lo_12[1377]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo_hi_1 = {regroupV0_lo_12[1389], regroupV0_lo_12[1385]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo_5 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo_hi_1, regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi_lo_1 = {regroupV0_lo_12[1397], regroupV0_lo_12[1393]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi_hi_1 = {regroupV0_lo_12[1405], regroupV0_lo_12[1401]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi_5 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi_hi_1, regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_9 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi_5, regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_lo_hi_12 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_9, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_9};
  wire [31:0]        regroupV0_lo_lo_hi_lo_hi_lo_12 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_12, regroupV0_lo_lo_hi_lo_hi_lo_lo_12};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo_lo_1 = {regroupV0_lo_12[1413], regroupV0_lo_12[1409]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo_hi_1 = {regroupV0_lo_12[1421], regroupV0_lo_12[1417]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo_5 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo_hi_1, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi_lo_1 = {regroupV0_lo_12[1429], regroupV0_lo_12[1425]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi_hi_1 = {regroupV0_lo_12[1437], regroupV0_lo_12[1433]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi_5 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi_hi_1, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_9 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi_5, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo_lo_1 = {regroupV0_lo_12[1445], regroupV0_lo_12[1441]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo_hi_1 = {regroupV0_lo_12[1453], regroupV0_lo_12[1449]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo_5 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo_hi_1, regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi_lo_1 = {regroupV0_lo_12[1461], regroupV0_lo_12[1457]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi_hi_1 = {regroupV0_lo_12[1469], regroupV0_lo_12[1465]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi_5 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi_hi_1, regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_9 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi_5, regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_hi_lo_12 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_9, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_9};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo_lo_1 = {regroupV0_lo_12[1477], regroupV0_lo_12[1473]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo_hi_1 = {regroupV0_lo_12[1485], regroupV0_lo_12[1481]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo_5 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo_hi_1, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi_lo_1 = {regroupV0_lo_12[1493], regroupV0_lo_12[1489]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi_hi_1 = {regroupV0_lo_12[1501], regroupV0_lo_12[1497]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi_5 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi_hi_1, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_9 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi_5, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo_lo_1 = {regroupV0_lo_12[1509], regroupV0_lo_12[1505]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo_hi_1 = {regroupV0_lo_12[1517], regroupV0_lo_12[1513]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo_5 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo_hi_1, regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi_lo_1 = {regroupV0_lo_12[1525], regroupV0_lo_12[1521]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi_hi_1 = {regroupV0_lo_12[1533], regroupV0_lo_12[1529]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi_5 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi_hi_1, regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_9 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi_5, regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_hi_hi_12 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_9, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_9};
  wire [31:0]        regroupV0_lo_lo_hi_lo_hi_hi_12 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_12, regroupV0_lo_lo_hi_lo_hi_hi_lo_12};
  wire [63:0]        regroupV0_lo_lo_hi_lo_hi_12 = {regroupV0_lo_lo_hi_lo_hi_hi_12, regroupV0_lo_lo_hi_lo_hi_lo_12};
  wire [127:0]       regroupV0_lo_lo_hi_lo_12 = {regroupV0_lo_lo_hi_lo_hi_12, regroupV0_lo_lo_hi_lo_lo_12};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo_lo_1 = {regroupV0_lo_12[1541], regroupV0_lo_12[1537]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo_hi_1 = {regroupV0_lo_12[1549], regroupV0_lo_12[1545]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo_5 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo_hi_1, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi_lo_1 = {regroupV0_lo_12[1557], regroupV0_lo_12[1553]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi_hi_1 = {regroupV0_lo_12[1565], regroupV0_lo_12[1561]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi_5 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi_hi_1, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_9 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi_5, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo_lo_1 = {regroupV0_lo_12[1573], regroupV0_lo_12[1569]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo_hi_1 = {regroupV0_lo_12[1581], regroupV0_lo_12[1577]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo_5 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo_hi_1, regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi_lo_1 = {regroupV0_lo_12[1589], regroupV0_lo_12[1585]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi_hi_1 = {regroupV0_lo_12[1597], regroupV0_lo_12[1593]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi_5 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi_hi_1, regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_9 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi_5, regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_lo_lo_12 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_9, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_9};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo_lo_1 = {regroupV0_lo_12[1605], regroupV0_lo_12[1601]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo_hi_1 = {regroupV0_lo_12[1613], regroupV0_lo_12[1609]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo_5 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo_hi_1, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi_lo_1 = {regroupV0_lo_12[1621], regroupV0_lo_12[1617]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi_hi_1 = {regroupV0_lo_12[1629], regroupV0_lo_12[1625]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi_5 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi_hi_1, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_9 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi_5, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo_lo_1 = {regroupV0_lo_12[1637], regroupV0_lo_12[1633]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo_hi_1 = {regroupV0_lo_12[1645], regroupV0_lo_12[1641]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo_5 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo_hi_1, regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi_lo_1 = {regroupV0_lo_12[1653], regroupV0_lo_12[1649]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi_hi_1 = {regroupV0_lo_12[1661], regroupV0_lo_12[1657]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi_5 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi_hi_1, regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_9 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi_5, regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_lo_hi_12 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_9, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_9};
  wire [31:0]        regroupV0_lo_lo_hi_hi_lo_lo_12 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_12, regroupV0_lo_lo_hi_hi_lo_lo_lo_12};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo_lo_1 = {regroupV0_lo_12[1669], regroupV0_lo_12[1665]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo_hi_1 = {regroupV0_lo_12[1677], regroupV0_lo_12[1673]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo_5 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo_hi_1, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi_lo_1 = {regroupV0_lo_12[1685], regroupV0_lo_12[1681]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi_hi_1 = {regroupV0_lo_12[1693], regroupV0_lo_12[1689]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi_5 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi_hi_1, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_9 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi_5, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo_lo_1 = {regroupV0_lo_12[1701], regroupV0_lo_12[1697]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo_hi_1 = {regroupV0_lo_12[1709], regroupV0_lo_12[1705]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo_5 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo_hi_1, regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi_lo_1 = {regroupV0_lo_12[1717], regroupV0_lo_12[1713]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi_hi_1 = {regroupV0_lo_12[1725], regroupV0_lo_12[1721]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi_5 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi_hi_1, regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_9 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi_5, regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_hi_lo_12 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_9, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_9};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo_lo_1 = {regroupV0_lo_12[1733], regroupV0_lo_12[1729]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo_hi_1 = {regroupV0_lo_12[1741], regroupV0_lo_12[1737]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo_5 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo_hi_1, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi_lo_1 = {regroupV0_lo_12[1749], regroupV0_lo_12[1745]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi_hi_1 = {regroupV0_lo_12[1757], regroupV0_lo_12[1753]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi_5 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi_hi_1, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_9 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi_5, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo_lo_1 = {regroupV0_lo_12[1765], regroupV0_lo_12[1761]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo_hi_1 = {regroupV0_lo_12[1773], regroupV0_lo_12[1769]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo_5 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo_hi_1, regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi_lo_1 = {regroupV0_lo_12[1781], regroupV0_lo_12[1777]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi_hi_1 = {regroupV0_lo_12[1789], regroupV0_lo_12[1785]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi_5 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi_hi_1, regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_9 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi_5, regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_hi_hi_12 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_9, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_9};
  wire [31:0]        regroupV0_lo_lo_hi_hi_lo_hi_12 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_12, regroupV0_lo_lo_hi_hi_lo_hi_lo_12};
  wire [63:0]        regroupV0_lo_lo_hi_hi_lo_12 = {regroupV0_lo_lo_hi_hi_lo_hi_12, regroupV0_lo_lo_hi_hi_lo_lo_12};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo_lo_1 = {regroupV0_lo_12[1797], regroupV0_lo_12[1793]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo_hi_1 = {regroupV0_lo_12[1805], regroupV0_lo_12[1801]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo_5 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo_hi_1, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi_lo_1 = {regroupV0_lo_12[1813], regroupV0_lo_12[1809]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi_hi_1 = {regroupV0_lo_12[1821], regroupV0_lo_12[1817]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi_5 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi_hi_1, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_9 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi_5, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo_lo_1 = {regroupV0_lo_12[1829], regroupV0_lo_12[1825]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo_hi_1 = {regroupV0_lo_12[1837], regroupV0_lo_12[1833]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo_5 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo_hi_1, regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi_lo_1 = {regroupV0_lo_12[1845], regroupV0_lo_12[1841]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi_hi_1 = {regroupV0_lo_12[1853], regroupV0_lo_12[1849]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi_5 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi_hi_1, regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_9 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi_5, regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_lo_lo_12 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_9, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_9};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo_lo_1 = {regroupV0_lo_12[1861], regroupV0_lo_12[1857]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo_hi_1 = {regroupV0_lo_12[1869], regroupV0_lo_12[1865]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo_5 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo_hi_1, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi_lo_1 = {regroupV0_lo_12[1877], regroupV0_lo_12[1873]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi_hi_1 = {regroupV0_lo_12[1885], regroupV0_lo_12[1881]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi_5 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi_hi_1, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_9 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi_5, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo_lo_1 = {regroupV0_lo_12[1893], regroupV0_lo_12[1889]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo_hi_1 = {regroupV0_lo_12[1901], regroupV0_lo_12[1897]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo_5 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo_hi_1, regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi_lo_1 = {regroupV0_lo_12[1909], regroupV0_lo_12[1905]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi_hi_1 = {regroupV0_lo_12[1917], regroupV0_lo_12[1913]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi_5 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi_hi_1, regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_9 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi_5, regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_lo_hi_12 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_9, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_9};
  wire [31:0]        regroupV0_lo_lo_hi_hi_hi_lo_12 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_12, regroupV0_lo_lo_hi_hi_hi_lo_lo_12};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo_lo_1 = {regroupV0_lo_12[1925], regroupV0_lo_12[1921]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo_hi_1 = {regroupV0_lo_12[1933], regroupV0_lo_12[1929]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo_5 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo_hi_1, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi_lo_1 = {regroupV0_lo_12[1941], regroupV0_lo_12[1937]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi_hi_1 = {regroupV0_lo_12[1949], regroupV0_lo_12[1945]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi_5 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi_hi_1, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_9 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi_5, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo_lo_1 = {regroupV0_lo_12[1957], regroupV0_lo_12[1953]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo_hi_1 = {regroupV0_lo_12[1965], regroupV0_lo_12[1961]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo_5 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo_hi_1, regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi_lo_1 = {regroupV0_lo_12[1973], regroupV0_lo_12[1969]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi_hi_1 = {regroupV0_lo_12[1981], regroupV0_lo_12[1977]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi_5 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi_hi_1, regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_9 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi_5, regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_hi_lo_12 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_9, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_9};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo_lo_1 = {regroupV0_lo_12[1989], regroupV0_lo_12[1985]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo_hi_1 = {regroupV0_lo_12[1997], regroupV0_lo_12[1993]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo_5 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo_hi_1, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi_lo_1 = {regroupV0_lo_12[2005], regroupV0_lo_12[2001]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi_hi_1 = {regroupV0_lo_12[2013], regroupV0_lo_12[2009]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi_5 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi_hi_1, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_9 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi_5, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo_lo_1 = {regroupV0_lo_12[2021], regroupV0_lo_12[2017]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo_hi_1 = {regroupV0_lo_12[2029], regroupV0_lo_12[2025]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo_5 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo_hi_1, regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi_lo_1 = {regroupV0_lo_12[2037], regroupV0_lo_12[2033]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi_hi_1 = {regroupV0_lo_12[2045], regroupV0_lo_12[2041]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi_5 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi_hi_1, regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_9 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi_5, regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_hi_hi_12 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_9, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_9};
  wire [31:0]        regroupV0_lo_lo_hi_hi_hi_hi_12 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_12, regroupV0_lo_lo_hi_hi_hi_hi_lo_12};
  wire [63:0]        regroupV0_lo_lo_hi_hi_hi_12 = {regroupV0_lo_lo_hi_hi_hi_hi_12, regroupV0_lo_lo_hi_hi_hi_lo_12};
  wire [127:0]       regroupV0_lo_lo_hi_hi_12 = {regroupV0_lo_lo_hi_hi_hi_12, regroupV0_lo_lo_hi_hi_lo_12};
  wire [255:0]       regroupV0_lo_lo_hi_12 = {regroupV0_lo_lo_hi_hi_12, regroupV0_lo_lo_hi_lo_12};
  wire [511:0]       regroupV0_lo_lo_12 = {regroupV0_lo_lo_hi_12, regroupV0_lo_lo_lo_12};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo_lo_1 = {regroupV0_lo_12[2053], regroupV0_lo_12[2049]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo_hi_1 = {regroupV0_lo_12[2061], regroupV0_lo_12[2057]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo_5 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo_hi_1, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi_lo_1 = {regroupV0_lo_12[2069], regroupV0_lo_12[2065]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi_hi_1 = {regroupV0_lo_12[2077], regroupV0_lo_12[2073]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi_5 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi_hi_1, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_9 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi_5, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo_lo_1 = {regroupV0_lo_12[2085], regroupV0_lo_12[2081]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo_hi_1 = {regroupV0_lo_12[2093], regroupV0_lo_12[2089]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo_5 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo_hi_1, regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi_lo_1 = {regroupV0_lo_12[2101], regroupV0_lo_12[2097]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi_hi_1 = {regroupV0_lo_12[2109], regroupV0_lo_12[2105]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi_5 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi_hi_1, regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_9 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi_5, regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_lo_lo_12 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_9, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_9};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo_lo_1 = {regroupV0_lo_12[2117], regroupV0_lo_12[2113]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo_hi_1 = {regroupV0_lo_12[2125], regroupV0_lo_12[2121]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo_5 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo_hi_1, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi_lo_1 = {regroupV0_lo_12[2133], regroupV0_lo_12[2129]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi_hi_1 = {regroupV0_lo_12[2141], regroupV0_lo_12[2137]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi_5 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi_hi_1, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_9 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi_5, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo_lo_1 = {regroupV0_lo_12[2149], regroupV0_lo_12[2145]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo_hi_1 = {regroupV0_lo_12[2157], regroupV0_lo_12[2153]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo_5 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo_hi_1, regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi_lo_1 = {regroupV0_lo_12[2165], regroupV0_lo_12[2161]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi_hi_1 = {regroupV0_lo_12[2173], regroupV0_lo_12[2169]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi_5 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi_hi_1, regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_9 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi_5, regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_lo_hi_12 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_9, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_9};
  wire [31:0]        regroupV0_lo_hi_lo_lo_lo_lo_12 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_12, regroupV0_lo_hi_lo_lo_lo_lo_lo_12};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo_lo_1 = {regroupV0_lo_12[2181], regroupV0_lo_12[2177]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo_hi_1 = {regroupV0_lo_12[2189], regroupV0_lo_12[2185]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo_5 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo_hi_1, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi_lo_1 = {regroupV0_lo_12[2197], regroupV0_lo_12[2193]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi_hi_1 = {regroupV0_lo_12[2205], regroupV0_lo_12[2201]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi_5 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi_hi_1, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_9 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi_5, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo_lo_1 = {regroupV0_lo_12[2213], regroupV0_lo_12[2209]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo_hi_1 = {regroupV0_lo_12[2221], regroupV0_lo_12[2217]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo_5 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo_hi_1, regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi_lo_1 = {regroupV0_lo_12[2229], regroupV0_lo_12[2225]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi_hi_1 = {regroupV0_lo_12[2237], regroupV0_lo_12[2233]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi_5 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi_hi_1, regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_9 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi_5, regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_hi_lo_12 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_9, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_9};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo_lo_1 = {regroupV0_lo_12[2245], regroupV0_lo_12[2241]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo_hi_1 = {regroupV0_lo_12[2253], regroupV0_lo_12[2249]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo_5 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo_hi_1, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi_lo_1 = {regroupV0_lo_12[2261], regroupV0_lo_12[2257]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi_hi_1 = {regroupV0_lo_12[2269], regroupV0_lo_12[2265]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi_5 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi_hi_1, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_9 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi_5, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo_lo_1 = {regroupV0_lo_12[2277], regroupV0_lo_12[2273]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo_hi_1 = {regroupV0_lo_12[2285], regroupV0_lo_12[2281]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo_5 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo_hi_1, regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi_lo_1 = {regroupV0_lo_12[2293], regroupV0_lo_12[2289]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi_hi_1 = {regroupV0_lo_12[2301], regroupV0_lo_12[2297]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi_5 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi_hi_1, regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_9 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi_5, regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_hi_hi_12 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_9, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_9};
  wire [31:0]        regroupV0_lo_hi_lo_lo_lo_hi_12 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_12, regroupV0_lo_hi_lo_lo_lo_hi_lo_12};
  wire [63:0]        regroupV0_lo_hi_lo_lo_lo_12 = {regroupV0_lo_hi_lo_lo_lo_hi_12, regroupV0_lo_hi_lo_lo_lo_lo_12};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo_lo_1 = {regroupV0_lo_12[2309], regroupV0_lo_12[2305]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo_hi_1 = {regroupV0_lo_12[2317], regroupV0_lo_12[2313]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo_5 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo_hi_1, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi_lo_1 = {regroupV0_lo_12[2325], regroupV0_lo_12[2321]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi_hi_1 = {regroupV0_lo_12[2333], regroupV0_lo_12[2329]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi_5 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi_hi_1, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_9 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi_5, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo_lo_1 = {regroupV0_lo_12[2341], regroupV0_lo_12[2337]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo_hi_1 = {regroupV0_lo_12[2349], regroupV0_lo_12[2345]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo_5 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo_hi_1, regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi_lo_1 = {regroupV0_lo_12[2357], regroupV0_lo_12[2353]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi_hi_1 = {regroupV0_lo_12[2365], regroupV0_lo_12[2361]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi_5 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi_hi_1, regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_9 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi_5, regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_lo_lo_12 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_9, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_9};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo_lo_1 = {regroupV0_lo_12[2373], regroupV0_lo_12[2369]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo_hi_1 = {regroupV0_lo_12[2381], regroupV0_lo_12[2377]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo_5 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo_hi_1, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi_lo_1 = {regroupV0_lo_12[2389], regroupV0_lo_12[2385]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi_hi_1 = {regroupV0_lo_12[2397], regroupV0_lo_12[2393]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi_5 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi_hi_1, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_9 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi_5, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo_lo_1 = {regroupV0_lo_12[2405], regroupV0_lo_12[2401]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo_hi_1 = {regroupV0_lo_12[2413], regroupV0_lo_12[2409]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo_5 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo_hi_1, regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi_lo_1 = {regroupV0_lo_12[2421], regroupV0_lo_12[2417]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi_hi_1 = {regroupV0_lo_12[2429], regroupV0_lo_12[2425]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi_5 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi_hi_1, regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_9 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi_5, regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_lo_hi_12 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_9, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_9};
  wire [31:0]        regroupV0_lo_hi_lo_lo_hi_lo_12 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_12, regroupV0_lo_hi_lo_lo_hi_lo_lo_12};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo_lo_1 = {regroupV0_lo_12[2437], regroupV0_lo_12[2433]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo_hi_1 = {regroupV0_lo_12[2445], regroupV0_lo_12[2441]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo_5 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo_hi_1, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi_lo_1 = {regroupV0_lo_12[2453], regroupV0_lo_12[2449]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi_hi_1 = {regroupV0_lo_12[2461], regroupV0_lo_12[2457]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi_5 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi_hi_1, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_9 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi_5, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo_lo_1 = {regroupV0_lo_12[2469], regroupV0_lo_12[2465]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo_hi_1 = {regroupV0_lo_12[2477], regroupV0_lo_12[2473]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo_5 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo_hi_1, regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi_lo_1 = {regroupV0_lo_12[2485], regroupV0_lo_12[2481]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi_hi_1 = {regroupV0_lo_12[2493], regroupV0_lo_12[2489]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi_5 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi_hi_1, regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_9 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi_5, regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_hi_lo_12 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_9, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_9};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo_lo_1 = {regroupV0_lo_12[2501], regroupV0_lo_12[2497]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo_hi_1 = {regroupV0_lo_12[2509], regroupV0_lo_12[2505]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo_5 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo_hi_1, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi_lo_1 = {regroupV0_lo_12[2517], regroupV0_lo_12[2513]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi_hi_1 = {regroupV0_lo_12[2525], regroupV0_lo_12[2521]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi_5 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi_hi_1, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_9 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi_5, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo_lo_1 = {regroupV0_lo_12[2533], regroupV0_lo_12[2529]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo_hi_1 = {regroupV0_lo_12[2541], regroupV0_lo_12[2537]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo_5 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo_hi_1, regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi_lo_1 = {regroupV0_lo_12[2549], regroupV0_lo_12[2545]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi_hi_1 = {regroupV0_lo_12[2557], regroupV0_lo_12[2553]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi_5 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi_hi_1, regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_9 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi_5, regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_hi_hi_12 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_9, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_9};
  wire [31:0]        regroupV0_lo_hi_lo_lo_hi_hi_12 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_12, regroupV0_lo_hi_lo_lo_hi_hi_lo_12};
  wire [63:0]        regroupV0_lo_hi_lo_lo_hi_12 = {regroupV0_lo_hi_lo_lo_hi_hi_12, regroupV0_lo_hi_lo_lo_hi_lo_12};
  wire [127:0]       regroupV0_lo_hi_lo_lo_12 = {regroupV0_lo_hi_lo_lo_hi_12, regroupV0_lo_hi_lo_lo_lo_12};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo_lo_1 = {regroupV0_lo_12[2565], regroupV0_lo_12[2561]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo_hi_1 = {regroupV0_lo_12[2573], regroupV0_lo_12[2569]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo_5 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo_hi_1, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi_lo_1 = {regroupV0_lo_12[2581], regroupV0_lo_12[2577]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi_hi_1 = {regroupV0_lo_12[2589], regroupV0_lo_12[2585]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi_5 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi_hi_1, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_9 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi_5, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo_lo_1 = {regroupV0_lo_12[2597], regroupV0_lo_12[2593]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo_hi_1 = {regroupV0_lo_12[2605], regroupV0_lo_12[2601]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo_5 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo_hi_1, regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi_lo_1 = {regroupV0_lo_12[2613], regroupV0_lo_12[2609]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi_hi_1 = {regroupV0_lo_12[2621], regroupV0_lo_12[2617]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi_5 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi_hi_1, regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_9 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi_5, regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_lo_lo_12 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_9, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_9};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo_lo_1 = {regroupV0_lo_12[2629], regroupV0_lo_12[2625]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo_hi_1 = {regroupV0_lo_12[2637], regroupV0_lo_12[2633]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo_5 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo_hi_1, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi_lo_1 = {regroupV0_lo_12[2645], regroupV0_lo_12[2641]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi_hi_1 = {regroupV0_lo_12[2653], regroupV0_lo_12[2649]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi_5 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi_hi_1, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_9 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi_5, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo_lo_1 = {regroupV0_lo_12[2661], regroupV0_lo_12[2657]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo_hi_1 = {regroupV0_lo_12[2669], regroupV0_lo_12[2665]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo_5 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo_hi_1, regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi_lo_1 = {regroupV0_lo_12[2677], regroupV0_lo_12[2673]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi_hi_1 = {regroupV0_lo_12[2685], regroupV0_lo_12[2681]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi_5 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi_hi_1, regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_9 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi_5, regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_lo_hi_12 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_9, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_9};
  wire [31:0]        regroupV0_lo_hi_lo_hi_lo_lo_12 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_12, regroupV0_lo_hi_lo_hi_lo_lo_lo_12};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo_lo_1 = {regroupV0_lo_12[2693], regroupV0_lo_12[2689]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo_hi_1 = {regroupV0_lo_12[2701], regroupV0_lo_12[2697]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo_5 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo_hi_1, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi_lo_1 = {regroupV0_lo_12[2709], regroupV0_lo_12[2705]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi_hi_1 = {regroupV0_lo_12[2717], regroupV0_lo_12[2713]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi_5 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi_hi_1, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_9 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi_5, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo_lo_1 = {regroupV0_lo_12[2725], regroupV0_lo_12[2721]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo_hi_1 = {regroupV0_lo_12[2733], regroupV0_lo_12[2729]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo_5 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo_hi_1, regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi_lo_1 = {regroupV0_lo_12[2741], regroupV0_lo_12[2737]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi_hi_1 = {regroupV0_lo_12[2749], regroupV0_lo_12[2745]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi_5 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi_hi_1, regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_9 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi_5, regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_hi_lo_12 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_9, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_9};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo_lo_1 = {regroupV0_lo_12[2757], regroupV0_lo_12[2753]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo_hi_1 = {regroupV0_lo_12[2765], regroupV0_lo_12[2761]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo_5 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo_hi_1, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi_lo_1 = {regroupV0_lo_12[2773], regroupV0_lo_12[2769]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi_hi_1 = {regroupV0_lo_12[2781], regroupV0_lo_12[2777]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi_5 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi_hi_1, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_9 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi_5, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo_lo_1 = {regroupV0_lo_12[2789], regroupV0_lo_12[2785]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo_hi_1 = {regroupV0_lo_12[2797], regroupV0_lo_12[2793]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo_5 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo_hi_1, regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi_lo_1 = {regroupV0_lo_12[2805], regroupV0_lo_12[2801]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi_hi_1 = {regroupV0_lo_12[2813], regroupV0_lo_12[2809]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi_5 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi_hi_1, regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_9 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi_5, regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_hi_hi_12 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_9, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_9};
  wire [31:0]        regroupV0_lo_hi_lo_hi_lo_hi_12 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_12, regroupV0_lo_hi_lo_hi_lo_hi_lo_12};
  wire [63:0]        regroupV0_lo_hi_lo_hi_lo_12 = {regroupV0_lo_hi_lo_hi_lo_hi_12, regroupV0_lo_hi_lo_hi_lo_lo_12};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo_lo_1 = {regroupV0_lo_12[2821], regroupV0_lo_12[2817]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo_hi_1 = {regroupV0_lo_12[2829], regroupV0_lo_12[2825]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo_5 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo_hi_1, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi_lo_1 = {regroupV0_lo_12[2837], regroupV0_lo_12[2833]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi_hi_1 = {regroupV0_lo_12[2845], regroupV0_lo_12[2841]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi_5 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi_hi_1, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_9 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi_5, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo_lo_1 = {regroupV0_lo_12[2853], regroupV0_lo_12[2849]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo_hi_1 = {regroupV0_lo_12[2861], regroupV0_lo_12[2857]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo_5 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo_hi_1, regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi_lo_1 = {regroupV0_lo_12[2869], regroupV0_lo_12[2865]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi_hi_1 = {regroupV0_lo_12[2877], regroupV0_lo_12[2873]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi_5 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi_hi_1, regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_9 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi_5, regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_lo_lo_12 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_9, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_9};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo_lo_1 = {regroupV0_lo_12[2885], regroupV0_lo_12[2881]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo_hi_1 = {regroupV0_lo_12[2893], regroupV0_lo_12[2889]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo_5 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo_hi_1, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi_lo_1 = {regroupV0_lo_12[2901], regroupV0_lo_12[2897]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi_hi_1 = {regroupV0_lo_12[2909], regroupV0_lo_12[2905]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi_5 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi_hi_1, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_9 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi_5, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo_lo_1 = {regroupV0_lo_12[2917], regroupV0_lo_12[2913]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo_hi_1 = {regroupV0_lo_12[2925], regroupV0_lo_12[2921]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo_5 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo_hi_1, regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi_lo_1 = {regroupV0_lo_12[2933], regroupV0_lo_12[2929]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi_hi_1 = {regroupV0_lo_12[2941], regroupV0_lo_12[2937]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi_5 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi_hi_1, regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_9 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi_5, regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_lo_hi_12 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_9, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_9};
  wire [31:0]        regroupV0_lo_hi_lo_hi_hi_lo_12 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_12, regroupV0_lo_hi_lo_hi_hi_lo_lo_12};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo_lo_1 = {regroupV0_lo_12[2949], regroupV0_lo_12[2945]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo_hi_1 = {regroupV0_lo_12[2957], regroupV0_lo_12[2953]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo_5 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo_hi_1, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi_lo_1 = {regroupV0_lo_12[2965], regroupV0_lo_12[2961]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi_hi_1 = {regroupV0_lo_12[2973], regroupV0_lo_12[2969]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi_5 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi_hi_1, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_9 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi_5, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo_lo_1 = {regroupV0_lo_12[2981], regroupV0_lo_12[2977]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo_hi_1 = {regroupV0_lo_12[2989], regroupV0_lo_12[2985]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo_5 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo_hi_1, regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi_lo_1 = {regroupV0_lo_12[2997], regroupV0_lo_12[2993]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi_hi_1 = {regroupV0_lo_12[3005], regroupV0_lo_12[3001]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi_5 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi_hi_1, regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_9 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi_5, regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_hi_lo_12 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_9, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_9};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo_lo_1 = {regroupV0_lo_12[3013], regroupV0_lo_12[3009]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo_hi_1 = {regroupV0_lo_12[3021], regroupV0_lo_12[3017]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo_5 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo_hi_1, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi_lo_1 = {regroupV0_lo_12[3029], regroupV0_lo_12[3025]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi_hi_1 = {regroupV0_lo_12[3037], regroupV0_lo_12[3033]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi_5 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi_hi_1, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_9 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi_5, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo_lo_1 = {regroupV0_lo_12[3045], regroupV0_lo_12[3041]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo_hi_1 = {regroupV0_lo_12[3053], regroupV0_lo_12[3049]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo_5 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo_hi_1, regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi_lo_1 = {regroupV0_lo_12[3061], regroupV0_lo_12[3057]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi_hi_1 = {regroupV0_lo_12[3069], regroupV0_lo_12[3065]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi_5 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi_hi_1, regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_9 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi_5, regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_hi_hi_12 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_9, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_9};
  wire [31:0]        regroupV0_lo_hi_lo_hi_hi_hi_12 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_12, regroupV0_lo_hi_lo_hi_hi_hi_lo_12};
  wire [63:0]        regroupV0_lo_hi_lo_hi_hi_12 = {regroupV0_lo_hi_lo_hi_hi_hi_12, regroupV0_lo_hi_lo_hi_hi_lo_12};
  wire [127:0]       regroupV0_lo_hi_lo_hi_12 = {regroupV0_lo_hi_lo_hi_hi_12, regroupV0_lo_hi_lo_hi_lo_12};
  wire [255:0]       regroupV0_lo_hi_lo_12 = {regroupV0_lo_hi_lo_hi_12, regroupV0_lo_hi_lo_lo_12};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo_lo_1 = {regroupV0_lo_12[3077], regroupV0_lo_12[3073]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo_hi_1 = {regroupV0_lo_12[3085], regroupV0_lo_12[3081]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo_5 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo_hi_1, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi_lo_1 = {regroupV0_lo_12[3093], regroupV0_lo_12[3089]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi_hi_1 = {regroupV0_lo_12[3101], regroupV0_lo_12[3097]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi_5 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi_hi_1, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_9 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi_5, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo_lo_1 = {regroupV0_lo_12[3109], regroupV0_lo_12[3105]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo_hi_1 = {regroupV0_lo_12[3117], regroupV0_lo_12[3113]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo_5 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo_hi_1, regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi_lo_1 = {regroupV0_lo_12[3125], regroupV0_lo_12[3121]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi_hi_1 = {regroupV0_lo_12[3133], regroupV0_lo_12[3129]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi_5 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi_hi_1, regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_9 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi_5, regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_lo_lo_12 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_9, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_9};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo_lo_1 = {regroupV0_lo_12[3141], regroupV0_lo_12[3137]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo_hi_1 = {regroupV0_lo_12[3149], regroupV0_lo_12[3145]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo_5 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo_hi_1, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi_lo_1 = {regroupV0_lo_12[3157], regroupV0_lo_12[3153]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi_hi_1 = {regroupV0_lo_12[3165], regroupV0_lo_12[3161]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi_5 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi_hi_1, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_9 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi_5, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo_lo_1 = {regroupV0_lo_12[3173], regroupV0_lo_12[3169]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo_hi_1 = {regroupV0_lo_12[3181], regroupV0_lo_12[3177]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo_5 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo_hi_1, regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi_lo_1 = {regroupV0_lo_12[3189], regroupV0_lo_12[3185]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi_hi_1 = {regroupV0_lo_12[3197], regroupV0_lo_12[3193]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi_5 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi_hi_1, regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_9 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi_5, regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_lo_hi_12 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_9, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_9};
  wire [31:0]        regroupV0_lo_hi_hi_lo_lo_lo_12 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_12, regroupV0_lo_hi_hi_lo_lo_lo_lo_12};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo_lo_1 = {regroupV0_lo_12[3205], regroupV0_lo_12[3201]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo_hi_1 = {regroupV0_lo_12[3213], regroupV0_lo_12[3209]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo_5 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo_hi_1, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi_lo_1 = {regroupV0_lo_12[3221], regroupV0_lo_12[3217]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi_hi_1 = {regroupV0_lo_12[3229], regroupV0_lo_12[3225]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi_5 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi_hi_1, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_9 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi_5, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo_lo_1 = {regroupV0_lo_12[3237], regroupV0_lo_12[3233]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo_hi_1 = {regroupV0_lo_12[3245], regroupV0_lo_12[3241]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo_5 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo_hi_1, regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi_lo_1 = {regroupV0_lo_12[3253], regroupV0_lo_12[3249]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi_hi_1 = {regroupV0_lo_12[3261], regroupV0_lo_12[3257]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi_5 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi_hi_1, regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_9 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi_5, regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_hi_lo_12 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_9, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_9};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo_lo_1 = {regroupV0_lo_12[3269], regroupV0_lo_12[3265]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo_hi_1 = {regroupV0_lo_12[3277], regroupV0_lo_12[3273]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo_5 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo_hi_1, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi_lo_1 = {regroupV0_lo_12[3285], regroupV0_lo_12[3281]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi_hi_1 = {regroupV0_lo_12[3293], regroupV0_lo_12[3289]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi_5 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi_hi_1, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_9 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi_5, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo_lo_1 = {regroupV0_lo_12[3301], regroupV0_lo_12[3297]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo_hi_1 = {regroupV0_lo_12[3309], regroupV0_lo_12[3305]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo_5 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo_hi_1, regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi_lo_1 = {regroupV0_lo_12[3317], regroupV0_lo_12[3313]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi_hi_1 = {regroupV0_lo_12[3325], regroupV0_lo_12[3321]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi_5 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi_hi_1, regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_9 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi_5, regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_hi_hi_12 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_9, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_9};
  wire [31:0]        regroupV0_lo_hi_hi_lo_lo_hi_12 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_12, regroupV0_lo_hi_hi_lo_lo_hi_lo_12};
  wire [63:0]        regroupV0_lo_hi_hi_lo_lo_12 = {regroupV0_lo_hi_hi_lo_lo_hi_12, regroupV0_lo_hi_hi_lo_lo_lo_12};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo_lo_1 = {regroupV0_lo_12[3333], regroupV0_lo_12[3329]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo_hi_1 = {regroupV0_lo_12[3341], regroupV0_lo_12[3337]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo_5 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo_hi_1, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi_lo_1 = {regroupV0_lo_12[3349], regroupV0_lo_12[3345]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi_hi_1 = {regroupV0_lo_12[3357], regroupV0_lo_12[3353]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi_5 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi_hi_1, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_9 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi_5, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo_lo_1 = {regroupV0_lo_12[3365], regroupV0_lo_12[3361]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo_hi_1 = {regroupV0_lo_12[3373], regroupV0_lo_12[3369]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo_5 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo_hi_1, regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi_lo_1 = {regroupV0_lo_12[3381], regroupV0_lo_12[3377]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi_hi_1 = {regroupV0_lo_12[3389], regroupV0_lo_12[3385]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi_5 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi_hi_1, regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_9 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi_5, regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_lo_lo_12 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_9, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_9};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo_lo_1 = {regroupV0_lo_12[3397], regroupV0_lo_12[3393]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo_hi_1 = {regroupV0_lo_12[3405], regroupV0_lo_12[3401]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo_5 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo_hi_1, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi_lo_1 = {regroupV0_lo_12[3413], regroupV0_lo_12[3409]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi_hi_1 = {regroupV0_lo_12[3421], regroupV0_lo_12[3417]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi_5 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi_hi_1, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_9 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi_5, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo_lo_1 = {regroupV0_lo_12[3429], regroupV0_lo_12[3425]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo_hi_1 = {regroupV0_lo_12[3437], regroupV0_lo_12[3433]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo_5 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo_hi_1, regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi_lo_1 = {regroupV0_lo_12[3445], regroupV0_lo_12[3441]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi_hi_1 = {regroupV0_lo_12[3453], regroupV0_lo_12[3449]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi_5 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi_hi_1, regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_9 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi_5, regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_lo_hi_12 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_9, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_9};
  wire [31:0]        regroupV0_lo_hi_hi_lo_hi_lo_12 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_12, regroupV0_lo_hi_hi_lo_hi_lo_lo_12};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo_lo_1 = {regroupV0_lo_12[3461], regroupV0_lo_12[3457]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo_hi_1 = {regroupV0_lo_12[3469], regroupV0_lo_12[3465]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo_5 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo_hi_1, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi_lo_1 = {regroupV0_lo_12[3477], regroupV0_lo_12[3473]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi_hi_1 = {regroupV0_lo_12[3485], regroupV0_lo_12[3481]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi_5 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi_hi_1, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_9 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi_5, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo_lo_1 = {regroupV0_lo_12[3493], regroupV0_lo_12[3489]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo_hi_1 = {regroupV0_lo_12[3501], regroupV0_lo_12[3497]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo_5 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo_hi_1, regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi_lo_1 = {regroupV0_lo_12[3509], regroupV0_lo_12[3505]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi_hi_1 = {regroupV0_lo_12[3517], regroupV0_lo_12[3513]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi_5 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi_hi_1, regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_9 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi_5, regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_hi_lo_12 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_9, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_9};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo_lo_1 = {regroupV0_lo_12[3525], regroupV0_lo_12[3521]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo_hi_1 = {regroupV0_lo_12[3533], regroupV0_lo_12[3529]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo_5 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo_hi_1, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi_lo_1 = {regroupV0_lo_12[3541], regroupV0_lo_12[3537]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi_hi_1 = {regroupV0_lo_12[3549], regroupV0_lo_12[3545]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi_5 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi_hi_1, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_9 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi_5, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo_lo_1 = {regroupV0_lo_12[3557], regroupV0_lo_12[3553]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo_hi_1 = {regroupV0_lo_12[3565], regroupV0_lo_12[3561]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo_5 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo_hi_1, regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi_lo_1 = {regroupV0_lo_12[3573], regroupV0_lo_12[3569]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi_hi_1 = {regroupV0_lo_12[3581], regroupV0_lo_12[3577]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi_5 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi_hi_1, regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_9 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi_5, regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_hi_hi_12 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_9, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_9};
  wire [31:0]        regroupV0_lo_hi_hi_lo_hi_hi_12 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_12, regroupV0_lo_hi_hi_lo_hi_hi_lo_12};
  wire [63:0]        regroupV0_lo_hi_hi_lo_hi_12 = {regroupV0_lo_hi_hi_lo_hi_hi_12, regroupV0_lo_hi_hi_lo_hi_lo_12};
  wire [127:0]       regroupV0_lo_hi_hi_lo_12 = {regroupV0_lo_hi_hi_lo_hi_12, regroupV0_lo_hi_hi_lo_lo_12};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo_lo_1 = {regroupV0_lo_12[3589], regroupV0_lo_12[3585]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo_hi_1 = {regroupV0_lo_12[3597], regroupV0_lo_12[3593]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo_5 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo_hi_1, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi_lo_1 = {regroupV0_lo_12[3605], regroupV0_lo_12[3601]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi_hi_1 = {regroupV0_lo_12[3613], regroupV0_lo_12[3609]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi_5 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi_hi_1, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_9 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi_5, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo_lo_1 = {regroupV0_lo_12[3621], regroupV0_lo_12[3617]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo_hi_1 = {regroupV0_lo_12[3629], regroupV0_lo_12[3625]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo_5 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo_hi_1, regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi_lo_1 = {regroupV0_lo_12[3637], regroupV0_lo_12[3633]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi_hi_1 = {regroupV0_lo_12[3645], regroupV0_lo_12[3641]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi_5 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi_hi_1, regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_9 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi_5, regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_lo_lo_12 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_9, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_9};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo_lo_1 = {regroupV0_lo_12[3653], regroupV0_lo_12[3649]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo_hi_1 = {regroupV0_lo_12[3661], regroupV0_lo_12[3657]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo_5 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo_hi_1, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi_lo_1 = {regroupV0_lo_12[3669], regroupV0_lo_12[3665]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi_hi_1 = {regroupV0_lo_12[3677], regroupV0_lo_12[3673]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi_5 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi_hi_1, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_9 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi_5, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo_lo_1 = {regroupV0_lo_12[3685], regroupV0_lo_12[3681]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo_hi_1 = {regroupV0_lo_12[3693], regroupV0_lo_12[3689]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo_5 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo_hi_1, regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi_lo_1 = {regroupV0_lo_12[3701], regroupV0_lo_12[3697]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi_hi_1 = {regroupV0_lo_12[3709], regroupV0_lo_12[3705]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi_5 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi_hi_1, regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_9 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi_5, regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_lo_hi_12 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_9, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_9};
  wire [31:0]        regroupV0_lo_hi_hi_hi_lo_lo_12 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_12, regroupV0_lo_hi_hi_hi_lo_lo_lo_12};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo_lo_1 = {regroupV0_lo_12[3717], regroupV0_lo_12[3713]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo_hi_1 = {regroupV0_lo_12[3725], regroupV0_lo_12[3721]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo_5 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo_hi_1, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi_lo_1 = {regroupV0_lo_12[3733], regroupV0_lo_12[3729]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi_hi_1 = {regroupV0_lo_12[3741], regroupV0_lo_12[3737]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi_5 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi_hi_1, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_9 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi_5, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo_lo_1 = {regroupV0_lo_12[3749], regroupV0_lo_12[3745]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo_hi_1 = {regroupV0_lo_12[3757], regroupV0_lo_12[3753]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo_5 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo_hi_1, regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi_lo_1 = {regroupV0_lo_12[3765], regroupV0_lo_12[3761]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi_hi_1 = {regroupV0_lo_12[3773], regroupV0_lo_12[3769]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi_5 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi_hi_1, regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_9 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi_5, regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_hi_lo_12 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_9, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_9};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo_lo_1 = {regroupV0_lo_12[3781], regroupV0_lo_12[3777]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo_hi_1 = {regroupV0_lo_12[3789], regroupV0_lo_12[3785]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo_5 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo_hi_1, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi_lo_1 = {regroupV0_lo_12[3797], regroupV0_lo_12[3793]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi_hi_1 = {regroupV0_lo_12[3805], regroupV0_lo_12[3801]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi_5 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi_hi_1, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_9 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi_5, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo_lo_1 = {regroupV0_lo_12[3813], regroupV0_lo_12[3809]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo_hi_1 = {regroupV0_lo_12[3821], regroupV0_lo_12[3817]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo_5 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo_hi_1, regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi_lo_1 = {regroupV0_lo_12[3829], regroupV0_lo_12[3825]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi_hi_1 = {regroupV0_lo_12[3837], regroupV0_lo_12[3833]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi_5 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi_hi_1, regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_9 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi_5, regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_hi_hi_12 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_9, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_9};
  wire [31:0]        regroupV0_lo_hi_hi_hi_lo_hi_12 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_12, regroupV0_lo_hi_hi_hi_lo_hi_lo_12};
  wire [63:0]        regroupV0_lo_hi_hi_hi_lo_12 = {regroupV0_lo_hi_hi_hi_lo_hi_12, regroupV0_lo_hi_hi_hi_lo_lo_12};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo_lo_1 = {regroupV0_lo_12[3845], regroupV0_lo_12[3841]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo_hi_1 = {regroupV0_lo_12[3853], regroupV0_lo_12[3849]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo_5 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo_hi_1, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi_lo_1 = {regroupV0_lo_12[3861], regroupV0_lo_12[3857]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi_hi_1 = {regroupV0_lo_12[3869], regroupV0_lo_12[3865]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi_5 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi_hi_1, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_9 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi_5, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo_lo_1 = {regroupV0_lo_12[3877], regroupV0_lo_12[3873]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo_hi_1 = {regroupV0_lo_12[3885], regroupV0_lo_12[3881]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo_5 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo_hi_1, regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi_lo_1 = {regroupV0_lo_12[3893], regroupV0_lo_12[3889]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi_hi_1 = {regroupV0_lo_12[3901], regroupV0_lo_12[3897]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi_5 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi_hi_1, regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_9 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi_5, regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_lo_lo_12 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_9, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_9};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo_lo_1 = {regroupV0_lo_12[3909], regroupV0_lo_12[3905]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo_hi_1 = {regroupV0_lo_12[3917], regroupV0_lo_12[3913]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo_5 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo_hi_1, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi_lo_1 = {regroupV0_lo_12[3925], regroupV0_lo_12[3921]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi_hi_1 = {regroupV0_lo_12[3933], regroupV0_lo_12[3929]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi_5 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi_hi_1, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_9 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi_5, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo_lo_1 = {regroupV0_lo_12[3941], regroupV0_lo_12[3937]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo_hi_1 = {regroupV0_lo_12[3949], regroupV0_lo_12[3945]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo_5 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo_hi_1, regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi_lo_1 = {regroupV0_lo_12[3957], regroupV0_lo_12[3953]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi_hi_1 = {regroupV0_lo_12[3965], regroupV0_lo_12[3961]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi_5 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi_hi_1, regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_9 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi_5, regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_lo_hi_12 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_9, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_9};
  wire [31:0]        regroupV0_lo_hi_hi_hi_hi_lo_12 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_12, regroupV0_lo_hi_hi_hi_hi_lo_lo_12};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo_lo_1 = {regroupV0_lo_12[3973], regroupV0_lo_12[3969]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo_hi_1 = {regroupV0_lo_12[3981], regroupV0_lo_12[3977]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo_5 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo_hi_1, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi_lo_1 = {regroupV0_lo_12[3989], regroupV0_lo_12[3985]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi_hi_1 = {regroupV0_lo_12[3997], regroupV0_lo_12[3993]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi_5 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi_hi_1, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_9 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi_5, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo_lo_1 = {regroupV0_lo_12[4005], regroupV0_lo_12[4001]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo_hi_1 = {regroupV0_lo_12[4013], regroupV0_lo_12[4009]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo_5 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo_hi_1, regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi_lo_1 = {regroupV0_lo_12[4021], regroupV0_lo_12[4017]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi_hi_1 = {regroupV0_lo_12[4029], regroupV0_lo_12[4025]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi_5 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi_hi_1, regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_9 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi_5, regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_hi_lo_12 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_9, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_9};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo_lo_1 = {regroupV0_lo_12[4037], regroupV0_lo_12[4033]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo_hi_1 = {regroupV0_lo_12[4045], regroupV0_lo_12[4041]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo_5 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo_hi_1, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi_lo_1 = {regroupV0_lo_12[4053], regroupV0_lo_12[4049]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi_hi_1 = {regroupV0_lo_12[4061], regroupV0_lo_12[4057]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi_5 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi_hi_1, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_9 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi_5, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo_lo_1 = {regroupV0_lo_12[4069], regroupV0_lo_12[4065]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo_hi_1 = {regroupV0_lo_12[4077], regroupV0_lo_12[4073]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo_5 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo_hi_1, regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi_lo_1 = {regroupV0_lo_12[4085], regroupV0_lo_12[4081]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi_hi_1 = {regroupV0_lo_12[4093], regroupV0_lo_12[4089]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi_5 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi_hi_1, regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_9 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi_5, regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_hi_hi_12 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_9, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_9};
  wire [31:0]        regroupV0_lo_hi_hi_hi_hi_hi_12 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_12, regroupV0_lo_hi_hi_hi_hi_hi_lo_12};
  wire [63:0]        regroupV0_lo_hi_hi_hi_hi_12 = {regroupV0_lo_hi_hi_hi_hi_hi_12, regroupV0_lo_hi_hi_hi_hi_lo_12};
  wire [127:0]       regroupV0_lo_hi_hi_hi_12 = {regroupV0_lo_hi_hi_hi_hi_12, regroupV0_lo_hi_hi_hi_lo_12};
  wire [255:0]       regroupV0_lo_hi_hi_12 = {regroupV0_lo_hi_hi_hi_12, regroupV0_lo_hi_hi_lo_12};
  wire [511:0]       regroupV0_lo_hi_12 = {regroupV0_lo_hi_hi_12, regroupV0_lo_hi_lo_12};
  wire [1023:0]      regroupV0_lo_14 = {regroupV0_lo_hi_12, regroupV0_lo_lo_12};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo_lo_1 = {regroupV0_hi_12[5], regroupV0_hi_12[1]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo_hi_1 = {regroupV0_hi_12[13], regroupV0_hi_12[9]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo_5 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi_lo_1 = {regroupV0_hi_12[21], regroupV0_hi_12[17]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi_hi_1 = {regroupV0_hi_12[29], regroupV0_hi_12[25]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi_5 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi_hi_1, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_9 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi_5, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo_lo_1 = {regroupV0_hi_12[37], regroupV0_hi_12[33]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo_hi_1 = {regroupV0_hi_12[45], regroupV0_hi_12[41]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo_5 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo_hi_1, regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi_lo_1 = {regroupV0_hi_12[53], regroupV0_hi_12[49]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi_hi_1 = {regroupV0_hi_12[61], regroupV0_hi_12[57]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi_5 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi_hi_1, regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_9 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi_5, regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_lo_lo_12 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_9, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_9};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo_lo_1 = {regroupV0_hi_12[69], regroupV0_hi_12[65]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo_hi_1 = {regroupV0_hi_12[77], regroupV0_hi_12[73]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo_5 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi_lo_1 = {regroupV0_hi_12[85], regroupV0_hi_12[81]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi_hi_1 = {regroupV0_hi_12[93], regroupV0_hi_12[89]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi_5 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi_hi_1, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_9 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi_5, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo_lo_1 = {regroupV0_hi_12[101], regroupV0_hi_12[97]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo_hi_1 = {regroupV0_hi_12[109], regroupV0_hi_12[105]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo_5 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo_hi_1, regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi_lo_1 = {regroupV0_hi_12[117], regroupV0_hi_12[113]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi_hi_1 = {regroupV0_hi_12[125], regroupV0_hi_12[121]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi_5 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi_hi_1, regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_9 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi_5, regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_lo_hi_12 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_9, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_9};
  wire [31:0]        regroupV0_hi_lo_lo_lo_lo_lo_12 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_12, regroupV0_hi_lo_lo_lo_lo_lo_lo_12};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo_lo_1 = {regroupV0_hi_12[133], regroupV0_hi_12[129]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo_hi_1 = {regroupV0_hi_12[141], regroupV0_hi_12[137]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo_5 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi_lo_1 = {regroupV0_hi_12[149], regroupV0_hi_12[145]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi_hi_1 = {regroupV0_hi_12[157], regroupV0_hi_12[153]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi_5 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi_hi_1, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_9 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi_5, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo_lo_1 = {regroupV0_hi_12[165], regroupV0_hi_12[161]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo_hi_1 = {regroupV0_hi_12[173], regroupV0_hi_12[169]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo_5 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo_hi_1, regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi_lo_1 = {regroupV0_hi_12[181], regroupV0_hi_12[177]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi_hi_1 = {regroupV0_hi_12[189], regroupV0_hi_12[185]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi_5 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi_hi_1, regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_9 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi_5, regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_hi_lo_12 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_9, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_9};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo_lo_1 = {regroupV0_hi_12[197], regroupV0_hi_12[193]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo_hi_1 = {regroupV0_hi_12[205], regroupV0_hi_12[201]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo_5 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi_lo_1 = {regroupV0_hi_12[213], regroupV0_hi_12[209]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi_hi_1 = {regroupV0_hi_12[221], regroupV0_hi_12[217]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi_5 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi_hi_1, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_9 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi_5, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo_lo_1 = {regroupV0_hi_12[229], regroupV0_hi_12[225]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo_hi_1 = {regroupV0_hi_12[237], regroupV0_hi_12[233]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo_5 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo_hi_1, regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi_lo_1 = {regroupV0_hi_12[245], regroupV0_hi_12[241]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi_hi_1 = {regroupV0_hi_12[253], regroupV0_hi_12[249]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi_5 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi_hi_1, regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_9 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi_5, regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_hi_hi_12 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_9, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_9};
  wire [31:0]        regroupV0_hi_lo_lo_lo_lo_hi_12 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_12, regroupV0_hi_lo_lo_lo_lo_hi_lo_12};
  wire [63:0]        regroupV0_hi_lo_lo_lo_lo_12 = {regroupV0_hi_lo_lo_lo_lo_hi_12, regroupV0_hi_lo_lo_lo_lo_lo_12};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo_lo_1 = {regroupV0_hi_12[261], regroupV0_hi_12[257]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo_hi_1 = {regroupV0_hi_12[269], regroupV0_hi_12[265]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo_5 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi_lo_1 = {regroupV0_hi_12[277], regroupV0_hi_12[273]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi_hi_1 = {regroupV0_hi_12[285], regroupV0_hi_12[281]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi_5 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi_hi_1, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_9 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi_5, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo_lo_1 = {regroupV0_hi_12[293], regroupV0_hi_12[289]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo_hi_1 = {regroupV0_hi_12[301], regroupV0_hi_12[297]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo_5 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo_hi_1, regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi_lo_1 = {regroupV0_hi_12[309], regroupV0_hi_12[305]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi_hi_1 = {regroupV0_hi_12[317], regroupV0_hi_12[313]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi_5 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi_hi_1, regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_9 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi_5, regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_lo_lo_12 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_9, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_9};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo_lo_1 = {regroupV0_hi_12[325], regroupV0_hi_12[321]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo_hi_1 = {regroupV0_hi_12[333], regroupV0_hi_12[329]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo_5 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi_lo_1 = {regroupV0_hi_12[341], regroupV0_hi_12[337]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi_hi_1 = {regroupV0_hi_12[349], regroupV0_hi_12[345]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi_5 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi_hi_1, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_9 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi_5, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo_lo_1 = {regroupV0_hi_12[357], regroupV0_hi_12[353]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo_hi_1 = {regroupV0_hi_12[365], regroupV0_hi_12[361]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo_5 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo_hi_1, regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi_lo_1 = {regroupV0_hi_12[373], regroupV0_hi_12[369]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi_hi_1 = {regroupV0_hi_12[381], regroupV0_hi_12[377]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi_5 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi_hi_1, regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_9 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi_5, regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_lo_hi_12 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_9, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_9};
  wire [31:0]        regroupV0_hi_lo_lo_lo_hi_lo_12 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_12, regroupV0_hi_lo_lo_lo_hi_lo_lo_12};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo_lo_1 = {regroupV0_hi_12[389], regroupV0_hi_12[385]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo_hi_1 = {regroupV0_hi_12[397], regroupV0_hi_12[393]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo_5 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi_lo_1 = {regroupV0_hi_12[405], regroupV0_hi_12[401]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi_hi_1 = {regroupV0_hi_12[413], regroupV0_hi_12[409]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi_5 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi_hi_1, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_9 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi_5, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo_lo_1 = {regroupV0_hi_12[421], regroupV0_hi_12[417]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo_hi_1 = {regroupV0_hi_12[429], regroupV0_hi_12[425]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo_5 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo_hi_1, regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi_lo_1 = {regroupV0_hi_12[437], regroupV0_hi_12[433]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi_hi_1 = {regroupV0_hi_12[445], regroupV0_hi_12[441]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi_5 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi_hi_1, regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_9 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi_5, regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_hi_lo_12 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_9, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_9};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo_lo_1 = {regroupV0_hi_12[453], regroupV0_hi_12[449]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo_hi_1 = {regroupV0_hi_12[461], regroupV0_hi_12[457]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo_5 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi_lo_1 = {regroupV0_hi_12[469], regroupV0_hi_12[465]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi_hi_1 = {regroupV0_hi_12[477], regroupV0_hi_12[473]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi_5 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi_hi_1, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_9 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi_5, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo_lo_1 = {regroupV0_hi_12[485], regroupV0_hi_12[481]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo_hi_1 = {regroupV0_hi_12[493], regroupV0_hi_12[489]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo_5 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo_hi_1, regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi_lo_1 = {regroupV0_hi_12[501], regroupV0_hi_12[497]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi_hi_1 = {regroupV0_hi_12[509], regroupV0_hi_12[505]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi_5 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi_hi_1, regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_9 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi_5, regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_hi_hi_12 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_9, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_9};
  wire [31:0]        regroupV0_hi_lo_lo_lo_hi_hi_12 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_12, regroupV0_hi_lo_lo_lo_hi_hi_lo_12};
  wire [63:0]        regroupV0_hi_lo_lo_lo_hi_12 = {regroupV0_hi_lo_lo_lo_hi_hi_12, regroupV0_hi_lo_lo_lo_hi_lo_12};
  wire [127:0]       regroupV0_hi_lo_lo_lo_12 = {regroupV0_hi_lo_lo_lo_hi_12, regroupV0_hi_lo_lo_lo_lo_12};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo_lo_1 = {regroupV0_hi_12[517], regroupV0_hi_12[513]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo_hi_1 = {regroupV0_hi_12[525], regroupV0_hi_12[521]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo_5 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo_hi_1, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi_lo_1 = {regroupV0_hi_12[533], regroupV0_hi_12[529]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi_hi_1 = {regroupV0_hi_12[541], regroupV0_hi_12[537]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi_5 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi_hi_1, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_9 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi_5, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo_lo_1 = {regroupV0_hi_12[549], regroupV0_hi_12[545]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo_hi_1 = {regroupV0_hi_12[557], regroupV0_hi_12[553]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo_5 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo_hi_1, regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi_lo_1 = {regroupV0_hi_12[565], regroupV0_hi_12[561]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi_hi_1 = {regroupV0_hi_12[573], regroupV0_hi_12[569]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi_5 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi_hi_1, regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_9 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi_5, regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_lo_lo_12 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_9, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_9};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo_lo_1 = {regroupV0_hi_12[581], regroupV0_hi_12[577]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo_hi_1 = {regroupV0_hi_12[589], regroupV0_hi_12[585]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo_5 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo_hi_1, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi_lo_1 = {regroupV0_hi_12[597], regroupV0_hi_12[593]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi_hi_1 = {regroupV0_hi_12[605], regroupV0_hi_12[601]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi_5 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi_hi_1, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_9 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi_5, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo_lo_1 = {regroupV0_hi_12[613], regroupV0_hi_12[609]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo_hi_1 = {regroupV0_hi_12[621], regroupV0_hi_12[617]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo_5 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo_hi_1, regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi_lo_1 = {regroupV0_hi_12[629], regroupV0_hi_12[625]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi_hi_1 = {regroupV0_hi_12[637], regroupV0_hi_12[633]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi_5 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi_hi_1, regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_9 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi_5, regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_lo_hi_12 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_9, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_9};
  wire [31:0]        regroupV0_hi_lo_lo_hi_lo_lo_12 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_12, regroupV0_hi_lo_lo_hi_lo_lo_lo_12};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo_lo_1 = {regroupV0_hi_12[645], regroupV0_hi_12[641]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo_hi_1 = {regroupV0_hi_12[653], regroupV0_hi_12[649]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo_5 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo_hi_1, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi_lo_1 = {regroupV0_hi_12[661], regroupV0_hi_12[657]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi_hi_1 = {regroupV0_hi_12[669], regroupV0_hi_12[665]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi_5 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi_hi_1, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_9 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi_5, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo_lo_1 = {regroupV0_hi_12[677], regroupV0_hi_12[673]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo_hi_1 = {regroupV0_hi_12[685], regroupV0_hi_12[681]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo_5 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo_hi_1, regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi_lo_1 = {regroupV0_hi_12[693], regroupV0_hi_12[689]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi_hi_1 = {regroupV0_hi_12[701], regroupV0_hi_12[697]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi_5 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi_hi_1, regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_9 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi_5, regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_hi_lo_12 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_9, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_9};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo_lo_1 = {regroupV0_hi_12[709], regroupV0_hi_12[705]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo_hi_1 = {regroupV0_hi_12[717], regroupV0_hi_12[713]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo_5 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo_hi_1, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi_lo_1 = {regroupV0_hi_12[725], regroupV0_hi_12[721]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi_hi_1 = {regroupV0_hi_12[733], regroupV0_hi_12[729]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi_5 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi_hi_1, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_9 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi_5, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo_lo_1 = {regroupV0_hi_12[741], regroupV0_hi_12[737]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo_hi_1 = {regroupV0_hi_12[749], regroupV0_hi_12[745]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo_5 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo_hi_1, regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi_lo_1 = {regroupV0_hi_12[757], regroupV0_hi_12[753]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi_hi_1 = {regroupV0_hi_12[765], regroupV0_hi_12[761]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi_5 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi_hi_1, regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_9 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi_5, regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_hi_hi_12 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_9, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_9};
  wire [31:0]        regroupV0_hi_lo_lo_hi_lo_hi_12 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_12, regroupV0_hi_lo_lo_hi_lo_hi_lo_12};
  wire [63:0]        regroupV0_hi_lo_lo_hi_lo_12 = {regroupV0_hi_lo_lo_hi_lo_hi_12, regroupV0_hi_lo_lo_hi_lo_lo_12};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo_lo_1 = {regroupV0_hi_12[773], regroupV0_hi_12[769]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo_hi_1 = {regroupV0_hi_12[781], regroupV0_hi_12[777]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo_5 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo_hi_1, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi_lo_1 = {regroupV0_hi_12[789], regroupV0_hi_12[785]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi_hi_1 = {regroupV0_hi_12[797], regroupV0_hi_12[793]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi_5 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi_hi_1, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_9 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi_5, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo_lo_1 = {regroupV0_hi_12[805], regroupV0_hi_12[801]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo_hi_1 = {regroupV0_hi_12[813], regroupV0_hi_12[809]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo_5 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo_hi_1, regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi_lo_1 = {regroupV0_hi_12[821], regroupV0_hi_12[817]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi_hi_1 = {regroupV0_hi_12[829], regroupV0_hi_12[825]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi_5 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi_hi_1, regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_9 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi_5, regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_lo_lo_12 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_9, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_9};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo_lo_1 = {regroupV0_hi_12[837], regroupV0_hi_12[833]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo_hi_1 = {regroupV0_hi_12[845], regroupV0_hi_12[841]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo_5 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo_hi_1, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi_lo_1 = {regroupV0_hi_12[853], regroupV0_hi_12[849]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi_hi_1 = {regroupV0_hi_12[861], regroupV0_hi_12[857]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi_5 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi_hi_1, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_9 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi_5, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo_lo_1 = {regroupV0_hi_12[869], regroupV0_hi_12[865]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo_hi_1 = {regroupV0_hi_12[877], regroupV0_hi_12[873]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo_5 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo_hi_1, regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi_lo_1 = {regroupV0_hi_12[885], regroupV0_hi_12[881]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi_hi_1 = {regroupV0_hi_12[893], regroupV0_hi_12[889]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi_5 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi_hi_1, regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_9 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi_5, regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_lo_hi_12 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_9, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_9};
  wire [31:0]        regroupV0_hi_lo_lo_hi_hi_lo_12 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_12, regroupV0_hi_lo_lo_hi_hi_lo_lo_12};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo_lo_1 = {regroupV0_hi_12[901], regroupV0_hi_12[897]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo_hi_1 = {regroupV0_hi_12[909], regroupV0_hi_12[905]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo_5 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo_hi_1, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi_lo_1 = {regroupV0_hi_12[917], regroupV0_hi_12[913]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi_hi_1 = {regroupV0_hi_12[925], regroupV0_hi_12[921]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi_5 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi_hi_1, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_9 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi_5, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo_lo_1 = {regroupV0_hi_12[933], regroupV0_hi_12[929]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo_hi_1 = {regroupV0_hi_12[941], regroupV0_hi_12[937]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo_5 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo_hi_1, regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi_lo_1 = {regroupV0_hi_12[949], regroupV0_hi_12[945]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi_hi_1 = {regroupV0_hi_12[957], regroupV0_hi_12[953]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi_5 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi_hi_1, regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_9 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi_5, regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_hi_lo_12 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_9, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_9};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo_lo_1 = {regroupV0_hi_12[965], regroupV0_hi_12[961]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo_hi_1 = {regroupV0_hi_12[973], regroupV0_hi_12[969]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo_5 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo_hi_1, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi_lo_1 = {regroupV0_hi_12[981], regroupV0_hi_12[977]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi_hi_1 = {regroupV0_hi_12[989], regroupV0_hi_12[985]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi_5 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi_hi_1, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_9 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi_5, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo_lo_1 = {regroupV0_hi_12[997], regroupV0_hi_12[993]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo_hi_1 = {regroupV0_hi_12[1005], regroupV0_hi_12[1001]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo_5 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo_hi_1, regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi_lo_1 = {regroupV0_hi_12[1013], regroupV0_hi_12[1009]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi_hi_1 = {regroupV0_hi_12[1021], regroupV0_hi_12[1017]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi_5 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi_hi_1, regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_9 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi_5, regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_hi_hi_12 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_9, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_9};
  wire [31:0]        regroupV0_hi_lo_lo_hi_hi_hi_12 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_12, regroupV0_hi_lo_lo_hi_hi_hi_lo_12};
  wire [63:0]        regroupV0_hi_lo_lo_hi_hi_12 = {regroupV0_hi_lo_lo_hi_hi_hi_12, regroupV0_hi_lo_lo_hi_hi_lo_12};
  wire [127:0]       regroupV0_hi_lo_lo_hi_12 = {regroupV0_hi_lo_lo_hi_hi_12, regroupV0_hi_lo_lo_hi_lo_12};
  wire [255:0]       regroupV0_hi_lo_lo_12 = {regroupV0_hi_lo_lo_hi_12, regroupV0_hi_lo_lo_lo_12};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo_lo_1 = {regroupV0_hi_12[1029], regroupV0_hi_12[1025]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo_hi_1 = {regroupV0_hi_12[1037], regroupV0_hi_12[1033]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo_5 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo_hi_1, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi_lo_1 = {regroupV0_hi_12[1045], regroupV0_hi_12[1041]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi_hi_1 = {regroupV0_hi_12[1053], regroupV0_hi_12[1049]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi_5 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi_hi_1, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_9 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi_5, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo_lo_1 = {regroupV0_hi_12[1061], regroupV0_hi_12[1057]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo_hi_1 = {regroupV0_hi_12[1069], regroupV0_hi_12[1065]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo_5 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo_hi_1, regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi_lo_1 = {regroupV0_hi_12[1077], regroupV0_hi_12[1073]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi_hi_1 = {regroupV0_hi_12[1085], regroupV0_hi_12[1081]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi_5 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi_hi_1, regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_9 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi_5, regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_lo_lo_12 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_9, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_9};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo_lo_1 = {regroupV0_hi_12[1093], regroupV0_hi_12[1089]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo_hi_1 = {regroupV0_hi_12[1101], regroupV0_hi_12[1097]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo_5 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo_hi_1, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi_lo_1 = {regroupV0_hi_12[1109], regroupV0_hi_12[1105]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi_hi_1 = {regroupV0_hi_12[1117], regroupV0_hi_12[1113]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi_5 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi_hi_1, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_9 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi_5, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo_lo_1 = {regroupV0_hi_12[1125], regroupV0_hi_12[1121]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo_hi_1 = {regroupV0_hi_12[1133], regroupV0_hi_12[1129]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo_5 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo_hi_1, regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi_lo_1 = {regroupV0_hi_12[1141], regroupV0_hi_12[1137]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi_hi_1 = {regroupV0_hi_12[1149], regroupV0_hi_12[1145]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi_5 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi_hi_1, regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_9 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi_5, regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_lo_hi_12 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_9, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_9};
  wire [31:0]        regroupV0_hi_lo_hi_lo_lo_lo_12 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_12, regroupV0_hi_lo_hi_lo_lo_lo_lo_12};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo_lo_1 = {regroupV0_hi_12[1157], regroupV0_hi_12[1153]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo_hi_1 = {regroupV0_hi_12[1165], regroupV0_hi_12[1161]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo_5 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo_hi_1, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi_lo_1 = {regroupV0_hi_12[1173], regroupV0_hi_12[1169]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi_hi_1 = {regroupV0_hi_12[1181], regroupV0_hi_12[1177]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi_5 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi_hi_1, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_9 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi_5, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo_lo_1 = {regroupV0_hi_12[1189], regroupV0_hi_12[1185]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo_hi_1 = {regroupV0_hi_12[1197], regroupV0_hi_12[1193]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo_5 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo_hi_1, regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi_lo_1 = {regroupV0_hi_12[1205], regroupV0_hi_12[1201]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi_hi_1 = {regroupV0_hi_12[1213], regroupV0_hi_12[1209]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi_5 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi_hi_1, regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_9 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi_5, regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_hi_lo_12 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_9, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_9};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo_lo_1 = {regroupV0_hi_12[1221], regroupV0_hi_12[1217]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo_hi_1 = {regroupV0_hi_12[1229], regroupV0_hi_12[1225]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo_5 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo_hi_1, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi_lo_1 = {regroupV0_hi_12[1237], regroupV0_hi_12[1233]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi_hi_1 = {regroupV0_hi_12[1245], regroupV0_hi_12[1241]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi_5 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi_hi_1, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_9 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi_5, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo_lo_1 = {regroupV0_hi_12[1253], regroupV0_hi_12[1249]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo_hi_1 = {regroupV0_hi_12[1261], regroupV0_hi_12[1257]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo_5 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo_hi_1, regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi_lo_1 = {regroupV0_hi_12[1269], regroupV0_hi_12[1265]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi_hi_1 = {regroupV0_hi_12[1277], regroupV0_hi_12[1273]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi_5 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi_hi_1, regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_9 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi_5, regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_hi_hi_12 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_9, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_9};
  wire [31:0]        regroupV0_hi_lo_hi_lo_lo_hi_12 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_12, regroupV0_hi_lo_hi_lo_lo_hi_lo_12};
  wire [63:0]        regroupV0_hi_lo_hi_lo_lo_12 = {regroupV0_hi_lo_hi_lo_lo_hi_12, regroupV0_hi_lo_hi_lo_lo_lo_12};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo_lo_1 = {regroupV0_hi_12[1285], regroupV0_hi_12[1281]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo_hi_1 = {regroupV0_hi_12[1293], regroupV0_hi_12[1289]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo_5 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo_hi_1, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi_lo_1 = {regroupV0_hi_12[1301], regroupV0_hi_12[1297]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi_hi_1 = {regroupV0_hi_12[1309], regroupV0_hi_12[1305]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi_5 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi_hi_1, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_9 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi_5, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo_lo_1 = {regroupV0_hi_12[1317], regroupV0_hi_12[1313]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo_hi_1 = {regroupV0_hi_12[1325], regroupV0_hi_12[1321]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo_5 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo_hi_1, regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi_lo_1 = {regroupV0_hi_12[1333], regroupV0_hi_12[1329]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi_hi_1 = {regroupV0_hi_12[1341], regroupV0_hi_12[1337]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi_5 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi_hi_1, regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_9 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi_5, regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_lo_lo_12 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_9, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_9};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo_lo_1 = {regroupV0_hi_12[1349], regroupV0_hi_12[1345]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo_hi_1 = {regroupV0_hi_12[1357], regroupV0_hi_12[1353]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo_5 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo_hi_1, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi_lo_1 = {regroupV0_hi_12[1365], regroupV0_hi_12[1361]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi_hi_1 = {regroupV0_hi_12[1373], regroupV0_hi_12[1369]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi_5 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi_hi_1, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_9 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi_5, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo_lo_1 = {regroupV0_hi_12[1381], regroupV0_hi_12[1377]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo_hi_1 = {regroupV0_hi_12[1389], regroupV0_hi_12[1385]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo_5 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo_hi_1, regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi_lo_1 = {regroupV0_hi_12[1397], regroupV0_hi_12[1393]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi_hi_1 = {regroupV0_hi_12[1405], regroupV0_hi_12[1401]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi_5 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi_hi_1, regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_9 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi_5, regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_lo_hi_12 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_9, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_9};
  wire [31:0]        regroupV0_hi_lo_hi_lo_hi_lo_12 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_12, regroupV0_hi_lo_hi_lo_hi_lo_lo_12};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo_lo_1 = {regroupV0_hi_12[1413], regroupV0_hi_12[1409]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo_hi_1 = {regroupV0_hi_12[1421], regroupV0_hi_12[1417]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo_5 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo_hi_1, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi_lo_1 = {regroupV0_hi_12[1429], regroupV0_hi_12[1425]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi_hi_1 = {regroupV0_hi_12[1437], regroupV0_hi_12[1433]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi_5 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi_hi_1, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_9 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi_5, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo_lo_1 = {regroupV0_hi_12[1445], regroupV0_hi_12[1441]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo_hi_1 = {regroupV0_hi_12[1453], regroupV0_hi_12[1449]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo_5 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo_hi_1, regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi_lo_1 = {regroupV0_hi_12[1461], regroupV0_hi_12[1457]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi_hi_1 = {regroupV0_hi_12[1469], regroupV0_hi_12[1465]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi_5 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi_hi_1, regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_9 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi_5, regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_hi_lo_12 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_9, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_9};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo_lo_1 = {regroupV0_hi_12[1477], regroupV0_hi_12[1473]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo_hi_1 = {regroupV0_hi_12[1485], regroupV0_hi_12[1481]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo_5 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo_hi_1, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi_lo_1 = {regroupV0_hi_12[1493], regroupV0_hi_12[1489]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi_hi_1 = {regroupV0_hi_12[1501], regroupV0_hi_12[1497]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi_5 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi_hi_1, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_9 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi_5, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo_lo_1 = {regroupV0_hi_12[1509], regroupV0_hi_12[1505]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo_hi_1 = {regroupV0_hi_12[1517], regroupV0_hi_12[1513]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo_5 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo_hi_1, regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi_lo_1 = {regroupV0_hi_12[1525], regroupV0_hi_12[1521]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi_hi_1 = {regroupV0_hi_12[1533], regroupV0_hi_12[1529]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi_5 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi_hi_1, regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_9 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi_5, regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_hi_hi_12 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_9, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_9};
  wire [31:0]        regroupV0_hi_lo_hi_lo_hi_hi_12 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_12, regroupV0_hi_lo_hi_lo_hi_hi_lo_12};
  wire [63:0]        regroupV0_hi_lo_hi_lo_hi_12 = {regroupV0_hi_lo_hi_lo_hi_hi_12, regroupV0_hi_lo_hi_lo_hi_lo_12};
  wire [127:0]       regroupV0_hi_lo_hi_lo_12 = {regroupV0_hi_lo_hi_lo_hi_12, regroupV0_hi_lo_hi_lo_lo_12};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo_lo_1 = {regroupV0_hi_12[1541], regroupV0_hi_12[1537]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo_hi_1 = {regroupV0_hi_12[1549], regroupV0_hi_12[1545]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo_5 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo_hi_1, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi_lo_1 = {regroupV0_hi_12[1557], regroupV0_hi_12[1553]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi_hi_1 = {regroupV0_hi_12[1565], regroupV0_hi_12[1561]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi_5 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi_hi_1, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_9 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi_5, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo_lo_1 = {regroupV0_hi_12[1573], regroupV0_hi_12[1569]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo_hi_1 = {regroupV0_hi_12[1581], regroupV0_hi_12[1577]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo_5 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo_hi_1, regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi_lo_1 = {regroupV0_hi_12[1589], regroupV0_hi_12[1585]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi_hi_1 = {regroupV0_hi_12[1597], regroupV0_hi_12[1593]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi_5 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi_hi_1, regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_9 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi_5, regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_lo_lo_12 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_9, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_9};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo_lo_1 = {regroupV0_hi_12[1605], regroupV0_hi_12[1601]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo_hi_1 = {regroupV0_hi_12[1613], regroupV0_hi_12[1609]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo_5 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo_hi_1, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi_lo_1 = {regroupV0_hi_12[1621], regroupV0_hi_12[1617]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi_hi_1 = {regroupV0_hi_12[1629], regroupV0_hi_12[1625]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi_5 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi_hi_1, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_9 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi_5, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo_lo_1 = {regroupV0_hi_12[1637], regroupV0_hi_12[1633]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo_hi_1 = {regroupV0_hi_12[1645], regroupV0_hi_12[1641]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo_5 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo_hi_1, regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi_lo_1 = {regroupV0_hi_12[1653], regroupV0_hi_12[1649]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi_hi_1 = {regroupV0_hi_12[1661], regroupV0_hi_12[1657]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi_5 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi_hi_1, regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_9 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi_5, regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_lo_hi_12 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_9, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_9};
  wire [31:0]        regroupV0_hi_lo_hi_hi_lo_lo_12 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_12, regroupV0_hi_lo_hi_hi_lo_lo_lo_12};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo_lo_1 = {regroupV0_hi_12[1669], regroupV0_hi_12[1665]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo_hi_1 = {regroupV0_hi_12[1677], regroupV0_hi_12[1673]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo_5 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo_hi_1, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi_lo_1 = {regroupV0_hi_12[1685], regroupV0_hi_12[1681]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi_hi_1 = {regroupV0_hi_12[1693], regroupV0_hi_12[1689]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi_5 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi_hi_1, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_9 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi_5, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo_lo_1 = {regroupV0_hi_12[1701], regroupV0_hi_12[1697]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo_hi_1 = {regroupV0_hi_12[1709], regroupV0_hi_12[1705]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo_5 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo_hi_1, regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi_lo_1 = {regroupV0_hi_12[1717], regroupV0_hi_12[1713]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi_hi_1 = {regroupV0_hi_12[1725], regroupV0_hi_12[1721]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi_5 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi_hi_1, regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_9 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi_5, regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_hi_lo_12 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_9, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_9};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo_lo_1 = {regroupV0_hi_12[1733], regroupV0_hi_12[1729]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo_hi_1 = {regroupV0_hi_12[1741], regroupV0_hi_12[1737]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo_5 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo_hi_1, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi_lo_1 = {regroupV0_hi_12[1749], regroupV0_hi_12[1745]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi_hi_1 = {regroupV0_hi_12[1757], regroupV0_hi_12[1753]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi_5 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi_hi_1, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_9 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi_5, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo_lo_1 = {regroupV0_hi_12[1765], regroupV0_hi_12[1761]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo_hi_1 = {regroupV0_hi_12[1773], regroupV0_hi_12[1769]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo_5 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo_hi_1, regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi_lo_1 = {regroupV0_hi_12[1781], regroupV0_hi_12[1777]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi_hi_1 = {regroupV0_hi_12[1789], regroupV0_hi_12[1785]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi_5 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi_hi_1, regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_9 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi_5, regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_hi_hi_12 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_9, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_9};
  wire [31:0]        regroupV0_hi_lo_hi_hi_lo_hi_12 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_12, regroupV0_hi_lo_hi_hi_lo_hi_lo_12};
  wire [63:0]        regroupV0_hi_lo_hi_hi_lo_12 = {regroupV0_hi_lo_hi_hi_lo_hi_12, regroupV0_hi_lo_hi_hi_lo_lo_12};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo_lo_1 = {regroupV0_hi_12[1797], regroupV0_hi_12[1793]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo_hi_1 = {regroupV0_hi_12[1805], regroupV0_hi_12[1801]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo_5 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo_hi_1, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi_lo_1 = {regroupV0_hi_12[1813], regroupV0_hi_12[1809]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi_hi_1 = {regroupV0_hi_12[1821], regroupV0_hi_12[1817]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi_5 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi_hi_1, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_9 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi_5, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo_lo_1 = {regroupV0_hi_12[1829], regroupV0_hi_12[1825]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo_hi_1 = {regroupV0_hi_12[1837], regroupV0_hi_12[1833]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo_5 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo_hi_1, regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi_lo_1 = {regroupV0_hi_12[1845], regroupV0_hi_12[1841]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi_hi_1 = {regroupV0_hi_12[1853], regroupV0_hi_12[1849]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi_5 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi_hi_1, regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_9 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi_5, regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_lo_lo_12 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_9, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_9};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo_lo_1 = {regroupV0_hi_12[1861], regroupV0_hi_12[1857]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo_hi_1 = {regroupV0_hi_12[1869], regroupV0_hi_12[1865]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo_5 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo_hi_1, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi_lo_1 = {regroupV0_hi_12[1877], regroupV0_hi_12[1873]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi_hi_1 = {regroupV0_hi_12[1885], regroupV0_hi_12[1881]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi_5 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi_hi_1, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_9 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi_5, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo_lo_1 = {regroupV0_hi_12[1893], regroupV0_hi_12[1889]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo_hi_1 = {regroupV0_hi_12[1901], regroupV0_hi_12[1897]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo_5 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo_hi_1, regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi_lo_1 = {regroupV0_hi_12[1909], regroupV0_hi_12[1905]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi_hi_1 = {regroupV0_hi_12[1917], regroupV0_hi_12[1913]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi_5 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi_hi_1, regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_9 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi_5, regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_lo_hi_12 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_9, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_9};
  wire [31:0]        regroupV0_hi_lo_hi_hi_hi_lo_12 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_12, regroupV0_hi_lo_hi_hi_hi_lo_lo_12};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo_lo_1 = {regroupV0_hi_12[1925], regroupV0_hi_12[1921]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo_hi_1 = {regroupV0_hi_12[1933], regroupV0_hi_12[1929]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo_5 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo_hi_1, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi_lo_1 = {regroupV0_hi_12[1941], regroupV0_hi_12[1937]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi_hi_1 = {regroupV0_hi_12[1949], regroupV0_hi_12[1945]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi_5 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi_hi_1, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_9 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi_5, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo_lo_1 = {regroupV0_hi_12[1957], regroupV0_hi_12[1953]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo_hi_1 = {regroupV0_hi_12[1965], regroupV0_hi_12[1961]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo_5 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo_hi_1, regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi_lo_1 = {regroupV0_hi_12[1973], regroupV0_hi_12[1969]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi_hi_1 = {regroupV0_hi_12[1981], regroupV0_hi_12[1977]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi_5 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi_hi_1, regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_9 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi_5, regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_hi_lo_12 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_9, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_9};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo_lo_1 = {regroupV0_hi_12[1989], regroupV0_hi_12[1985]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo_hi_1 = {regroupV0_hi_12[1997], regroupV0_hi_12[1993]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo_5 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo_hi_1, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi_lo_1 = {regroupV0_hi_12[2005], regroupV0_hi_12[2001]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi_hi_1 = {regroupV0_hi_12[2013], regroupV0_hi_12[2009]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi_5 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi_hi_1, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_9 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi_5, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo_lo_1 = {regroupV0_hi_12[2021], regroupV0_hi_12[2017]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo_hi_1 = {regroupV0_hi_12[2029], regroupV0_hi_12[2025]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo_5 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo_hi_1, regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi_lo_1 = {regroupV0_hi_12[2037], regroupV0_hi_12[2033]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi_hi_1 = {regroupV0_hi_12[2045], regroupV0_hi_12[2041]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi_5 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi_hi_1, regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_9 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi_5, regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_hi_hi_12 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_9, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_9};
  wire [31:0]        regroupV0_hi_lo_hi_hi_hi_hi_12 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_12, regroupV0_hi_lo_hi_hi_hi_hi_lo_12};
  wire [63:0]        regroupV0_hi_lo_hi_hi_hi_12 = {regroupV0_hi_lo_hi_hi_hi_hi_12, regroupV0_hi_lo_hi_hi_hi_lo_12};
  wire [127:0]       regroupV0_hi_lo_hi_hi_12 = {regroupV0_hi_lo_hi_hi_hi_12, regroupV0_hi_lo_hi_hi_lo_12};
  wire [255:0]       regroupV0_hi_lo_hi_12 = {regroupV0_hi_lo_hi_hi_12, regroupV0_hi_lo_hi_lo_12};
  wire [511:0]       regroupV0_hi_lo_12 = {regroupV0_hi_lo_hi_12, regroupV0_hi_lo_lo_12};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo_lo_1 = {regroupV0_hi_12[2053], regroupV0_hi_12[2049]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo_hi_1 = {regroupV0_hi_12[2061], regroupV0_hi_12[2057]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo_5 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo_hi_1, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi_lo_1 = {regroupV0_hi_12[2069], regroupV0_hi_12[2065]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi_hi_1 = {regroupV0_hi_12[2077], regroupV0_hi_12[2073]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi_5 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi_hi_1, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_9 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi_5, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo_lo_1 = {regroupV0_hi_12[2085], regroupV0_hi_12[2081]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo_hi_1 = {regroupV0_hi_12[2093], regroupV0_hi_12[2089]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo_5 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo_hi_1, regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi_lo_1 = {regroupV0_hi_12[2101], regroupV0_hi_12[2097]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi_hi_1 = {regroupV0_hi_12[2109], regroupV0_hi_12[2105]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi_5 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi_hi_1, regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_9 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi_5, regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_lo_lo_12 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_9, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_9};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo_lo_1 = {regroupV0_hi_12[2117], regroupV0_hi_12[2113]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo_hi_1 = {regroupV0_hi_12[2125], regroupV0_hi_12[2121]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo_5 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo_hi_1, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi_lo_1 = {regroupV0_hi_12[2133], regroupV0_hi_12[2129]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi_hi_1 = {regroupV0_hi_12[2141], regroupV0_hi_12[2137]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi_5 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi_hi_1, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_9 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi_5, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo_lo_1 = {regroupV0_hi_12[2149], regroupV0_hi_12[2145]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo_hi_1 = {regroupV0_hi_12[2157], regroupV0_hi_12[2153]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo_5 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo_hi_1, regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi_lo_1 = {regroupV0_hi_12[2165], regroupV0_hi_12[2161]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi_hi_1 = {regroupV0_hi_12[2173], regroupV0_hi_12[2169]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi_5 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi_hi_1, regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_9 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi_5, regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_lo_hi_12 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_9, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_9};
  wire [31:0]        regroupV0_hi_hi_lo_lo_lo_lo_12 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_12, regroupV0_hi_hi_lo_lo_lo_lo_lo_12};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo_lo_1 = {regroupV0_hi_12[2181], regroupV0_hi_12[2177]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo_hi_1 = {regroupV0_hi_12[2189], regroupV0_hi_12[2185]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo_5 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo_hi_1, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi_lo_1 = {regroupV0_hi_12[2197], regroupV0_hi_12[2193]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi_hi_1 = {regroupV0_hi_12[2205], regroupV0_hi_12[2201]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi_5 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi_hi_1, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_9 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi_5, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo_lo_1 = {regroupV0_hi_12[2213], regroupV0_hi_12[2209]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo_hi_1 = {regroupV0_hi_12[2221], regroupV0_hi_12[2217]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo_5 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo_hi_1, regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi_lo_1 = {regroupV0_hi_12[2229], regroupV0_hi_12[2225]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi_hi_1 = {regroupV0_hi_12[2237], regroupV0_hi_12[2233]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi_5 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi_hi_1, regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_9 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi_5, regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_hi_lo_12 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_9, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_9};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo_lo_1 = {regroupV0_hi_12[2245], regroupV0_hi_12[2241]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo_hi_1 = {regroupV0_hi_12[2253], regroupV0_hi_12[2249]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo_5 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo_hi_1, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi_lo_1 = {regroupV0_hi_12[2261], regroupV0_hi_12[2257]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi_hi_1 = {regroupV0_hi_12[2269], regroupV0_hi_12[2265]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi_5 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi_hi_1, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_9 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi_5, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo_lo_1 = {regroupV0_hi_12[2277], regroupV0_hi_12[2273]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo_hi_1 = {regroupV0_hi_12[2285], regroupV0_hi_12[2281]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo_5 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo_hi_1, regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi_lo_1 = {regroupV0_hi_12[2293], regroupV0_hi_12[2289]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi_hi_1 = {regroupV0_hi_12[2301], regroupV0_hi_12[2297]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi_5 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi_hi_1, regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_9 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi_5, regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_hi_hi_12 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_9, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_9};
  wire [31:0]        regroupV0_hi_hi_lo_lo_lo_hi_12 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_12, regroupV0_hi_hi_lo_lo_lo_hi_lo_12};
  wire [63:0]        regroupV0_hi_hi_lo_lo_lo_12 = {regroupV0_hi_hi_lo_lo_lo_hi_12, regroupV0_hi_hi_lo_lo_lo_lo_12};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo_lo_1 = {regroupV0_hi_12[2309], regroupV0_hi_12[2305]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo_hi_1 = {regroupV0_hi_12[2317], regroupV0_hi_12[2313]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo_5 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo_hi_1, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi_lo_1 = {regroupV0_hi_12[2325], regroupV0_hi_12[2321]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi_hi_1 = {regroupV0_hi_12[2333], regroupV0_hi_12[2329]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi_5 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi_hi_1, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_9 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi_5, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo_lo_1 = {regroupV0_hi_12[2341], regroupV0_hi_12[2337]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo_hi_1 = {regroupV0_hi_12[2349], regroupV0_hi_12[2345]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo_5 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo_hi_1, regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi_lo_1 = {regroupV0_hi_12[2357], regroupV0_hi_12[2353]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi_hi_1 = {regroupV0_hi_12[2365], regroupV0_hi_12[2361]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi_5 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi_hi_1, regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_9 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi_5, regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_lo_lo_12 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_9, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_9};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo_lo_1 = {regroupV0_hi_12[2373], regroupV0_hi_12[2369]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo_hi_1 = {regroupV0_hi_12[2381], regroupV0_hi_12[2377]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo_5 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo_hi_1, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi_lo_1 = {regroupV0_hi_12[2389], regroupV0_hi_12[2385]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi_hi_1 = {regroupV0_hi_12[2397], regroupV0_hi_12[2393]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi_5 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi_hi_1, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_9 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi_5, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo_lo_1 = {regroupV0_hi_12[2405], regroupV0_hi_12[2401]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo_hi_1 = {regroupV0_hi_12[2413], regroupV0_hi_12[2409]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo_5 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo_hi_1, regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi_lo_1 = {regroupV0_hi_12[2421], regroupV0_hi_12[2417]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi_hi_1 = {regroupV0_hi_12[2429], regroupV0_hi_12[2425]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi_5 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi_hi_1, regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_9 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi_5, regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_lo_hi_12 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_9, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_9};
  wire [31:0]        regroupV0_hi_hi_lo_lo_hi_lo_12 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_12, regroupV0_hi_hi_lo_lo_hi_lo_lo_12};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo_lo_1 = {regroupV0_hi_12[2437], regroupV0_hi_12[2433]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo_hi_1 = {regroupV0_hi_12[2445], regroupV0_hi_12[2441]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo_5 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo_hi_1, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi_lo_1 = {regroupV0_hi_12[2453], regroupV0_hi_12[2449]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi_hi_1 = {regroupV0_hi_12[2461], regroupV0_hi_12[2457]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi_5 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi_hi_1, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_9 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi_5, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo_lo_1 = {regroupV0_hi_12[2469], regroupV0_hi_12[2465]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo_hi_1 = {regroupV0_hi_12[2477], regroupV0_hi_12[2473]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo_5 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo_hi_1, regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi_lo_1 = {regroupV0_hi_12[2485], regroupV0_hi_12[2481]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi_hi_1 = {regroupV0_hi_12[2493], regroupV0_hi_12[2489]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi_5 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi_hi_1, regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_9 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi_5, regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_hi_lo_12 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_9, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_9};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo_lo_1 = {regroupV0_hi_12[2501], regroupV0_hi_12[2497]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo_hi_1 = {regroupV0_hi_12[2509], regroupV0_hi_12[2505]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo_5 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo_hi_1, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi_lo_1 = {regroupV0_hi_12[2517], regroupV0_hi_12[2513]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi_hi_1 = {regroupV0_hi_12[2525], regroupV0_hi_12[2521]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi_5 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi_hi_1, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_9 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi_5, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo_lo_1 = {regroupV0_hi_12[2533], regroupV0_hi_12[2529]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo_hi_1 = {regroupV0_hi_12[2541], regroupV0_hi_12[2537]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo_5 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo_hi_1, regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi_lo_1 = {regroupV0_hi_12[2549], regroupV0_hi_12[2545]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi_hi_1 = {regroupV0_hi_12[2557], regroupV0_hi_12[2553]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi_5 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi_hi_1, regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_9 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi_5, regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_hi_hi_12 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_9, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_9};
  wire [31:0]        regroupV0_hi_hi_lo_lo_hi_hi_12 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_12, regroupV0_hi_hi_lo_lo_hi_hi_lo_12};
  wire [63:0]        regroupV0_hi_hi_lo_lo_hi_12 = {regroupV0_hi_hi_lo_lo_hi_hi_12, regroupV0_hi_hi_lo_lo_hi_lo_12};
  wire [127:0]       regroupV0_hi_hi_lo_lo_12 = {regroupV0_hi_hi_lo_lo_hi_12, regroupV0_hi_hi_lo_lo_lo_12};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo_lo_1 = {regroupV0_hi_12[2565], regroupV0_hi_12[2561]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo_hi_1 = {regroupV0_hi_12[2573], regroupV0_hi_12[2569]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo_5 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo_hi_1, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi_lo_1 = {regroupV0_hi_12[2581], regroupV0_hi_12[2577]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi_hi_1 = {regroupV0_hi_12[2589], regroupV0_hi_12[2585]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi_5 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi_hi_1, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_9 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi_5, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo_lo_1 = {regroupV0_hi_12[2597], regroupV0_hi_12[2593]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo_hi_1 = {regroupV0_hi_12[2605], regroupV0_hi_12[2601]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo_5 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo_hi_1, regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi_lo_1 = {regroupV0_hi_12[2613], regroupV0_hi_12[2609]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi_hi_1 = {regroupV0_hi_12[2621], regroupV0_hi_12[2617]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi_5 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi_hi_1, regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_9 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi_5, regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_lo_lo_12 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_9, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_9};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo_lo_1 = {regroupV0_hi_12[2629], regroupV0_hi_12[2625]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo_hi_1 = {regroupV0_hi_12[2637], regroupV0_hi_12[2633]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo_5 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo_hi_1, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi_lo_1 = {regroupV0_hi_12[2645], regroupV0_hi_12[2641]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi_hi_1 = {regroupV0_hi_12[2653], regroupV0_hi_12[2649]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi_5 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi_hi_1, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_9 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi_5, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo_lo_1 = {regroupV0_hi_12[2661], regroupV0_hi_12[2657]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo_hi_1 = {regroupV0_hi_12[2669], regroupV0_hi_12[2665]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo_5 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo_hi_1, regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi_lo_1 = {regroupV0_hi_12[2677], regroupV0_hi_12[2673]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi_hi_1 = {regroupV0_hi_12[2685], regroupV0_hi_12[2681]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi_5 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi_hi_1, regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_9 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi_5, regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_lo_hi_12 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_9, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_9};
  wire [31:0]        regroupV0_hi_hi_lo_hi_lo_lo_12 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_12, regroupV0_hi_hi_lo_hi_lo_lo_lo_12};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo_lo_1 = {regroupV0_hi_12[2693], regroupV0_hi_12[2689]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo_hi_1 = {regroupV0_hi_12[2701], regroupV0_hi_12[2697]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo_5 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo_hi_1, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi_lo_1 = {regroupV0_hi_12[2709], regroupV0_hi_12[2705]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi_hi_1 = {regroupV0_hi_12[2717], regroupV0_hi_12[2713]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi_5 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi_hi_1, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_9 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi_5, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo_lo_1 = {regroupV0_hi_12[2725], regroupV0_hi_12[2721]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo_hi_1 = {regroupV0_hi_12[2733], regroupV0_hi_12[2729]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo_5 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo_hi_1, regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi_lo_1 = {regroupV0_hi_12[2741], regroupV0_hi_12[2737]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi_hi_1 = {regroupV0_hi_12[2749], regroupV0_hi_12[2745]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi_5 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi_hi_1, regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_9 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi_5, regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_hi_lo_12 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_9, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_9};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo_lo_1 = {regroupV0_hi_12[2757], regroupV0_hi_12[2753]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo_hi_1 = {regroupV0_hi_12[2765], regroupV0_hi_12[2761]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo_5 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo_hi_1, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi_lo_1 = {regroupV0_hi_12[2773], regroupV0_hi_12[2769]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi_hi_1 = {regroupV0_hi_12[2781], regroupV0_hi_12[2777]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi_5 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi_hi_1, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_9 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi_5, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo_lo_1 = {regroupV0_hi_12[2789], regroupV0_hi_12[2785]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo_hi_1 = {regroupV0_hi_12[2797], regroupV0_hi_12[2793]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo_5 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo_hi_1, regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi_lo_1 = {regroupV0_hi_12[2805], regroupV0_hi_12[2801]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi_hi_1 = {regroupV0_hi_12[2813], regroupV0_hi_12[2809]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi_5 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi_hi_1, regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_9 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi_5, regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_hi_hi_12 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_9, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_9};
  wire [31:0]        regroupV0_hi_hi_lo_hi_lo_hi_12 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_12, regroupV0_hi_hi_lo_hi_lo_hi_lo_12};
  wire [63:0]        regroupV0_hi_hi_lo_hi_lo_12 = {regroupV0_hi_hi_lo_hi_lo_hi_12, regroupV0_hi_hi_lo_hi_lo_lo_12};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo_lo_1 = {regroupV0_hi_12[2821], regroupV0_hi_12[2817]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo_hi_1 = {regroupV0_hi_12[2829], regroupV0_hi_12[2825]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo_5 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo_hi_1, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi_lo_1 = {regroupV0_hi_12[2837], regroupV0_hi_12[2833]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi_hi_1 = {regroupV0_hi_12[2845], regroupV0_hi_12[2841]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi_5 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi_hi_1, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_9 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi_5, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo_lo_1 = {regroupV0_hi_12[2853], regroupV0_hi_12[2849]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo_hi_1 = {regroupV0_hi_12[2861], regroupV0_hi_12[2857]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo_5 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo_hi_1, regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi_lo_1 = {regroupV0_hi_12[2869], regroupV0_hi_12[2865]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi_hi_1 = {regroupV0_hi_12[2877], regroupV0_hi_12[2873]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi_5 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi_hi_1, regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_9 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi_5, regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_lo_lo_12 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_9, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_9};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo_lo_1 = {regroupV0_hi_12[2885], regroupV0_hi_12[2881]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo_hi_1 = {regroupV0_hi_12[2893], regroupV0_hi_12[2889]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo_5 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo_hi_1, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi_lo_1 = {regroupV0_hi_12[2901], regroupV0_hi_12[2897]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi_hi_1 = {regroupV0_hi_12[2909], regroupV0_hi_12[2905]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi_5 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi_hi_1, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_9 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi_5, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo_lo_1 = {regroupV0_hi_12[2917], regroupV0_hi_12[2913]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo_hi_1 = {regroupV0_hi_12[2925], regroupV0_hi_12[2921]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo_5 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo_hi_1, regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi_lo_1 = {regroupV0_hi_12[2933], regroupV0_hi_12[2929]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi_hi_1 = {regroupV0_hi_12[2941], regroupV0_hi_12[2937]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi_5 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi_hi_1, regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_9 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi_5, regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_lo_hi_12 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_9, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_9};
  wire [31:0]        regroupV0_hi_hi_lo_hi_hi_lo_12 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_12, regroupV0_hi_hi_lo_hi_hi_lo_lo_12};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo_lo_1 = {regroupV0_hi_12[2949], regroupV0_hi_12[2945]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo_hi_1 = {regroupV0_hi_12[2957], regroupV0_hi_12[2953]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo_5 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo_hi_1, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi_lo_1 = {regroupV0_hi_12[2965], regroupV0_hi_12[2961]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi_hi_1 = {regroupV0_hi_12[2973], regroupV0_hi_12[2969]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi_5 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi_hi_1, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_9 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi_5, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo_lo_1 = {regroupV0_hi_12[2981], regroupV0_hi_12[2977]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo_hi_1 = {regroupV0_hi_12[2989], regroupV0_hi_12[2985]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo_5 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo_hi_1, regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi_lo_1 = {regroupV0_hi_12[2997], regroupV0_hi_12[2993]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi_hi_1 = {regroupV0_hi_12[3005], regroupV0_hi_12[3001]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi_5 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi_hi_1, regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_9 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi_5, regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_hi_lo_12 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_9, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_9};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo_lo_1 = {regroupV0_hi_12[3013], regroupV0_hi_12[3009]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo_hi_1 = {regroupV0_hi_12[3021], regroupV0_hi_12[3017]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo_5 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo_hi_1, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi_lo_1 = {regroupV0_hi_12[3029], regroupV0_hi_12[3025]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi_hi_1 = {regroupV0_hi_12[3037], regroupV0_hi_12[3033]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi_5 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi_hi_1, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_9 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi_5, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo_lo_1 = {regroupV0_hi_12[3045], regroupV0_hi_12[3041]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo_hi_1 = {regroupV0_hi_12[3053], regroupV0_hi_12[3049]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo_5 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo_hi_1, regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi_lo_1 = {regroupV0_hi_12[3061], regroupV0_hi_12[3057]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi_hi_1 = {regroupV0_hi_12[3069], regroupV0_hi_12[3065]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi_5 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi_hi_1, regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_9 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi_5, regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_hi_hi_12 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_9, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_9};
  wire [31:0]        regroupV0_hi_hi_lo_hi_hi_hi_12 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_12, regroupV0_hi_hi_lo_hi_hi_hi_lo_12};
  wire [63:0]        regroupV0_hi_hi_lo_hi_hi_12 = {regroupV0_hi_hi_lo_hi_hi_hi_12, regroupV0_hi_hi_lo_hi_hi_lo_12};
  wire [127:0]       regroupV0_hi_hi_lo_hi_12 = {regroupV0_hi_hi_lo_hi_hi_12, regroupV0_hi_hi_lo_hi_lo_12};
  wire [255:0]       regroupV0_hi_hi_lo_12 = {regroupV0_hi_hi_lo_hi_12, regroupV0_hi_hi_lo_lo_12};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo_lo_1 = {regroupV0_hi_12[3077], regroupV0_hi_12[3073]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo_hi_1 = {regroupV0_hi_12[3085], regroupV0_hi_12[3081]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo_5 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo_hi_1, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi_lo_1 = {regroupV0_hi_12[3093], regroupV0_hi_12[3089]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi_hi_1 = {regroupV0_hi_12[3101], regroupV0_hi_12[3097]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi_5 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi_hi_1, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_9 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi_5, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo_lo_1 = {regroupV0_hi_12[3109], regroupV0_hi_12[3105]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo_hi_1 = {regroupV0_hi_12[3117], regroupV0_hi_12[3113]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo_5 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo_hi_1, regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi_lo_1 = {regroupV0_hi_12[3125], regroupV0_hi_12[3121]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi_hi_1 = {regroupV0_hi_12[3133], regroupV0_hi_12[3129]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi_5 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi_hi_1, regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_9 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi_5, regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_lo_lo_12 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_9, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_9};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo_lo_1 = {regroupV0_hi_12[3141], regroupV0_hi_12[3137]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo_hi_1 = {regroupV0_hi_12[3149], regroupV0_hi_12[3145]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo_5 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo_hi_1, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi_lo_1 = {regroupV0_hi_12[3157], regroupV0_hi_12[3153]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi_hi_1 = {regroupV0_hi_12[3165], regroupV0_hi_12[3161]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi_5 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi_hi_1, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_9 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi_5, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo_lo_1 = {regroupV0_hi_12[3173], regroupV0_hi_12[3169]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo_hi_1 = {regroupV0_hi_12[3181], regroupV0_hi_12[3177]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo_5 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo_hi_1, regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi_lo_1 = {regroupV0_hi_12[3189], regroupV0_hi_12[3185]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi_hi_1 = {regroupV0_hi_12[3197], regroupV0_hi_12[3193]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi_5 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_9 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi_5, regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_lo_hi_12 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_9, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_9};
  wire [31:0]        regroupV0_hi_hi_hi_lo_lo_lo_12 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_12, regroupV0_hi_hi_hi_lo_lo_lo_lo_12};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo_lo_1 = {regroupV0_hi_12[3205], regroupV0_hi_12[3201]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo_hi_1 = {regroupV0_hi_12[3213], regroupV0_hi_12[3209]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo_5 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo_hi_1, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi_lo_1 = {regroupV0_hi_12[3221], regroupV0_hi_12[3217]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi_hi_1 = {regroupV0_hi_12[3229], regroupV0_hi_12[3225]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi_5 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi_hi_1, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_9 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi_5, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo_lo_1 = {regroupV0_hi_12[3237], regroupV0_hi_12[3233]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo_hi_1 = {regroupV0_hi_12[3245], regroupV0_hi_12[3241]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo_5 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo_hi_1, regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi_lo_1 = {regroupV0_hi_12[3253], regroupV0_hi_12[3249]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi_hi_1 = {regroupV0_hi_12[3261], regroupV0_hi_12[3257]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi_5 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi_hi_1, regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_9 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi_5, regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_hi_lo_12 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_9, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_9};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo_lo_1 = {regroupV0_hi_12[3269], regroupV0_hi_12[3265]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo_hi_1 = {regroupV0_hi_12[3277], regroupV0_hi_12[3273]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo_5 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo_hi_1, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi_lo_1 = {regroupV0_hi_12[3285], regroupV0_hi_12[3281]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi_hi_1 = {regroupV0_hi_12[3293], regroupV0_hi_12[3289]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi_5 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi_hi_1, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_9 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi_5, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo_lo_1 = {regroupV0_hi_12[3301], regroupV0_hi_12[3297]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo_hi_1 = {regroupV0_hi_12[3309], regroupV0_hi_12[3305]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo_5 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo_hi_1, regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi_lo_1 = {regroupV0_hi_12[3317], regroupV0_hi_12[3313]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi_hi_1 = {regroupV0_hi_12[3325], regroupV0_hi_12[3321]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi_5 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_9 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi_5, regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_hi_hi_12 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_9, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_9};
  wire [31:0]        regroupV0_hi_hi_hi_lo_lo_hi_12 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_12, regroupV0_hi_hi_hi_lo_lo_hi_lo_12};
  wire [63:0]        regroupV0_hi_hi_hi_lo_lo_12 = {regroupV0_hi_hi_hi_lo_lo_hi_12, regroupV0_hi_hi_hi_lo_lo_lo_12};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo_lo_1 = {regroupV0_hi_12[3333], regroupV0_hi_12[3329]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo_hi_1 = {regroupV0_hi_12[3341], regroupV0_hi_12[3337]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo_5 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo_hi_1, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi_lo_1 = {regroupV0_hi_12[3349], regroupV0_hi_12[3345]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi_hi_1 = {regroupV0_hi_12[3357], regroupV0_hi_12[3353]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi_5 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi_hi_1, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_9 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi_5, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo_lo_1 = {regroupV0_hi_12[3365], regroupV0_hi_12[3361]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo_hi_1 = {regroupV0_hi_12[3373], regroupV0_hi_12[3369]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo_5 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo_hi_1, regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi_lo_1 = {regroupV0_hi_12[3381], regroupV0_hi_12[3377]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi_hi_1 = {regroupV0_hi_12[3389], regroupV0_hi_12[3385]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi_5 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi_hi_1, regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_9 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi_5, regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_lo_lo_12 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_9, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_9};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo_lo_1 = {regroupV0_hi_12[3397], regroupV0_hi_12[3393]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo_hi_1 = {regroupV0_hi_12[3405], regroupV0_hi_12[3401]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo_5 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo_hi_1, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi_lo_1 = {regroupV0_hi_12[3413], regroupV0_hi_12[3409]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi_hi_1 = {regroupV0_hi_12[3421], regroupV0_hi_12[3417]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi_5 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi_hi_1, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_9 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi_5, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo_lo_1 = {regroupV0_hi_12[3429], regroupV0_hi_12[3425]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo_hi_1 = {regroupV0_hi_12[3437], regroupV0_hi_12[3433]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo_5 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo_hi_1, regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi_lo_1 = {regroupV0_hi_12[3445], regroupV0_hi_12[3441]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi_hi_1 = {regroupV0_hi_12[3453], regroupV0_hi_12[3449]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi_5 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_9 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi_5, regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_lo_hi_12 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_9, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_9};
  wire [31:0]        regroupV0_hi_hi_hi_lo_hi_lo_12 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_12, regroupV0_hi_hi_hi_lo_hi_lo_lo_12};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo_lo_1 = {regroupV0_hi_12[3461], regroupV0_hi_12[3457]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo_hi_1 = {regroupV0_hi_12[3469], regroupV0_hi_12[3465]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo_5 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo_hi_1, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi_lo_1 = {regroupV0_hi_12[3477], regroupV0_hi_12[3473]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi_hi_1 = {regroupV0_hi_12[3485], regroupV0_hi_12[3481]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi_5 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi_hi_1, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_9 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi_5, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo_lo_1 = {regroupV0_hi_12[3493], regroupV0_hi_12[3489]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo_hi_1 = {regroupV0_hi_12[3501], regroupV0_hi_12[3497]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo_5 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo_hi_1, regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi_lo_1 = {regroupV0_hi_12[3509], regroupV0_hi_12[3505]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi_hi_1 = {regroupV0_hi_12[3517], regroupV0_hi_12[3513]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi_5 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi_hi_1, regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_9 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi_5, regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_hi_lo_12 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_9, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_9};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo_lo_1 = {regroupV0_hi_12[3525], regroupV0_hi_12[3521]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo_hi_1 = {regroupV0_hi_12[3533], regroupV0_hi_12[3529]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo_5 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo_hi_1, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi_lo_1 = {regroupV0_hi_12[3541], regroupV0_hi_12[3537]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi_hi_1 = {regroupV0_hi_12[3549], regroupV0_hi_12[3545]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi_5 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi_hi_1, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_9 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi_5, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo_lo_1 = {regroupV0_hi_12[3557], regroupV0_hi_12[3553]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo_hi_1 = {regroupV0_hi_12[3565], regroupV0_hi_12[3561]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo_5 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo_hi_1, regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi_lo_1 = {regroupV0_hi_12[3573], regroupV0_hi_12[3569]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi_hi_1 = {regroupV0_hi_12[3581], regroupV0_hi_12[3577]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi_5 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_9 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi_5, regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_hi_hi_12 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_9, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_9};
  wire [31:0]        regroupV0_hi_hi_hi_lo_hi_hi_12 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_12, regroupV0_hi_hi_hi_lo_hi_hi_lo_12};
  wire [63:0]        regroupV0_hi_hi_hi_lo_hi_12 = {regroupV0_hi_hi_hi_lo_hi_hi_12, regroupV0_hi_hi_hi_lo_hi_lo_12};
  wire [127:0]       regroupV0_hi_hi_hi_lo_12 = {regroupV0_hi_hi_hi_lo_hi_12, regroupV0_hi_hi_hi_lo_lo_12};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo_lo_1 = {regroupV0_hi_12[3589], regroupV0_hi_12[3585]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo_hi_1 = {regroupV0_hi_12[3597], regroupV0_hi_12[3593]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo_5 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo_hi_1, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi_lo_1 = {regroupV0_hi_12[3605], regroupV0_hi_12[3601]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi_hi_1 = {regroupV0_hi_12[3613], regroupV0_hi_12[3609]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi_5 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi_hi_1, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_9 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi_5, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo_lo_1 = {regroupV0_hi_12[3621], regroupV0_hi_12[3617]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo_hi_1 = {regroupV0_hi_12[3629], regroupV0_hi_12[3625]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo_5 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo_hi_1, regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi_lo_1 = {regroupV0_hi_12[3637], regroupV0_hi_12[3633]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi_hi_1 = {regroupV0_hi_12[3645], regroupV0_hi_12[3641]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi_5 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi_hi_1, regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_9 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi_5, regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_lo_lo_12 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_9, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_9};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo_lo_1 = {regroupV0_hi_12[3653], regroupV0_hi_12[3649]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo_hi_1 = {regroupV0_hi_12[3661], regroupV0_hi_12[3657]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo_5 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo_hi_1, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi_lo_1 = {regroupV0_hi_12[3669], regroupV0_hi_12[3665]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi_hi_1 = {regroupV0_hi_12[3677], regroupV0_hi_12[3673]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi_5 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi_hi_1, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_9 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi_5, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo_lo_1 = {regroupV0_hi_12[3685], regroupV0_hi_12[3681]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo_hi_1 = {regroupV0_hi_12[3693], regroupV0_hi_12[3689]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo_5 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo_hi_1, regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi_lo_1 = {regroupV0_hi_12[3701], regroupV0_hi_12[3697]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi_hi_1 = {regroupV0_hi_12[3709], regroupV0_hi_12[3705]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi_5 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_9 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi_5, regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_lo_hi_12 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_9, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_9};
  wire [31:0]        regroupV0_hi_hi_hi_hi_lo_lo_12 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_12, regroupV0_hi_hi_hi_hi_lo_lo_lo_12};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo_lo_1 = {regroupV0_hi_12[3717], regroupV0_hi_12[3713]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo_hi_1 = {regroupV0_hi_12[3725], regroupV0_hi_12[3721]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo_5 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo_hi_1, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi_lo_1 = {regroupV0_hi_12[3733], regroupV0_hi_12[3729]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi_hi_1 = {regroupV0_hi_12[3741], regroupV0_hi_12[3737]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi_5 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi_hi_1, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_9 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi_5, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo_lo_1 = {regroupV0_hi_12[3749], regroupV0_hi_12[3745]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo_hi_1 = {regroupV0_hi_12[3757], regroupV0_hi_12[3753]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo_5 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo_hi_1, regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi_lo_1 = {regroupV0_hi_12[3765], regroupV0_hi_12[3761]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi_hi_1 = {regroupV0_hi_12[3773], regroupV0_hi_12[3769]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi_5 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi_hi_1, regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_9 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi_5, regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_hi_lo_12 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_9, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_9};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo_lo_1 = {regroupV0_hi_12[3781], regroupV0_hi_12[3777]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo_hi_1 = {regroupV0_hi_12[3789], regroupV0_hi_12[3785]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo_5 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo_hi_1, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi_lo_1 = {regroupV0_hi_12[3797], regroupV0_hi_12[3793]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi_hi_1 = {regroupV0_hi_12[3805], regroupV0_hi_12[3801]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi_5 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi_hi_1, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_9 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi_5, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo_lo_1 = {regroupV0_hi_12[3813], regroupV0_hi_12[3809]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo_hi_1 = {regroupV0_hi_12[3821], regroupV0_hi_12[3817]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo_5 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo_hi_1, regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi_lo_1 = {regroupV0_hi_12[3829], regroupV0_hi_12[3825]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi_hi_1 = {regroupV0_hi_12[3837], regroupV0_hi_12[3833]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi_5 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_9 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi_5, regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_hi_hi_12 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_9, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_9};
  wire [31:0]        regroupV0_hi_hi_hi_hi_lo_hi_12 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_12, regroupV0_hi_hi_hi_hi_lo_hi_lo_12};
  wire [63:0]        regroupV0_hi_hi_hi_hi_lo_12 = {regroupV0_hi_hi_hi_hi_lo_hi_12, regroupV0_hi_hi_hi_hi_lo_lo_12};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo_lo_1 = {regroupV0_hi_12[3845], regroupV0_hi_12[3841]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo_hi_1 = {regroupV0_hi_12[3853], regroupV0_hi_12[3849]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo_5 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo_hi_1, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi_lo_1 = {regroupV0_hi_12[3861], regroupV0_hi_12[3857]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi_hi_1 = {regroupV0_hi_12[3869], regroupV0_hi_12[3865]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi_5 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi_hi_1, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_9 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi_5, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo_lo_1 = {regroupV0_hi_12[3877], regroupV0_hi_12[3873]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo_hi_1 = {regroupV0_hi_12[3885], regroupV0_hi_12[3881]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo_5 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo_hi_1, regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi_lo_1 = {regroupV0_hi_12[3893], regroupV0_hi_12[3889]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi_hi_1 = {regroupV0_hi_12[3901], regroupV0_hi_12[3897]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi_5 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi_hi_1, regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_9 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi_5, regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_lo_lo_12 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_9, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_9};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo_lo_1 = {regroupV0_hi_12[3909], regroupV0_hi_12[3905]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo_hi_1 = {regroupV0_hi_12[3917], regroupV0_hi_12[3913]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo_5 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo_hi_1, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi_lo_1 = {regroupV0_hi_12[3925], regroupV0_hi_12[3921]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi_hi_1 = {regroupV0_hi_12[3933], regroupV0_hi_12[3929]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi_5 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi_hi_1, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_9 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi_5, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo_lo_1 = {regroupV0_hi_12[3941], regroupV0_hi_12[3937]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo_hi_1 = {regroupV0_hi_12[3949], regroupV0_hi_12[3945]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo_5 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo_hi_1, regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi_lo_1 = {regroupV0_hi_12[3957], regroupV0_hi_12[3953]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi_hi_1 = {regroupV0_hi_12[3965], regroupV0_hi_12[3961]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi_5 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_9 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi_5, regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_lo_hi_12 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_9, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_9};
  wire [31:0]        regroupV0_hi_hi_hi_hi_hi_lo_12 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_12, regroupV0_hi_hi_hi_hi_hi_lo_lo_12};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo_lo_1 = {regroupV0_hi_12[3973], regroupV0_hi_12[3969]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo_hi_1 = {regroupV0_hi_12[3981], regroupV0_hi_12[3977]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo_5 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo_hi_1, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi_lo_1 = {regroupV0_hi_12[3989], regroupV0_hi_12[3985]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi_hi_1 = {regroupV0_hi_12[3997], regroupV0_hi_12[3993]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi_5 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi_hi_1, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_9 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi_5, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo_lo_1 = {regroupV0_hi_12[4005], regroupV0_hi_12[4001]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo_hi_1 = {regroupV0_hi_12[4013], regroupV0_hi_12[4009]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo_5 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo_hi_1, regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi_lo_1 = {regroupV0_hi_12[4021], regroupV0_hi_12[4017]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi_hi_1 = {regroupV0_hi_12[4029], regroupV0_hi_12[4025]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi_5 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi_hi_1, regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_9 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi_5, regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_hi_lo_12 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_9, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_9};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo_lo_1 = {regroupV0_hi_12[4037], regroupV0_hi_12[4033]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo_hi_1 = {regroupV0_hi_12[4045], regroupV0_hi_12[4041]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo_5 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo_hi_1, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi_lo_1 = {regroupV0_hi_12[4053], regroupV0_hi_12[4049]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi_hi_1 = {regroupV0_hi_12[4061], regroupV0_hi_12[4057]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi_5 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi_hi_1, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_9 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi_5, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo_lo_1 = {regroupV0_hi_12[4069], regroupV0_hi_12[4065]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo_hi_1 = {regroupV0_hi_12[4077], regroupV0_hi_12[4073]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo_5 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo_hi_1, regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi_lo_1 = {regroupV0_hi_12[4085], regroupV0_hi_12[4081]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi_hi_1 = {regroupV0_hi_12[4093], regroupV0_hi_12[4089]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi_5 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_9 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi_5, regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_hi_hi_12 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_9, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_9};
  wire [31:0]        regroupV0_hi_hi_hi_hi_hi_hi_12 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_12, regroupV0_hi_hi_hi_hi_hi_hi_lo_12};
  wire [63:0]        regroupV0_hi_hi_hi_hi_hi_12 = {regroupV0_hi_hi_hi_hi_hi_hi_12, regroupV0_hi_hi_hi_hi_hi_lo_12};
  wire [127:0]       regroupV0_hi_hi_hi_hi_12 = {regroupV0_hi_hi_hi_hi_hi_12, regroupV0_hi_hi_hi_hi_lo_12};
  wire [255:0]       regroupV0_hi_hi_hi_12 = {regroupV0_hi_hi_hi_hi_12, regroupV0_hi_hi_hi_lo_12};
  wire [511:0]       regroupV0_hi_hi_12 = {regroupV0_hi_hi_hi_12, regroupV0_hi_hi_lo_12};
  wire [1023:0]      regroupV0_hi_14 = {regroupV0_hi_hi_12, regroupV0_hi_lo_12};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo_lo_2 = {regroupV0_lo_12[6], regroupV0_lo_12[2]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo_hi_2 = {regroupV0_lo_12[14], regroupV0_lo_12[10]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo_6 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi_lo_2 = {regroupV0_lo_12[22], regroupV0_lo_12[18]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi_hi_2 = {regroupV0_lo_12[30], regroupV0_lo_12[26]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi_6 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi_hi_2, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_10 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi_6, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo_lo_2 = {regroupV0_lo_12[38], regroupV0_lo_12[34]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo_hi_2 = {regroupV0_lo_12[46], regroupV0_lo_12[42]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo_6 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo_hi_2, regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi_lo_2 = {regroupV0_lo_12[54], regroupV0_lo_12[50]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi_hi_2 = {regroupV0_lo_12[62], regroupV0_lo_12[58]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi_6 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi_hi_2, regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_10 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi_6, regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_lo_lo_13 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_10, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_10};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo_lo_2 = {regroupV0_lo_12[70], regroupV0_lo_12[66]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo_hi_2 = {regroupV0_lo_12[78], regroupV0_lo_12[74]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo_6 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi_lo_2 = {regroupV0_lo_12[86], regroupV0_lo_12[82]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi_hi_2 = {regroupV0_lo_12[94], regroupV0_lo_12[90]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi_6 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi_hi_2, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_10 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi_6, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo_lo_2 = {regroupV0_lo_12[102], regroupV0_lo_12[98]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo_hi_2 = {regroupV0_lo_12[110], regroupV0_lo_12[106]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo_6 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo_hi_2, regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi_lo_2 = {regroupV0_lo_12[118], regroupV0_lo_12[114]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi_hi_2 = {regroupV0_lo_12[126], regroupV0_lo_12[122]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi_6 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi_hi_2, regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_10 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi_6, regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_lo_hi_13 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_10, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_10};
  wire [31:0]        regroupV0_lo_lo_lo_lo_lo_lo_13 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_13, regroupV0_lo_lo_lo_lo_lo_lo_lo_13};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo_lo_2 = {regroupV0_lo_12[134], regroupV0_lo_12[130]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo_hi_2 = {regroupV0_lo_12[142], regroupV0_lo_12[138]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo_6 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi_lo_2 = {regroupV0_lo_12[150], regroupV0_lo_12[146]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi_hi_2 = {regroupV0_lo_12[158], regroupV0_lo_12[154]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi_6 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi_hi_2, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_10 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi_6, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo_lo_2 = {regroupV0_lo_12[166], regroupV0_lo_12[162]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo_hi_2 = {regroupV0_lo_12[174], regroupV0_lo_12[170]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo_6 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo_hi_2, regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi_lo_2 = {regroupV0_lo_12[182], regroupV0_lo_12[178]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi_hi_2 = {regroupV0_lo_12[190], regroupV0_lo_12[186]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi_6 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi_hi_2, regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_10 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi_6, regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_hi_lo_13 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_10, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_10};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo_lo_2 = {regroupV0_lo_12[198], regroupV0_lo_12[194]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo_hi_2 = {regroupV0_lo_12[206], regroupV0_lo_12[202]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo_6 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi_lo_2 = {regroupV0_lo_12[214], regroupV0_lo_12[210]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi_hi_2 = {regroupV0_lo_12[222], regroupV0_lo_12[218]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi_6 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi_hi_2, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_10 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi_6, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo_lo_2 = {regroupV0_lo_12[230], regroupV0_lo_12[226]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo_hi_2 = {regroupV0_lo_12[238], regroupV0_lo_12[234]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo_6 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo_hi_2, regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi_lo_2 = {regroupV0_lo_12[246], regroupV0_lo_12[242]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi_hi_2 = {regroupV0_lo_12[254], regroupV0_lo_12[250]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi_6 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi_hi_2, regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_10 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi_6, regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_hi_hi_13 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_10, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_10};
  wire [31:0]        regroupV0_lo_lo_lo_lo_lo_hi_13 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_13, regroupV0_lo_lo_lo_lo_lo_hi_lo_13};
  wire [63:0]        regroupV0_lo_lo_lo_lo_lo_13 = {regroupV0_lo_lo_lo_lo_lo_hi_13, regroupV0_lo_lo_lo_lo_lo_lo_13};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo_lo_2 = {regroupV0_lo_12[262], regroupV0_lo_12[258]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo_hi_2 = {regroupV0_lo_12[270], regroupV0_lo_12[266]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo_6 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi_lo_2 = {regroupV0_lo_12[278], regroupV0_lo_12[274]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi_hi_2 = {regroupV0_lo_12[286], regroupV0_lo_12[282]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi_6 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi_hi_2, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_10 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi_6, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo_lo_2 = {regroupV0_lo_12[294], regroupV0_lo_12[290]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo_hi_2 = {regroupV0_lo_12[302], regroupV0_lo_12[298]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo_6 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo_hi_2, regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi_lo_2 = {regroupV0_lo_12[310], regroupV0_lo_12[306]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi_hi_2 = {regroupV0_lo_12[318], regroupV0_lo_12[314]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi_6 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi_hi_2, regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_10 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi_6, regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_lo_lo_13 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_10, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_10};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo_lo_2 = {regroupV0_lo_12[326], regroupV0_lo_12[322]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo_hi_2 = {regroupV0_lo_12[334], regroupV0_lo_12[330]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo_6 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi_lo_2 = {regroupV0_lo_12[342], regroupV0_lo_12[338]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi_hi_2 = {regroupV0_lo_12[350], regroupV0_lo_12[346]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi_6 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi_hi_2, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_10 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi_6, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo_lo_2 = {regroupV0_lo_12[358], regroupV0_lo_12[354]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo_hi_2 = {regroupV0_lo_12[366], regroupV0_lo_12[362]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo_6 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo_hi_2, regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi_lo_2 = {regroupV0_lo_12[374], regroupV0_lo_12[370]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi_hi_2 = {regroupV0_lo_12[382], regroupV0_lo_12[378]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi_6 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi_hi_2, regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_10 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi_6, regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_lo_hi_13 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_10, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_10};
  wire [31:0]        regroupV0_lo_lo_lo_lo_hi_lo_13 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_13, regroupV0_lo_lo_lo_lo_hi_lo_lo_13};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo_lo_2 = {regroupV0_lo_12[390], regroupV0_lo_12[386]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo_hi_2 = {regroupV0_lo_12[398], regroupV0_lo_12[394]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo_6 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi_lo_2 = {regroupV0_lo_12[406], regroupV0_lo_12[402]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi_hi_2 = {regroupV0_lo_12[414], regroupV0_lo_12[410]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi_6 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi_hi_2, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_10 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi_6, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo_lo_2 = {regroupV0_lo_12[422], regroupV0_lo_12[418]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo_hi_2 = {regroupV0_lo_12[430], regroupV0_lo_12[426]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo_6 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo_hi_2, regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi_lo_2 = {regroupV0_lo_12[438], regroupV0_lo_12[434]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi_hi_2 = {regroupV0_lo_12[446], regroupV0_lo_12[442]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi_6 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi_hi_2, regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_10 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi_6, regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_hi_lo_13 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_10, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_10};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo_lo_2 = {regroupV0_lo_12[454], regroupV0_lo_12[450]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo_hi_2 = {regroupV0_lo_12[462], regroupV0_lo_12[458]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo_6 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi_lo_2 = {regroupV0_lo_12[470], regroupV0_lo_12[466]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi_hi_2 = {regroupV0_lo_12[478], regroupV0_lo_12[474]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi_6 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi_hi_2, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_10 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi_6, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo_lo_2 = {regroupV0_lo_12[486], regroupV0_lo_12[482]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo_hi_2 = {regroupV0_lo_12[494], regroupV0_lo_12[490]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo_6 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo_hi_2, regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi_lo_2 = {regroupV0_lo_12[502], regroupV0_lo_12[498]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi_hi_2 = {regroupV0_lo_12[510], regroupV0_lo_12[506]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi_6 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi_hi_2, regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_10 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi_6, regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_hi_hi_13 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_10, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_10};
  wire [31:0]        regroupV0_lo_lo_lo_lo_hi_hi_13 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_13, regroupV0_lo_lo_lo_lo_hi_hi_lo_13};
  wire [63:0]        regroupV0_lo_lo_lo_lo_hi_13 = {regroupV0_lo_lo_lo_lo_hi_hi_13, regroupV0_lo_lo_lo_lo_hi_lo_13};
  wire [127:0]       regroupV0_lo_lo_lo_lo_13 = {regroupV0_lo_lo_lo_lo_hi_13, regroupV0_lo_lo_lo_lo_lo_13};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo_lo_2 = {regroupV0_lo_12[518], regroupV0_lo_12[514]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo_hi_2 = {regroupV0_lo_12[526], regroupV0_lo_12[522]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo_6 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi_lo_2 = {regroupV0_lo_12[534], regroupV0_lo_12[530]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi_hi_2 = {regroupV0_lo_12[542], regroupV0_lo_12[538]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi_6 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi_hi_2, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_10 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi_6, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo_lo_2 = {regroupV0_lo_12[550], regroupV0_lo_12[546]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo_hi_2 = {regroupV0_lo_12[558], regroupV0_lo_12[554]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo_6 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo_hi_2, regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi_lo_2 = {regroupV0_lo_12[566], regroupV0_lo_12[562]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi_hi_2 = {regroupV0_lo_12[574], regroupV0_lo_12[570]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi_6 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi_hi_2, regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_10 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi_6, regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_lo_lo_13 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_10, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_10};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo_lo_2 = {regroupV0_lo_12[582], regroupV0_lo_12[578]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo_hi_2 = {regroupV0_lo_12[590], regroupV0_lo_12[586]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo_6 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo_hi_2, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi_lo_2 = {regroupV0_lo_12[598], regroupV0_lo_12[594]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi_hi_2 = {regroupV0_lo_12[606], regroupV0_lo_12[602]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi_6 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi_hi_2, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_10 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi_6, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo_lo_2 = {regroupV0_lo_12[614], regroupV0_lo_12[610]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo_hi_2 = {regroupV0_lo_12[622], regroupV0_lo_12[618]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo_6 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo_hi_2, regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi_lo_2 = {regroupV0_lo_12[630], regroupV0_lo_12[626]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi_hi_2 = {regroupV0_lo_12[638], regroupV0_lo_12[634]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi_6 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi_hi_2, regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_10 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi_6, regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_lo_hi_13 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_10, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_10};
  wire [31:0]        regroupV0_lo_lo_lo_hi_lo_lo_13 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_13, regroupV0_lo_lo_lo_hi_lo_lo_lo_13};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo_lo_2 = {regroupV0_lo_12[646], regroupV0_lo_12[642]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo_hi_2 = {regroupV0_lo_12[654], regroupV0_lo_12[650]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo_6 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi_lo_2 = {regroupV0_lo_12[662], regroupV0_lo_12[658]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi_hi_2 = {regroupV0_lo_12[670], regroupV0_lo_12[666]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi_6 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi_hi_2, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_10 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi_6, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo_lo_2 = {regroupV0_lo_12[678], regroupV0_lo_12[674]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo_hi_2 = {regroupV0_lo_12[686], regroupV0_lo_12[682]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo_6 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo_hi_2, regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi_lo_2 = {regroupV0_lo_12[694], regroupV0_lo_12[690]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi_hi_2 = {regroupV0_lo_12[702], regroupV0_lo_12[698]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi_6 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi_hi_2, regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_10 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi_6, regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_hi_lo_13 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_10, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_10};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo_lo_2 = {regroupV0_lo_12[710], regroupV0_lo_12[706]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo_hi_2 = {regroupV0_lo_12[718], regroupV0_lo_12[714]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo_6 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo_hi_2, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi_lo_2 = {regroupV0_lo_12[726], regroupV0_lo_12[722]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi_hi_2 = {regroupV0_lo_12[734], regroupV0_lo_12[730]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi_6 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi_hi_2, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_10 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi_6, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo_lo_2 = {regroupV0_lo_12[742], regroupV0_lo_12[738]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo_hi_2 = {regroupV0_lo_12[750], regroupV0_lo_12[746]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo_6 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo_hi_2, regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi_lo_2 = {regroupV0_lo_12[758], regroupV0_lo_12[754]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi_hi_2 = {regroupV0_lo_12[766], regroupV0_lo_12[762]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi_6 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi_hi_2, regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_10 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi_6, regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_hi_hi_13 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_10, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_10};
  wire [31:0]        regroupV0_lo_lo_lo_hi_lo_hi_13 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_13, regroupV0_lo_lo_lo_hi_lo_hi_lo_13};
  wire [63:0]        regroupV0_lo_lo_lo_hi_lo_13 = {regroupV0_lo_lo_lo_hi_lo_hi_13, regroupV0_lo_lo_lo_hi_lo_lo_13};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo_lo_2 = {regroupV0_lo_12[774], regroupV0_lo_12[770]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo_hi_2 = {regroupV0_lo_12[782], regroupV0_lo_12[778]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo_6 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi_lo_2 = {regroupV0_lo_12[790], regroupV0_lo_12[786]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi_hi_2 = {regroupV0_lo_12[798], regroupV0_lo_12[794]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi_6 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi_hi_2, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_10 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi_6, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo_lo_2 = {regroupV0_lo_12[806], regroupV0_lo_12[802]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo_hi_2 = {regroupV0_lo_12[814], regroupV0_lo_12[810]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo_6 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo_hi_2, regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi_lo_2 = {regroupV0_lo_12[822], regroupV0_lo_12[818]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi_hi_2 = {regroupV0_lo_12[830], regroupV0_lo_12[826]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi_6 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi_hi_2, regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_10 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi_6, regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_lo_lo_13 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_10, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_10};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo_lo_2 = {regroupV0_lo_12[838], regroupV0_lo_12[834]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo_hi_2 = {regroupV0_lo_12[846], regroupV0_lo_12[842]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo_6 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo_hi_2, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi_lo_2 = {regroupV0_lo_12[854], regroupV0_lo_12[850]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi_hi_2 = {regroupV0_lo_12[862], regroupV0_lo_12[858]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi_6 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi_hi_2, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_10 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi_6, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo_lo_2 = {regroupV0_lo_12[870], regroupV0_lo_12[866]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo_hi_2 = {regroupV0_lo_12[878], regroupV0_lo_12[874]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo_6 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo_hi_2, regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi_lo_2 = {regroupV0_lo_12[886], regroupV0_lo_12[882]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi_hi_2 = {regroupV0_lo_12[894], regroupV0_lo_12[890]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi_6 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi_hi_2, regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_10 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi_6, regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_lo_hi_13 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_10, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_10};
  wire [31:0]        regroupV0_lo_lo_lo_hi_hi_lo_13 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_13, regroupV0_lo_lo_lo_hi_hi_lo_lo_13};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo_lo_2 = {regroupV0_lo_12[902], regroupV0_lo_12[898]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo_hi_2 = {regroupV0_lo_12[910], regroupV0_lo_12[906]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo_6 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi_lo_2 = {regroupV0_lo_12[918], regroupV0_lo_12[914]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi_hi_2 = {regroupV0_lo_12[926], regroupV0_lo_12[922]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi_6 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi_hi_2, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_10 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi_6, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo_lo_2 = {regroupV0_lo_12[934], regroupV0_lo_12[930]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo_hi_2 = {regroupV0_lo_12[942], regroupV0_lo_12[938]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo_6 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo_hi_2, regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi_lo_2 = {regroupV0_lo_12[950], regroupV0_lo_12[946]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi_hi_2 = {regroupV0_lo_12[958], regroupV0_lo_12[954]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi_6 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi_hi_2, regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_10 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi_6, regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_hi_lo_13 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_10, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_10};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo_lo_2 = {regroupV0_lo_12[966], regroupV0_lo_12[962]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo_hi_2 = {regroupV0_lo_12[974], regroupV0_lo_12[970]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo_6 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo_hi_2, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi_lo_2 = {regroupV0_lo_12[982], regroupV0_lo_12[978]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi_hi_2 = {regroupV0_lo_12[990], regroupV0_lo_12[986]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi_6 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi_hi_2, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_10 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi_6, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo_lo_2 = {regroupV0_lo_12[998], regroupV0_lo_12[994]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo_hi_2 = {regroupV0_lo_12[1006], regroupV0_lo_12[1002]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo_6 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo_hi_2, regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi_lo_2 = {regroupV0_lo_12[1014], regroupV0_lo_12[1010]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi_hi_2 = {regroupV0_lo_12[1022], regroupV0_lo_12[1018]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi_6 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi_hi_2, regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_10 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi_6, regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_hi_hi_13 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_10, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_10};
  wire [31:0]        regroupV0_lo_lo_lo_hi_hi_hi_13 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_13, regroupV0_lo_lo_lo_hi_hi_hi_lo_13};
  wire [63:0]        regroupV0_lo_lo_lo_hi_hi_13 = {regroupV0_lo_lo_lo_hi_hi_hi_13, regroupV0_lo_lo_lo_hi_hi_lo_13};
  wire [127:0]       regroupV0_lo_lo_lo_hi_13 = {regroupV0_lo_lo_lo_hi_hi_13, regroupV0_lo_lo_lo_hi_lo_13};
  wire [255:0]       regroupV0_lo_lo_lo_13 = {regroupV0_lo_lo_lo_hi_13, regroupV0_lo_lo_lo_lo_13};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo_lo_2 = {regroupV0_lo_12[1030], regroupV0_lo_12[1026]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo_hi_2 = {regroupV0_lo_12[1038], regroupV0_lo_12[1034]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo_6 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo_hi_2, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi_lo_2 = {regroupV0_lo_12[1046], regroupV0_lo_12[1042]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi_hi_2 = {regroupV0_lo_12[1054], regroupV0_lo_12[1050]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi_6 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi_hi_2, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_10 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi_6, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo_lo_2 = {regroupV0_lo_12[1062], regroupV0_lo_12[1058]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo_hi_2 = {regroupV0_lo_12[1070], regroupV0_lo_12[1066]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo_6 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo_hi_2, regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi_lo_2 = {regroupV0_lo_12[1078], regroupV0_lo_12[1074]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi_hi_2 = {regroupV0_lo_12[1086], regroupV0_lo_12[1082]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi_6 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi_hi_2, regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_10 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi_6, regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_lo_lo_13 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_10, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_10};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo_lo_2 = {regroupV0_lo_12[1094], regroupV0_lo_12[1090]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo_hi_2 = {regroupV0_lo_12[1102], regroupV0_lo_12[1098]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo_6 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo_hi_2, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi_lo_2 = {regroupV0_lo_12[1110], regroupV0_lo_12[1106]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi_hi_2 = {regroupV0_lo_12[1118], regroupV0_lo_12[1114]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi_6 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi_hi_2, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_10 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi_6, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo_lo_2 = {regroupV0_lo_12[1126], regroupV0_lo_12[1122]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo_hi_2 = {regroupV0_lo_12[1134], regroupV0_lo_12[1130]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo_6 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo_hi_2, regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi_lo_2 = {regroupV0_lo_12[1142], regroupV0_lo_12[1138]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi_hi_2 = {regroupV0_lo_12[1150], regroupV0_lo_12[1146]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi_6 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi_hi_2, regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_10 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi_6, regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_lo_hi_13 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_10, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_10};
  wire [31:0]        regroupV0_lo_lo_hi_lo_lo_lo_13 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_13, regroupV0_lo_lo_hi_lo_lo_lo_lo_13};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo_lo_2 = {regroupV0_lo_12[1158], regroupV0_lo_12[1154]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo_hi_2 = {regroupV0_lo_12[1166], regroupV0_lo_12[1162]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo_6 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo_hi_2, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi_lo_2 = {regroupV0_lo_12[1174], regroupV0_lo_12[1170]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi_hi_2 = {regroupV0_lo_12[1182], regroupV0_lo_12[1178]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi_6 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi_hi_2, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_10 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi_6, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo_lo_2 = {regroupV0_lo_12[1190], regroupV0_lo_12[1186]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo_hi_2 = {regroupV0_lo_12[1198], regroupV0_lo_12[1194]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo_6 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo_hi_2, regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi_lo_2 = {regroupV0_lo_12[1206], regroupV0_lo_12[1202]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi_hi_2 = {regroupV0_lo_12[1214], regroupV0_lo_12[1210]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi_6 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi_hi_2, regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_10 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi_6, regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_hi_lo_13 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_10, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_10};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo_lo_2 = {regroupV0_lo_12[1222], regroupV0_lo_12[1218]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo_hi_2 = {regroupV0_lo_12[1230], regroupV0_lo_12[1226]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo_6 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo_hi_2, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi_lo_2 = {regroupV0_lo_12[1238], regroupV0_lo_12[1234]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi_hi_2 = {regroupV0_lo_12[1246], regroupV0_lo_12[1242]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi_6 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi_hi_2, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_10 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi_6, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo_lo_2 = {regroupV0_lo_12[1254], regroupV0_lo_12[1250]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo_hi_2 = {regroupV0_lo_12[1262], regroupV0_lo_12[1258]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo_6 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo_hi_2, regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi_lo_2 = {regroupV0_lo_12[1270], regroupV0_lo_12[1266]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi_hi_2 = {regroupV0_lo_12[1278], regroupV0_lo_12[1274]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi_6 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi_hi_2, regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_10 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi_6, regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_hi_hi_13 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_10, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_10};
  wire [31:0]        regroupV0_lo_lo_hi_lo_lo_hi_13 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_13, regroupV0_lo_lo_hi_lo_lo_hi_lo_13};
  wire [63:0]        regroupV0_lo_lo_hi_lo_lo_13 = {regroupV0_lo_lo_hi_lo_lo_hi_13, regroupV0_lo_lo_hi_lo_lo_lo_13};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo_lo_2 = {regroupV0_lo_12[1286], regroupV0_lo_12[1282]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo_hi_2 = {regroupV0_lo_12[1294], regroupV0_lo_12[1290]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo_6 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo_hi_2, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi_lo_2 = {regroupV0_lo_12[1302], regroupV0_lo_12[1298]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi_hi_2 = {regroupV0_lo_12[1310], regroupV0_lo_12[1306]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi_6 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi_hi_2, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_10 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi_6, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo_lo_2 = {regroupV0_lo_12[1318], regroupV0_lo_12[1314]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo_hi_2 = {regroupV0_lo_12[1326], regroupV0_lo_12[1322]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo_6 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo_hi_2, regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi_lo_2 = {regroupV0_lo_12[1334], regroupV0_lo_12[1330]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi_hi_2 = {regroupV0_lo_12[1342], regroupV0_lo_12[1338]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi_6 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi_hi_2, regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_10 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi_6, regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_lo_lo_13 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_10, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_10};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo_lo_2 = {regroupV0_lo_12[1350], regroupV0_lo_12[1346]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo_hi_2 = {regroupV0_lo_12[1358], regroupV0_lo_12[1354]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo_6 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo_hi_2, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi_lo_2 = {regroupV0_lo_12[1366], regroupV0_lo_12[1362]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi_hi_2 = {regroupV0_lo_12[1374], regroupV0_lo_12[1370]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi_6 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi_hi_2, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_10 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi_6, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo_lo_2 = {regroupV0_lo_12[1382], regroupV0_lo_12[1378]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo_hi_2 = {regroupV0_lo_12[1390], regroupV0_lo_12[1386]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo_6 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo_hi_2, regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi_lo_2 = {regroupV0_lo_12[1398], regroupV0_lo_12[1394]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi_hi_2 = {regroupV0_lo_12[1406], regroupV0_lo_12[1402]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi_6 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi_hi_2, regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_10 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi_6, regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_lo_hi_13 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_10, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_10};
  wire [31:0]        regroupV0_lo_lo_hi_lo_hi_lo_13 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_13, regroupV0_lo_lo_hi_lo_hi_lo_lo_13};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo_lo_2 = {regroupV0_lo_12[1414], regroupV0_lo_12[1410]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo_hi_2 = {regroupV0_lo_12[1422], regroupV0_lo_12[1418]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo_6 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo_hi_2, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi_lo_2 = {regroupV0_lo_12[1430], regroupV0_lo_12[1426]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi_hi_2 = {regroupV0_lo_12[1438], regroupV0_lo_12[1434]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi_6 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi_hi_2, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_10 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi_6, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo_lo_2 = {regroupV0_lo_12[1446], regroupV0_lo_12[1442]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo_hi_2 = {regroupV0_lo_12[1454], regroupV0_lo_12[1450]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo_6 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo_hi_2, regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi_lo_2 = {regroupV0_lo_12[1462], regroupV0_lo_12[1458]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi_hi_2 = {regroupV0_lo_12[1470], regroupV0_lo_12[1466]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi_6 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi_hi_2, regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_10 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi_6, regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_hi_lo_13 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_10, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_10};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo_lo_2 = {regroupV0_lo_12[1478], regroupV0_lo_12[1474]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo_hi_2 = {regroupV0_lo_12[1486], regroupV0_lo_12[1482]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo_6 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo_hi_2, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi_lo_2 = {regroupV0_lo_12[1494], regroupV0_lo_12[1490]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi_hi_2 = {regroupV0_lo_12[1502], regroupV0_lo_12[1498]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi_6 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi_hi_2, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_10 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi_6, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo_lo_2 = {regroupV0_lo_12[1510], regroupV0_lo_12[1506]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo_hi_2 = {regroupV0_lo_12[1518], regroupV0_lo_12[1514]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo_6 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo_hi_2, regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi_lo_2 = {regroupV0_lo_12[1526], regroupV0_lo_12[1522]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi_hi_2 = {regroupV0_lo_12[1534], regroupV0_lo_12[1530]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi_6 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi_hi_2, regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_10 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi_6, regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_hi_hi_13 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_10, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_10};
  wire [31:0]        regroupV0_lo_lo_hi_lo_hi_hi_13 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_13, regroupV0_lo_lo_hi_lo_hi_hi_lo_13};
  wire [63:0]        regroupV0_lo_lo_hi_lo_hi_13 = {regroupV0_lo_lo_hi_lo_hi_hi_13, regroupV0_lo_lo_hi_lo_hi_lo_13};
  wire [127:0]       regroupV0_lo_lo_hi_lo_13 = {regroupV0_lo_lo_hi_lo_hi_13, regroupV0_lo_lo_hi_lo_lo_13};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo_lo_2 = {regroupV0_lo_12[1542], regroupV0_lo_12[1538]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo_hi_2 = {regroupV0_lo_12[1550], regroupV0_lo_12[1546]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo_6 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo_hi_2, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi_lo_2 = {regroupV0_lo_12[1558], regroupV0_lo_12[1554]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi_hi_2 = {regroupV0_lo_12[1566], regroupV0_lo_12[1562]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi_6 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi_hi_2, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_10 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi_6, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo_lo_2 = {regroupV0_lo_12[1574], regroupV0_lo_12[1570]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo_hi_2 = {regroupV0_lo_12[1582], regroupV0_lo_12[1578]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo_6 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo_hi_2, regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi_lo_2 = {regroupV0_lo_12[1590], regroupV0_lo_12[1586]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi_hi_2 = {regroupV0_lo_12[1598], regroupV0_lo_12[1594]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi_6 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi_hi_2, regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_10 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi_6, regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_lo_lo_13 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_10, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_10};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo_lo_2 = {regroupV0_lo_12[1606], regroupV0_lo_12[1602]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo_hi_2 = {regroupV0_lo_12[1614], regroupV0_lo_12[1610]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo_6 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo_hi_2, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi_lo_2 = {regroupV0_lo_12[1622], regroupV0_lo_12[1618]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi_hi_2 = {regroupV0_lo_12[1630], regroupV0_lo_12[1626]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi_6 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi_hi_2, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_10 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi_6, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo_lo_2 = {regroupV0_lo_12[1638], regroupV0_lo_12[1634]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo_hi_2 = {regroupV0_lo_12[1646], regroupV0_lo_12[1642]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo_6 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo_hi_2, regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi_lo_2 = {regroupV0_lo_12[1654], regroupV0_lo_12[1650]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi_hi_2 = {regroupV0_lo_12[1662], regroupV0_lo_12[1658]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi_6 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi_hi_2, regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_10 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi_6, regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_lo_hi_13 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_10, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_10};
  wire [31:0]        regroupV0_lo_lo_hi_hi_lo_lo_13 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_13, regroupV0_lo_lo_hi_hi_lo_lo_lo_13};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo_lo_2 = {regroupV0_lo_12[1670], regroupV0_lo_12[1666]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo_hi_2 = {regroupV0_lo_12[1678], regroupV0_lo_12[1674]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo_6 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo_hi_2, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi_lo_2 = {regroupV0_lo_12[1686], regroupV0_lo_12[1682]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi_hi_2 = {regroupV0_lo_12[1694], regroupV0_lo_12[1690]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi_6 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi_hi_2, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_10 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi_6, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo_lo_2 = {regroupV0_lo_12[1702], regroupV0_lo_12[1698]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo_hi_2 = {regroupV0_lo_12[1710], regroupV0_lo_12[1706]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo_6 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo_hi_2, regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi_lo_2 = {regroupV0_lo_12[1718], regroupV0_lo_12[1714]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi_hi_2 = {regroupV0_lo_12[1726], regroupV0_lo_12[1722]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi_6 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi_hi_2, regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_10 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi_6, regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_hi_lo_13 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_10, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_10};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo_lo_2 = {regroupV0_lo_12[1734], regroupV0_lo_12[1730]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo_hi_2 = {regroupV0_lo_12[1742], regroupV0_lo_12[1738]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo_6 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo_hi_2, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi_lo_2 = {regroupV0_lo_12[1750], regroupV0_lo_12[1746]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi_hi_2 = {regroupV0_lo_12[1758], regroupV0_lo_12[1754]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi_6 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi_hi_2, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_10 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi_6, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo_lo_2 = {regroupV0_lo_12[1766], regroupV0_lo_12[1762]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo_hi_2 = {regroupV0_lo_12[1774], regroupV0_lo_12[1770]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo_6 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo_hi_2, regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi_lo_2 = {regroupV0_lo_12[1782], regroupV0_lo_12[1778]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi_hi_2 = {regroupV0_lo_12[1790], regroupV0_lo_12[1786]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi_6 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi_hi_2, regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_10 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi_6, regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_hi_hi_13 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_10, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_10};
  wire [31:0]        regroupV0_lo_lo_hi_hi_lo_hi_13 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_13, regroupV0_lo_lo_hi_hi_lo_hi_lo_13};
  wire [63:0]        regroupV0_lo_lo_hi_hi_lo_13 = {regroupV0_lo_lo_hi_hi_lo_hi_13, regroupV0_lo_lo_hi_hi_lo_lo_13};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo_lo_2 = {regroupV0_lo_12[1798], regroupV0_lo_12[1794]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo_hi_2 = {regroupV0_lo_12[1806], regroupV0_lo_12[1802]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo_6 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo_hi_2, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi_lo_2 = {regroupV0_lo_12[1814], regroupV0_lo_12[1810]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi_hi_2 = {regroupV0_lo_12[1822], regroupV0_lo_12[1818]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi_6 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi_hi_2, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_10 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi_6, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo_lo_2 = {regroupV0_lo_12[1830], regroupV0_lo_12[1826]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo_hi_2 = {regroupV0_lo_12[1838], regroupV0_lo_12[1834]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo_6 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo_hi_2, regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi_lo_2 = {regroupV0_lo_12[1846], regroupV0_lo_12[1842]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi_hi_2 = {regroupV0_lo_12[1854], regroupV0_lo_12[1850]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi_6 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi_hi_2, regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_10 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi_6, regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_lo_lo_13 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_10, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_10};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo_lo_2 = {regroupV0_lo_12[1862], regroupV0_lo_12[1858]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo_hi_2 = {regroupV0_lo_12[1870], regroupV0_lo_12[1866]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo_6 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo_hi_2, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi_lo_2 = {regroupV0_lo_12[1878], regroupV0_lo_12[1874]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi_hi_2 = {regroupV0_lo_12[1886], regroupV0_lo_12[1882]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi_6 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi_hi_2, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_10 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi_6, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo_lo_2 = {regroupV0_lo_12[1894], regroupV0_lo_12[1890]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo_hi_2 = {regroupV0_lo_12[1902], regroupV0_lo_12[1898]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo_6 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo_hi_2, regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi_lo_2 = {regroupV0_lo_12[1910], regroupV0_lo_12[1906]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi_hi_2 = {regroupV0_lo_12[1918], regroupV0_lo_12[1914]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi_6 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi_hi_2, regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_10 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi_6, regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_lo_hi_13 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_10, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_10};
  wire [31:0]        regroupV0_lo_lo_hi_hi_hi_lo_13 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_13, regroupV0_lo_lo_hi_hi_hi_lo_lo_13};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo_lo_2 = {regroupV0_lo_12[1926], regroupV0_lo_12[1922]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo_hi_2 = {regroupV0_lo_12[1934], regroupV0_lo_12[1930]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo_6 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo_hi_2, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi_lo_2 = {regroupV0_lo_12[1942], regroupV0_lo_12[1938]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi_hi_2 = {regroupV0_lo_12[1950], regroupV0_lo_12[1946]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi_6 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi_hi_2, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_10 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi_6, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo_lo_2 = {regroupV0_lo_12[1958], regroupV0_lo_12[1954]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo_hi_2 = {regroupV0_lo_12[1966], regroupV0_lo_12[1962]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo_6 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo_hi_2, regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi_lo_2 = {regroupV0_lo_12[1974], regroupV0_lo_12[1970]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi_hi_2 = {regroupV0_lo_12[1982], regroupV0_lo_12[1978]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi_6 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi_hi_2, regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_10 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi_6, regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_hi_lo_13 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_10, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_10};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo_lo_2 = {regroupV0_lo_12[1990], regroupV0_lo_12[1986]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo_hi_2 = {regroupV0_lo_12[1998], regroupV0_lo_12[1994]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo_6 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo_hi_2, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi_lo_2 = {regroupV0_lo_12[2006], regroupV0_lo_12[2002]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi_hi_2 = {regroupV0_lo_12[2014], regroupV0_lo_12[2010]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi_6 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi_hi_2, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_10 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi_6, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo_lo_2 = {regroupV0_lo_12[2022], regroupV0_lo_12[2018]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo_hi_2 = {regroupV0_lo_12[2030], regroupV0_lo_12[2026]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo_6 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo_hi_2, regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi_lo_2 = {regroupV0_lo_12[2038], regroupV0_lo_12[2034]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi_hi_2 = {regroupV0_lo_12[2046], regroupV0_lo_12[2042]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi_6 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi_hi_2, regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_10 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi_6, regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_hi_hi_13 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_10, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_10};
  wire [31:0]        regroupV0_lo_lo_hi_hi_hi_hi_13 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_13, regroupV0_lo_lo_hi_hi_hi_hi_lo_13};
  wire [63:0]        regroupV0_lo_lo_hi_hi_hi_13 = {regroupV0_lo_lo_hi_hi_hi_hi_13, regroupV0_lo_lo_hi_hi_hi_lo_13};
  wire [127:0]       regroupV0_lo_lo_hi_hi_13 = {regroupV0_lo_lo_hi_hi_hi_13, regroupV0_lo_lo_hi_hi_lo_13};
  wire [255:0]       regroupV0_lo_lo_hi_13 = {regroupV0_lo_lo_hi_hi_13, regroupV0_lo_lo_hi_lo_13};
  wire [511:0]       regroupV0_lo_lo_13 = {regroupV0_lo_lo_hi_13, regroupV0_lo_lo_lo_13};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo_lo_2 = {regroupV0_lo_12[2054], regroupV0_lo_12[2050]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo_hi_2 = {regroupV0_lo_12[2062], regroupV0_lo_12[2058]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo_6 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo_hi_2, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi_lo_2 = {regroupV0_lo_12[2070], regroupV0_lo_12[2066]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi_hi_2 = {regroupV0_lo_12[2078], regroupV0_lo_12[2074]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi_6 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi_hi_2, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_10 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi_6, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo_lo_2 = {regroupV0_lo_12[2086], regroupV0_lo_12[2082]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo_hi_2 = {regroupV0_lo_12[2094], regroupV0_lo_12[2090]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo_6 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo_hi_2, regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi_lo_2 = {regroupV0_lo_12[2102], regroupV0_lo_12[2098]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi_hi_2 = {regroupV0_lo_12[2110], regroupV0_lo_12[2106]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi_6 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi_hi_2, regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_10 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi_6, regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_lo_lo_13 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_10, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_10};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo_lo_2 = {regroupV0_lo_12[2118], regroupV0_lo_12[2114]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo_hi_2 = {regroupV0_lo_12[2126], regroupV0_lo_12[2122]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo_6 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo_hi_2, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi_lo_2 = {regroupV0_lo_12[2134], regroupV0_lo_12[2130]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi_hi_2 = {regroupV0_lo_12[2142], regroupV0_lo_12[2138]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi_6 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi_hi_2, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_10 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi_6, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo_lo_2 = {regroupV0_lo_12[2150], regroupV0_lo_12[2146]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo_hi_2 = {regroupV0_lo_12[2158], regroupV0_lo_12[2154]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo_6 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo_hi_2, regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi_lo_2 = {regroupV0_lo_12[2166], regroupV0_lo_12[2162]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi_hi_2 = {regroupV0_lo_12[2174], regroupV0_lo_12[2170]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi_6 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi_hi_2, regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_10 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi_6, regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_lo_hi_13 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_10, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_10};
  wire [31:0]        regroupV0_lo_hi_lo_lo_lo_lo_13 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_13, regroupV0_lo_hi_lo_lo_lo_lo_lo_13};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo_lo_2 = {regroupV0_lo_12[2182], regroupV0_lo_12[2178]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo_hi_2 = {regroupV0_lo_12[2190], regroupV0_lo_12[2186]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo_6 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo_hi_2, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi_lo_2 = {regroupV0_lo_12[2198], regroupV0_lo_12[2194]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi_hi_2 = {regroupV0_lo_12[2206], regroupV0_lo_12[2202]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi_6 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi_hi_2, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_10 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi_6, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo_lo_2 = {regroupV0_lo_12[2214], regroupV0_lo_12[2210]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo_hi_2 = {regroupV0_lo_12[2222], regroupV0_lo_12[2218]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo_6 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo_hi_2, regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi_lo_2 = {regroupV0_lo_12[2230], regroupV0_lo_12[2226]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi_hi_2 = {regroupV0_lo_12[2238], regroupV0_lo_12[2234]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi_6 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi_hi_2, regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_10 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi_6, regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_hi_lo_13 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_10, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_10};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo_lo_2 = {regroupV0_lo_12[2246], regroupV0_lo_12[2242]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo_hi_2 = {regroupV0_lo_12[2254], regroupV0_lo_12[2250]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo_6 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo_hi_2, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi_lo_2 = {regroupV0_lo_12[2262], regroupV0_lo_12[2258]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi_hi_2 = {regroupV0_lo_12[2270], regroupV0_lo_12[2266]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi_6 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi_hi_2, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_10 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi_6, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo_lo_2 = {regroupV0_lo_12[2278], regroupV0_lo_12[2274]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo_hi_2 = {regroupV0_lo_12[2286], regroupV0_lo_12[2282]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo_6 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo_hi_2, regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi_lo_2 = {regroupV0_lo_12[2294], regroupV0_lo_12[2290]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi_hi_2 = {regroupV0_lo_12[2302], regroupV0_lo_12[2298]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi_6 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi_hi_2, regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_10 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi_6, regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_hi_hi_13 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_10, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_10};
  wire [31:0]        regroupV0_lo_hi_lo_lo_lo_hi_13 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_13, regroupV0_lo_hi_lo_lo_lo_hi_lo_13};
  wire [63:0]        regroupV0_lo_hi_lo_lo_lo_13 = {regroupV0_lo_hi_lo_lo_lo_hi_13, regroupV0_lo_hi_lo_lo_lo_lo_13};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo_lo_2 = {regroupV0_lo_12[2310], regroupV0_lo_12[2306]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo_hi_2 = {regroupV0_lo_12[2318], regroupV0_lo_12[2314]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo_6 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo_hi_2, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi_lo_2 = {regroupV0_lo_12[2326], regroupV0_lo_12[2322]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi_hi_2 = {regroupV0_lo_12[2334], regroupV0_lo_12[2330]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi_6 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi_hi_2, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_10 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi_6, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo_lo_2 = {regroupV0_lo_12[2342], regroupV0_lo_12[2338]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo_hi_2 = {regroupV0_lo_12[2350], regroupV0_lo_12[2346]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo_6 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo_hi_2, regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi_lo_2 = {regroupV0_lo_12[2358], regroupV0_lo_12[2354]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi_hi_2 = {regroupV0_lo_12[2366], regroupV0_lo_12[2362]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi_6 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi_hi_2, regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_10 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi_6, regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_lo_lo_13 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_10, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_10};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo_lo_2 = {regroupV0_lo_12[2374], regroupV0_lo_12[2370]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo_hi_2 = {regroupV0_lo_12[2382], regroupV0_lo_12[2378]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo_6 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo_hi_2, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi_lo_2 = {regroupV0_lo_12[2390], regroupV0_lo_12[2386]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi_hi_2 = {regroupV0_lo_12[2398], regroupV0_lo_12[2394]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi_6 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi_hi_2, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_10 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi_6, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo_lo_2 = {regroupV0_lo_12[2406], regroupV0_lo_12[2402]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo_hi_2 = {regroupV0_lo_12[2414], regroupV0_lo_12[2410]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo_6 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo_hi_2, regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi_lo_2 = {regroupV0_lo_12[2422], regroupV0_lo_12[2418]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi_hi_2 = {regroupV0_lo_12[2430], regroupV0_lo_12[2426]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi_6 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi_hi_2, regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_10 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi_6, regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_lo_hi_13 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_10, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_10};
  wire [31:0]        regroupV0_lo_hi_lo_lo_hi_lo_13 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_13, regroupV0_lo_hi_lo_lo_hi_lo_lo_13};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo_lo_2 = {regroupV0_lo_12[2438], regroupV0_lo_12[2434]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo_hi_2 = {regroupV0_lo_12[2446], regroupV0_lo_12[2442]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo_6 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo_hi_2, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi_lo_2 = {regroupV0_lo_12[2454], regroupV0_lo_12[2450]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi_hi_2 = {regroupV0_lo_12[2462], regroupV0_lo_12[2458]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi_6 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi_hi_2, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_10 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi_6, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo_lo_2 = {regroupV0_lo_12[2470], regroupV0_lo_12[2466]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo_hi_2 = {regroupV0_lo_12[2478], regroupV0_lo_12[2474]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo_6 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo_hi_2, regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi_lo_2 = {regroupV0_lo_12[2486], regroupV0_lo_12[2482]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi_hi_2 = {regroupV0_lo_12[2494], regroupV0_lo_12[2490]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi_6 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi_hi_2, regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_10 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi_6, regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_hi_lo_13 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_10, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_10};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo_lo_2 = {regroupV0_lo_12[2502], regroupV0_lo_12[2498]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo_hi_2 = {regroupV0_lo_12[2510], regroupV0_lo_12[2506]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo_6 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo_hi_2, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi_lo_2 = {regroupV0_lo_12[2518], regroupV0_lo_12[2514]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi_hi_2 = {regroupV0_lo_12[2526], regroupV0_lo_12[2522]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi_6 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi_hi_2, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_10 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi_6, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo_lo_2 = {regroupV0_lo_12[2534], regroupV0_lo_12[2530]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo_hi_2 = {regroupV0_lo_12[2542], regroupV0_lo_12[2538]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo_6 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo_hi_2, regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi_lo_2 = {regroupV0_lo_12[2550], regroupV0_lo_12[2546]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi_hi_2 = {regroupV0_lo_12[2558], regroupV0_lo_12[2554]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi_6 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi_hi_2, regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_10 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi_6, regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_hi_hi_13 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_10, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_10};
  wire [31:0]        regroupV0_lo_hi_lo_lo_hi_hi_13 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_13, regroupV0_lo_hi_lo_lo_hi_hi_lo_13};
  wire [63:0]        regroupV0_lo_hi_lo_lo_hi_13 = {regroupV0_lo_hi_lo_lo_hi_hi_13, regroupV0_lo_hi_lo_lo_hi_lo_13};
  wire [127:0]       regroupV0_lo_hi_lo_lo_13 = {regroupV0_lo_hi_lo_lo_hi_13, regroupV0_lo_hi_lo_lo_lo_13};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo_lo_2 = {regroupV0_lo_12[2566], regroupV0_lo_12[2562]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo_hi_2 = {regroupV0_lo_12[2574], regroupV0_lo_12[2570]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo_6 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo_hi_2, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi_lo_2 = {regroupV0_lo_12[2582], regroupV0_lo_12[2578]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi_hi_2 = {regroupV0_lo_12[2590], regroupV0_lo_12[2586]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi_6 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi_hi_2, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_10 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi_6, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo_lo_2 = {regroupV0_lo_12[2598], regroupV0_lo_12[2594]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo_hi_2 = {regroupV0_lo_12[2606], regroupV0_lo_12[2602]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo_6 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo_hi_2, regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi_lo_2 = {regroupV0_lo_12[2614], regroupV0_lo_12[2610]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi_hi_2 = {regroupV0_lo_12[2622], regroupV0_lo_12[2618]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi_6 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi_hi_2, regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_10 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi_6, regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_lo_lo_13 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_10, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_10};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo_lo_2 = {regroupV0_lo_12[2630], regroupV0_lo_12[2626]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo_hi_2 = {regroupV0_lo_12[2638], regroupV0_lo_12[2634]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo_6 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo_hi_2, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi_lo_2 = {regroupV0_lo_12[2646], regroupV0_lo_12[2642]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi_hi_2 = {regroupV0_lo_12[2654], regroupV0_lo_12[2650]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi_6 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi_hi_2, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_10 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi_6, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo_lo_2 = {regroupV0_lo_12[2662], regroupV0_lo_12[2658]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo_hi_2 = {regroupV0_lo_12[2670], regroupV0_lo_12[2666]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo_6 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo_hi_2, regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi_lo_2 = {regroupV0_lo_12[2678], regroupV0_lo_12[2674]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi_hi_2 = {regroupV0_lo_12[2686], regroupV0_lo_12[2682]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi_6 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi_hi_2, regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_10 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi_6, regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_lo_hi_13 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_10, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_10};
  wire [31:0]        regroupV0_lo_hi_lo_hi_lo_lo_13 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_13, regroupV0_lo_hi_lo_hi_lo_lo_lo_13};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo_lo_2 = {regroupV0_lo_12[2694], regroupV0_lo_12[2690]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo_hi_2 = {regroupV0_lo_12[2702], regroupV0_lo_12[2698]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo_6 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo_hi_2, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi_lo_2 = {regroupV0_lo_12[2710], regroupV0_lo_12[2706]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi_hi_2 = {regroupV0_lo_12[2718], regroupV0_lo_12[2714]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi_6 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi_hi_2, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_10 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi_6, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo_lo_2 = {regroupV0_lo_12[2726], regroupV0_lo_12[2722]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo_hi_2 = {regroupV0_lo_12[2734], regroupV0_lo_12[2730]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo_6 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo_hi_2, regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi_lo_2 = {regroupV0_lo_12[2742], regroupV0_lo_12[2738]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi_hi_2 = {regroupV0_lo_12[2750], regroupV0_lo_12[2746]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi_6 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi_hi_2, regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_10 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi_6, regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_hi_lo_13 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_10, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_10};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo_lo_2 = {regroupV0_lo_12[2758], regroupV0_lo_12[2754]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo_hi_2 = {regroupV0_lo_12[2766], regroupV0_lo_12[2762]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo_6 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo_hi_2, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi_lo_2 = {regroupV0_lo_12[2774], regroupV0_lo_12[2770]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi_hi_2 = {regroupV0_lo_12[2782], regroupV0_lo_12[2778]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi_6 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi_hi_2, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_10 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi_6, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo_lo_2 = {regroupV0_lo_12[2790], regroupV0_lo_12[2786]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo_hi_2 = {regroupV0_lo_12[2798], regroupV0_lo_12[2794]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo_6 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo_hi_2, regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi_lo_2 = {regroupV0_lo_12[2806], regroupV0_lo_12[2802]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi_hi_2 = {regroupV0_lo_12[2814], regroupV0_lo_12[2810]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi_6 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi_hi_2, regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_10 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi_6, regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_hi_hi_13 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_10, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_10};
  wire [31:0]        regroupV0_lo_hi_lo_hi_lo_hi_13 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_13, regroupV0_lo_hi_lo_hi_lo_hi_lo_13};
  wire [63:0]        regroupV0_lo_hi_lo_hi_lo_13 = {regroupV0_lo_hi_lo_hi_lo_hi_13, regroupV0_lo_hi_lo_hi_lo_lo_13};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo_lo_2 = {regroupV0_lo_12[2822], regroupV0_lo_12[2818]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo_hi_2 = {regroupV0_lo_12[2830], regroupV0_lo_12[2826]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo_6 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo_hi_2, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi_lo_2 = {regroupV0_lo_12[2838], regroupV0_lo_12[2834]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi_hi_2 = {regroupV0_lo_12[2846], regroupV0_lo_12[2842]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi_6 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi_hi_2, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_10 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi_6, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo_lo_2 = {regroupV0_lo_12[2854], regroupV0_lo_12[2850]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo_hi_2 = {regroupV0_lo_12[2862], regroupV0_lo_12[2858]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo_6 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo_hi_2, regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi_lo_2 = {regroupV0_lo_12[2870], regroupV0_lo_12[2866]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi_hi_2 = {regroupV0_lo_12[2878], regroupV0_lo_12[2874]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi_6 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi_hi_2, regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_10 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi_6, regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_lo_lo_13 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_10, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_10};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo_lo_2 = {regroupV0_lo_12[2886], regroupV0_lo_12[2882]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo_hi_2 = {regroupV0_lo_12[2894], regroupV0_lo_12[2890]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo_6 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo_hi_2, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi_lo_2 = {regroupV0_lo_12[2902], regroupV0_lo_12[2898]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi_hi_2 = {regroupV0_lo_12[2910], regroupV0_lo_12[2906]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi_6 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi_hi_2, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_10 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi_6, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo_lo_2 = {regroupV0_lo_12[2918], regroupV0_lo_12[2914]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo_hi_2 = {regroupV0_lo_12[2926], regroupV0_lo_12[2922]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo_6 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo_hi_2, regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi_lo_2 = {regroupV0_lo_12[2934], regroupV0_lo_12[2930]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi_hi_2 = {regroupV0_lo_12[2942], regroupV0_lo_12[2938]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi_6 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi_hi_2, regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_10 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi_6, regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_lo_hi_13 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_10, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_10};
  wire [31:0]        regroupV0_lo_hi_lo_hi_hi_lo_13 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_13, regroupV0_lo_hi_lo_hi_hi_lo_lo_13};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo_lo_2 = {regroupV0_lo_12[2950], regroupV0_lo_12[2946]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo_hi_2 = {regroupV0_lo_12[2958], regroupV0_lo_12[2954]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo_6 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo_hi_2, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi_lo_2 = {regroupV0_lo_12[2966], regroupV0_lo_12[2962]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi_hi_2 = {regroupV0_lo_12[2974], regroupV0_lo_12[2970]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi_6 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi_hi_2, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_10 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi_6, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo_lo_2 = {regroupV0_lo_12[2982], regroupV0_lo_12[2978]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo_hi_2 = {regroupV0_lo_12[2990], regroupV0_lo_12[2986]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo_6 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo_hi_2, regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi_lo_2 = {regroupV0_lo_12[2998], regroupV0_lo_12[2994]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi_hi_2 = {regroupV0_lo_12[3006], regroupV0_lo_12[3002]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi_6 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi_hi_2, regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_10 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi_6, regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_hi_lo_13 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_10, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_10};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo_lo_2 = {regroupV0_lo_12[3014], regroupV0_lo_12[3010]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo_hi_2 = {regroupV0_lo_12[3022], regroupV0_lo_12[3018]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo_6 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo_hi_2, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi_lo_2 = {regroupV0_lo_12[3030], regroupV0_lo_12[3026]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi_hi_2 = {regroupV0_lo_12[3038], regroupV0_lo_12[3034]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi_6 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi_hi_2, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_10 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi_6, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo_lo_2 = {regroupV0_lo_12[3046], regroupV0_lo_12[3042]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo_hi_2 = {regroupV0_lo_12[3054], regroupV0_lo_12[3050]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo_6 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo_hi_2, regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi_lo_2 = {regroupV0_lo_12[3062], regroupV0_lo_12[3058]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi_hi_2 = {regroupV0_lo_12[3070], regroupV0_lo_12[3066]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi_6 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi_hi_2, regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_10 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi_6, regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_hi_hi_13 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_10, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_10};
  wire [31:0]        regroupV0_lo_hi_lo_hi_hi_hi_13 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_13, regroupV0_lo_hi_lo_hi_hi_hi_lo_13};
  wire [63:0]        regroupV0_lo_hi_lo_hi_hi_13 = {regroupV0_lo_hi_lo_hi_hi_hi_13, regroupV0_lo_hi_lo_hi_hi_lo_13};
  wire [127:0]       regroupV0_lo_hi_lo_hi_13 = {regroupV0_lo_hi_lo_hi_hi_13, regroupV0_lo_hi_lo_hi_lo_13};
  wire [255:0]       regroupV0_lo_hi_lo_13 = {regroupV0_lo_hi_lo_hi_13, regroupV0_lo_hi_lo_lo_13};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo_lo_2 = {regroupV0_lo_12[3078], regroupV0_lo_12[3074]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo_hi_2 = {regroupV0_lo_12[3086], regroupV0_lo_12[3082]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo_6 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo_hi_2, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi_lo_2 = {regroupV0_lo_12[3094], regroupV0_lo_12[3090]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi_hi_2 = {regroupV0_lo_12[3102], regroupV0_lo_12[3098]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi_6 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi_hi_2, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_10 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi_6, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo_lo_2 = {regroupV0_lo_12[3110], regroupV0_lo_12[3106]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo_hi_2 = {regroupV0_lo_12[3118], regroupV0_lo_12[3114]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo_6 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo_hi_2, regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi_lo_2 = {regroupV0_lo_12[3126], regroupV0_lo_12[3122]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi_hi_2 = {regroupV0_lo_12[3134], regroupV0_lo_12[3130]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi_6 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi_hi_2, regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_10 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi_6, regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_lo_lo_13 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_10, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_10};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo_lo_2 = {regroupV0_lo_12[3142], regroupV0_lo_12[3138]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo_hi_2 = {regroupV0_lo_12[3150], regroupV0_lo_12[3146]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo_6 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo_hi_2, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi_lo_2 = {regroupV0_lo_12[3158], regroupV0_lo_12[3154]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi_hi_2 = {regroupV0_lo_12[3166], regroupV0_lo_12[3162]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi_6 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi_hi_2, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_10 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi_6, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo_lo_2 = {regroupV0_lo_12[3174], regroupV0_lo_12[3170]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo_hi_2 = {regroupV0_lo_12[3182], regroupV0_lo_12[3178]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo_6 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo_hi_2, regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi_lo_2 = {regroupV0_lo_12[3190], regroupV0_lo_12[3186]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi_hi_2 = {regroupV0_lo_12[3198], regroupV0_lo_12[3194]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi_6 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi_hi_2, regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_10 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi_6, regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_lo_hi_13 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_10, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_10};
  wire [31:0]        regroupV0_lo_hi_hi_lo_lo_lo_13 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_13, regroupV0_lo_hi_hi_lo_lo_lo_lo_13};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo_lo_2 = {regroupV0_lo_12[3206], regroupV0_lo_12[3202]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo_hi_2 = {regroupV0_lo_12[3214], regroupV0_lo_12[3210]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo_6 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo_hi_2, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi_lo_2 = {regroupV0_lo_12[3222], regroupV0_lo_12[3218]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi_hi_2 = {regroupV0_lo_12[3230], regroupV0_lo_12[3226]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi_6 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi_hi_2, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_10 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi_6, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo_lo_2 = {regroupV0_lo_12[3238], regroupV0_lo_12[3234]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo_hi_2 = {regroupV0_lo_12[3246], regroupV0_lo_12[3242]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo_6 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo_hi_2, regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi_lo_2 = {regroupV0_lo_12[3254], regroupV0_lo_12[3250]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi_hi_2 = {regroupV0_lo_12[3262], regroupV0_lo_12[3258]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi_6 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi_hi_2, regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_10 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi_6, regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_hi_lo_13 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_10, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_10};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo_lo_2 = {regroupV0_lo_12[3270], regroupV0_lo_12[3266]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo_hi_2 = {regroupV0_lo_12[3278], regroupV0_lo_12[3274]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo_6 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo_hi_2, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi_lo_2 = {regroupV0_lo_12[3286], regroupV0_lo_12[3282]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi_hi_2 = {regroupV0_lo_12[3294], regroupV0_lo_12[3290]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi_6 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi_hi_2, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_10 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi_6, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo_lo_2 = {regroupV0_lo_12[3302], regroupV0_lo_12[3298]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo_hi_2 = {regroupV0_lo_12[3310], regroupV0_lo_12[3306]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo_6 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo_hi_2, regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi_lo_2 = {regroupV0_lo_12[3318], regroupV0_lo_12[3314]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi_hi_2 = {regroupV0_lo_12[3326], regroupV0_lo_12[3322]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi_6 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi_hi_2, regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_10 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi_6, regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_hi_hi_13 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_10, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_10};
  wire [31:0]        regroupV0_lo_hi_hi_lo_lo_hi_13 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_13, regroupV0_lo_hi_hi_lo_lo_hi_lo_13};
  wire [63:0]        regroupV0_lo_hi_hi_lo_lo_13 = {regroupV0_lo_hi_hi_lo_lo_hi_13, regroupV0_lo_hi_hi_lo_lo_lo_13};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo_lo_2 = {regroupV0_lo_12[3334], regroupV0_lo_12[3330]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo_hi_2 = {regroupV0_lo_12[3342], regroupV0_lo_12[3338]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo_6 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo_hi_2, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi_lo_2 = {regroupV0_lo_12[3350], regroupV0_lo_12[3346]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi_hi_2 = {regroupV0_lo_12[3358], regroupV0_lo_12[3354]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi_6 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi_hi_2, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_10 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi_6, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo_lo_2 = {regroupV0_lo_12[3366], regroupV0_lo_12[3362]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo_hi_2 = {regroupV0_lo_12[3374], regroupV0_lo_12[3370]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo_6 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo_hi_2, regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi_lo_2 = {regroupV0_lo_12[3382], regroupV0_lo_12[3378]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi_hi_2 = {regroupV0_lo_12[3390], regroupV0_lo_12[3386]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi_6 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi_hi_2, regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_10 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi_6, regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_lo_lo_13 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_10, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_10};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo_lo_2 = {regroupV0_lo_12[3398], regroupV0_lo_12[3394]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo_hi_2 = {regroupV0_lo_12[3406], regroupV0_lo_12[3402]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo_6 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo_hi_2, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi_lo_2 = {regroupV0_lo_12[3414], regroupV0_lo_12[3410]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi_hi_2 = {regroupV0_lo_12[3422], regroupV0_lo_12[3418]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi_6 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi_hi_2, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_10 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi_6, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo_lo_2 = {regroupV0_lo_12[3430], regroupV0_lo_12[3426]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo_hi_2 = {regroupV0_lo_12[3438], regroupV0_lo_12[3434]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo_6 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo_hi_2, regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi_lo_2 = {regroupV0_lo_12[3446], regroupV0_lo_12[3442]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi_hi_2 = {regroupV0_lo_12[3454], regroupV0_lo_12[3450]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi_6 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi_hi_2, regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_10 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi_6, regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_lo_hi_13 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_10, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_10};
  wire [31:0]        regroupV0_lo_hi_hi_lo_hi_lo_13 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_13, regroupV0_lo_hi_hi_lo_hi_lo_lo_13};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo_lo_2 = {regroupV0_lo_12[3462], regroupV0_lo_12[3458]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo_hi_2 = {regroupV0_lo_12[3470], regroupV0_lo_12[3466]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo_6 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo_hi_2, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi_lo_2 = {regroupV0_lo_12[3478], regroupV0_lo_12[3474]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi_hi_2 = {regroupV0_lo_12[3486], regroupV0_lo_12[3482]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi_6 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi_hi_2, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_10 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi_6, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo_lo_2 = {regroupV0_lo_12[3494], regroupV0_lo_12[3490]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo_hi_2 = {regroupV0_lo_12[3502], regroupV0_lo_12[3498]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo_6 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo_hi_2, regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi_lo_2 = {regroupV0_lo_12[3510], regroupV0_lo_12[3506]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi_hi_2 = {regroupV0_lo_12[3518], regroupV0_lo_12[3514]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi_6 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi_hi_2, regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_10 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi_6, regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_hi_lo_13 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_10, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_10};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo_lo_2 = {regroupV0_lo_12[3526], regroupV0_lo_12[3522]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo_hi_2 = {regroupV0_lo_12[3534], regroupV0_lo_12[3530]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo_6 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo_hi_2, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi_lo_2 = {regroupV0_lo_12[3542], regroupV0_lo_12[3538]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi_hi_2 = {regroupV0_lo_12[3550], regroupV0_lo_12[3546]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi_6 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi_hi_2, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_10 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi_6, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo_lo_2 = {regroupV0_lo_12[3558], regroupV0_lo_12[3554]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo_hi_2 = {regroupV0_lo_12[3566], regroupV0_lo_12[3562]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo_6 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo_hi_2, regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi_lo_2 = {regroupV0_lo_12[3574], regroupV0_lo_12[3570]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi_hi_2 = {regroupV0_lo_12[3582], regroupV0_lo_12[3578]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi_6 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi_hi_2, regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_10 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi_6, regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_hi_hi_13 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_10, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_10};
  wire [31:0]        regroupV0_lo_hi_hi_lo_hi_hi_13 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_13, regroupV0_lo_hi_hi_lo_hi_hi_lo_13};
  wire [63:0]        regroupV0_lo_hi_hi_lo_hi_13 = {regroupV0_lo_hi_hi_lo_hi_hi_13, regroupV0_lo_hi_hi_lo_hi_lo_13};
  wire [127:0]       regroupV0_lo_hi_hi_lo_13 = {regroupV0_lo_hi_hi_lo_hi_13, regroupV0_lo_hi_hi_lo_lo_13};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo_lo_2 = {regroupV0_lo_12[3590], regroupV0_lo_12[3586]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo_hi_2 = {regroupV0_lo_12[3598], regroupV0_lo_12[3594]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo_6 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo_hi_2, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi_lo_2 = {regroupV0_lo_12[3606], regroupV0_lo_12[3602]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi_hi_2 = {regroupV0_lo_12[3614], regroupV0_lo_12[3610]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi_6 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi_hi_2, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_10 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi_6, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo_lo_2 = {regroupV0_lo_12[3622], regroupV0_lo_12[3618]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo_hi_2 = {regroupV0_lo_12[3630], regroupV0_lo_12[3626]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo_6 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo_hi_2, regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi_lo_2 = {regroupV0_lo_12[3638], regroupV0_lo_12[3634]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi_hi_2 = {regroupV0_lo_12[3646], regroupV0_lo_12[3642]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi_6 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi_hi_2, regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_10 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi_6, regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_lo_lo_13 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_10, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_10};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo_lo_2 = {regroupV0_lo_12[3654], regroupV0_lo_12[3650]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo_hi_2 = {regroupV0_lo_12[3662], regroupV0_lo_12[3658]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo_6 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo_hi_2, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi_lo_2 = {regroupV0_lo_12[3670], regroupV0_lo_12[3666]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi_hi_2 = {regroupV0_lo_12[3678], regroupV0_lo_12[3674]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi_6 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi_hi_2, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_10 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi_6, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo_lo_2 = {regroupV0_lo_12[3686], regroupV0_lo_12[3682]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo_hi_2 = {regroupV0_lo_12[3694], regroupV0_lo_12[3690]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo_6 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo_hi_2, regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi_lo_2 = {regroupV0_lo_12[3702], regroupV0_lo_12[3698]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi_hi_2 = {regroupV0_lo_12[3710], regroupV0_lo_12[3706]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi_6 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi_hi_2, regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_10 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi_6, regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_lo_hi_13 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_10, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_10};
  wire [31:0]        regroupV0_lo_hi_hi_hi_lo_lo_13 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_13, regroupV0_lo_hi_hi_hi_lo_lo_lo_13};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo_lo_2 = {regroupV0_lo_12[3718], regroupV0_lo_12[3714]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo_hi_2 = {regroupV0_lo_12[3726], regroupV0_lo_12[3722]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo_6 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo_hi_2, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi_lo_2 = {regroupV0_lo_12[3734], regroupV0_lo_12[3730]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi_hi_2 = {regroupV0_lo_12[3742], regroupV0_lo_12[3738]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi_6 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi_hi_2, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_10 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi_6, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo_lo_2 = {regroupV0_lo_12[3750], regroupV0_lo_12[3746]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo_hi_2 = {regroupV0_lo_12[3758], regroupV0_lo_12[3754]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo_6 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo_hi_2, regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi_lo_2 = {regroupV0_lo_12[3766], regroupV0_lo_12[3762]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi_hi_2 = {regroupV0_lo_12[3774], regroupV0_lo_12[3770]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi_6 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi_hi_2, regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_10 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi_6, regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_hi_lo_13 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_10, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_10};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo_lo_2 = {regroupV0_lo_12[3782], regroupV0_lo_12[3778]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo_hi_2 = {regroupV0_lo_12[3790], regroupV0_lo_12[3786]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo_6 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo_hi_2, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi_lo_2 = {regroupV0_lo_12[3798], regroupV0_lo_12[3794]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi_hi_2 = {regroupV0_lo_12[3806], regroupV0_lo_12[3802]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi_6 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi_hi_2, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_10 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi_6, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo_lo_2 = {regroupV0_lo_12[3814], regroupV0_lo_12[3810]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo_hi_2 = {regroupV0_lo_12[3822], regroupV0_lo_12[3818]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo_6 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo_hi_2, regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi_lo_2 = {regroupV0_lo_12[3830], regroupV0_lo_12[3826]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi_hi_2 = {regroupV0_lo_12[3838], regroupV0_lo_12[3834]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi_6 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi_hi_2, regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_10 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi_6, regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_hi_hi_13 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_10, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_10};
  wire [31:0]        regroupV0_lo_hi_hi_hi_lo_hi_13 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_13, regroupV0_lo_hi_hi_hi_lo_hi_lo_13};
  wire [63:0]        regroupV0_lo_hi_hi_hi_lo_13 = {regroupV0_lo_hi_hi_hi_lo_hi_13, regroupV0_lo_hi_hi_hi_lo_lo_13};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo_lo_2 = {regroupV0_lo_12[3846], regroupV0_lo_12[3842]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo_hi_2 = {regroupV0_lo_12[3854], regroupV0_lo_12[3850]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo_6 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo_hi_2, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi_lo_2 = {regroupV0_lo_12[3862], regroupV0_lo_12[3858]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi_hi_2 = {regroupV0_lo_12[3870], regroupV0_lo_12[3866]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi_6 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi_hi_2, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_10 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi_6, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo_lo_2 = {regroupV0_lo_12[3878], regroupV0_lo_12[3874]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo_hi_2 = {regroupV0_lo_12[3886], regroupV0_lo_12[3882]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo_6 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo_hi_2, regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi_lo_2 = {regroupV0_lo_12[3894], regroupV0_lo_12[3890]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi_hi_2 = {regroupV0_lo_12[3902], regroupV0_lo_12[3898]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi_6 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi_hi_2, regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_10 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi_6, regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_lo_lo_13 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_10, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_10};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo_lo_2 = {regroupV0_lo_12[3910], regroupV0_lo_12[3906]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo_hi_2 = {regroupV0_lo_12[3918], regroupV0_lo_12[3914]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo_6 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo_hi_2, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi_lo_2 = {regroupV0_lo_12[3926], regroupV0_lo_12[3922]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi_hi_2 = {regroupV0_lo_12[3934], regroupV0_lo_12[3930]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi_6 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi_hi_2, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_10 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi_6, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo_lo_2 = {regroupV0_lo_12[3942], regroupV0_lo_12[3938]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo_hi_2 = {regroupV0_lo_12[3950], regroupV0_lo_12[3946]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo_6 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo_hi_2, regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi_lo_2 = {regroupV0_lo_12[3958], regroupV0_lo_12[3954]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi_hi_2 = {regroupV0_lo_12[3966], regroupV0_lo_12[3962]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi_6 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi_hi_2, regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_10 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi_6, regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_lo_hi_13 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_10, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_10};
  wire [31:0]        regroupV0_lo_hi_hi_hi_hi_lo_13 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_13, regroupV0_lo_hi_hi_hi_hi_lo_lo_13};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo_lo_2 = {regroupV0_lo_12[3974], regroupV0_lo_12[3970]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo_hi_2 = {regroupV0_lo_12[3982], regroupV0_lo_12[3978]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo_6 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo_hi_2, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi_lo_2 = {regroupV0_lo_12[3990], regroupV0_lo_12[3986]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi_hi_2 = {regroupV0_lo_12[3998], regroupV0_lo_12[3994]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi_6 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi_hi_2, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_10 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi_6, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo_lo_2 = {regroupV0_lo_12[4006], regroupV0_lo_12[4002]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo_hi_2 = {regroupV0_lo_12[4014], regroupV0_lo_12[4010]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo_6 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo_hi_2, regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi_lo_2 = {regroupV0_lo_12[4022], regroupV0_lo_12[4018]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi_hi_2 = {regroupV0_lo_12[4030], regroupV0_lo_12[4026]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi_6 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi_hi_2, regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_10 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi_6, regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_hi_lo_13 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_10, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_10};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo_lo_2 = {regroupV0_lo_12[4038], regroupV0_lo_12[4034]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo_hi_2 = {regroupV0_lo_12[4046], regroupV0_lo_12[4042]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo_6 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo_hi_2, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi_lo_2 = {regroupV0_lo_12[4054], regroupV0_lo_12[4050]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi_hi_2 = {regroupV0_lo_12[4062], regroupV0_lo_12[4058]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi_6 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi_hi_2, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_10 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi_6, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo_lo_2 = {regroupV0_lo_12[4070], regroupV0_lo_12[4066]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo_hi_2 = {regroupV0_lo_12[4078], regroupV0_lo_12[4074]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo_6 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo_hi_2, regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi_lo_2 = {regroupV0_lo_12[4086], regroupV0_lo_12[4082]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi_hi_2 = {regroupV0_lo_12[4094], regroupV0_lo_12[4090]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi_6 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi_hi_2, regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_10 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi_6, regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_hi_hi_13 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_10, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_10};
  wire [31:0]        regroupV0_lo_hi_hi_hi_hi_hi_13 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_13, regroupV0_lo_hi_hi_hi_hi_hi_lo_13};
  wire [63:0]        regroupV0_lo_hi_hi_hi_hi_13 = {regroupV0_lo_hi_hi_hi_hi_hi_13, regroupV0_lo_hi_hi_hi_hi_lo_13};
  wire [127:0]       regroupV0_lo_hi_hi_hi_13 = {regroupV0_lo_hi_hi_hi_hi_13, regroupV0_lo_hi_hi_hi_lo_13};
  wire [255:0]       regroupV0_lo_hi_hi_13 = {regroupV0_lo_hi_hi_hi_13, regroupV0_lo_hi_hi_lo_13};
  wire [511:0]       regroupV0_lo_hi_13 = {regroupV0_lo_hi_hi_13, regroupV0_lo_hi_lo_13};
  wire [1023:0]      regroupV0_lo_15 = {regroupV0_lo_hi_13, regroupV0_lo_lo_13};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo_lo_2 = {regroupV0_hi_12[6], regroupV0_hi_12[2]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo_hi_2 = {regroupV0_hi_12[14], regroupV0_hi_12[10]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo_6 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi_lo_2 = {regroupV0_hi_12[22], regroupV0_hi_12[18]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi_hi_2 = {regroupV0_hi_12[30], regroupV0_hi_12[26]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi_6 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi_hi_2, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_10 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi_6, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo_lo_2 = {regroupV0_hi_12[38], regroupV0_hi_12[34]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo_hi_2 = {regroupV0_hi_12[46], regroupV0_hi_12[42]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo_6 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo_hi_2, regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi_lo_2 = {regroupV0_hi_12[54], regroupV0_hi_12[50]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi_hi_2 = {regroupV0_hi_12[62], regroupV0_hi_12[58]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi_6 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi_hi_2, regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_10 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi_6, regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_lo_lo_13 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_10, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_10};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo_lo_2 = {regroupV0_hi_12[70], regroupV0_hi_12[66]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo_hi_2 = {regroupV0_hi_12[78], regroupV0_hi_12[74]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo_6 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi_lo_2 = {regroupV0_hi_12[86], regroupV0_hi_12[82]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi_hi_2 = {regroupV0_hi_12[94], regroupV0_hi_12[90]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi_6 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi_hi_2, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_10 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi_6, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo_lo_2 = {regroupV0_hi_12[102], regroupV0_hi_12[98]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo_hi_2 = {regroupV0_hi_12[110], regroupV0_hi_12[106]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo_6 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo_hi_2, regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi_lo_2 = {regroupV0_hi_12[118], regroupV0_hi_12[114]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi_hi_2 = {regroupV0_hi_12[126], regroupV0_hi_12[122]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi_6 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi_hi_2, regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_10 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi_6, regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_lo_hi_13 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_10, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_10};
  wire [31:0]        regroupV0_hi_lo_lo_lo_lo_lo_13 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_13, regroupV0_hi_lo_lo_lo_lo_lo_lo_13};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo_lo_2 = {regroupV0_hi_12[134], regroupV0_hi_12[130]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo_hi_2 = {regroupV0_hi_12[142], regroupV0_hi_12[138]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo_6 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi_lo_2 = {regroupV0_hi_12[150], regroupV0_hi_12[146]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi_hi_2 = {regroupV0_hi_12[158], regroupV0_hi_12[154]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi_6 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi_hi_2, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_10 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi_6, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo_lo_2 = {regroupV0_hi_12[166], regroupV0_hi_12[162]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo_hi_2 = {regroupV0_hi_12[174], regroupV0_hi_12[170]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo_6 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo_hi_2, regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi_lo_2 = {regroupV0_hi_12[182], regroupV0_hi_12[178]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi_hi_2 = {regroupV0_hi_12[190], regroupV0_hi_12[186]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi_6 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi_hi_2, regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_10 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi_6, regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_hi_lo_13 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_10, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_10};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo_lo_2 = {regroupV0_hi_12[198], regroupV0_hi_12[194]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo_hi_2 = {regroupV0_hi_12[206], regroupV0_hi_12[202]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo_6 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi_lo_2 = {regroupV0_hi_12[214], regroupV0_hi_12[210]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi_hi_2 = {regroupV0_hi_12[222], regroupV0_hi_12[218]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi_6 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi_hi_2, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_10 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi_6, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo_lo_2 = {regroupV0_hi_12[230], regroupV0_hi_12[226]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo_hi_2 = {regroupV0_hi_12[238], regroupV0_hi_12[234]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo_6 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo_hi_2, regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi_lo_2 = {regroupV0_hi_12[246], regroupV0_hi_12[242]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi_hi_2 = {regroupV0_hi_12[254], regroupV0_hi_12[250]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi_6 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi_hi_2, regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_10 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi_6, regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_hi_hi_13 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_10, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_10};
  wire [31:0]        regroupV0_hi_lo_lo_lo_lo_hi_13 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_13, regroupV0_hi_lo_lo_lo_lo_hi_lo_13};
  wire [63:0]        regroupV0_hi_lo_lo_lo_lo_13 = {regroupV0_hi_lo_lo_lo_lo_hi_13, regroupV0_hi_lo_lo_lo_lo_lo_13};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo_lo_2 = {regroupV0_hi_12[262], regroupV0_hi_12[258]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo_hi_2 = {regroupV0_hi_12[270], regroupV0_hi_12[266]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo_6 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi_lo_2 = {regroupV0_hi_12[278], regroupV0_hi_12[274]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi_hi_2 = {regroupV0_hi_12[286], regroupV0_hi_12[282]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi_6 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi_hi_2, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_10 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi_6, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo_lo_2 = {regroupV0_hi_12[294], regroupV0_hi_12[290]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo_hi_2 = {regroupV0_hi_12[302], regroupV0_hi_12[298]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo_6 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo_hi_2, regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi_lo_2 = {regroupV0_hi_12[310], regroupV0_hi_12[306]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi_hi_2 = {regroupV0_hi_12[318], regroupV0_hi_12[314]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi_6 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi_hi_2, regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_10 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi_6, regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_lo_lo_13 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_10, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_10};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo_lo_2 = {regroupV0_hi_12[326], regroupV0_hi_12[322]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo_hi_2 = {regroupV0_hi_12[334], regroupV0_hi_12[330]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo_6 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi_lo_2 = {regroupV0_hi_12[342], regroupV0_hi_12[338]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi_hi_2 = {regroupV0_hi_12[350], regroupV0_hi_12[346]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi_6 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi_hi_2, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_10 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi_6, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo_lo_2 = {regroupV0_hi_12[358], regroupV0_hi_12[354]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo_hi_2 = {regroupV0_hi_12[366], regroupV0_hi_12[362]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo_6 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo_hi_2, regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi_lo_2 = {regroupV0_hi_12[374], regroupV0_hi_12[370]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi_hi_2 = {regroupV0_hi_12[382], regroupV0_hi_12[378]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi_6 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi_hi_2, regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_10 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi_6, regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_lo_hi_13 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_10, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_10};
  wire [31:0]        regroupV0_hi_lo_lo_lo_hi_lo_13 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_13, regroupV0_hi_lo_lo_lo_hi_lo_lo_13};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo_lo_2 = {regroupV0_hi_12[390], regroupV0_hi_12[386]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo_hi_2 = {regroupV0_hi_12[398], regroupV0_hi_12[394]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo_6 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi_lo_2 = {regroupV0_hi_12[406], regroupV0_hi_12[402]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi_hi_2 = {regroupV0_hi_12[414], regroupV0_hi_12[410]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi_6 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi_hi_2, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_10 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi_6, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo_lo_2 = {regroupV0_hi_12[422], regroupV0_hi_12[418]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo_hi_2 = {regroupV0_hi_12[430], regroupV0_hi_12[426]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo_6 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo_hi_2, regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi_lo_2 = {regroupV0_hi_12[438], regroupV0_hi_12[434]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi_hi_2 = {regroupV0_hi_12[446], regroupV0_hi_12[442]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi_6 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi_hi_2, regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_10 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi_6, regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_hi_lo_13 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_10, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_10};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo_lo_2 = {regroupV0_hi_12[454], regroupV0_hi_12[450]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo_hi_2 = {regroupV0_hi_12[462], regroupV0_hi_12[458]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo_6 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi_lo_2 = {regroupV0_hi_12[470], regroupV0_hi_12[466]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi_hi_2 = {regroupV0_hi_12[478], regroupV0_hi_12[474]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi_6 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi_hi_2, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_10 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi_6, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo_lo_2 = {regroupV0_hi_12[486], regroupV0_hi_12[482]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo_hi_2 = {regroupV0_hi_12[494], regroupV0_hi_12[490]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo_6 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo_hi_2, regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi_lo_2 = {regroupV0_hi_12[502], regroupV0_hi_12[498]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi_hi_2 = {regroupV0_hi_12[510], regroupV0_hi_12[506]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi_6 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi_hi_2, regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_10 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi_6, regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_hi_hi_13 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_10, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_10};
  wire [31:0]        regroupV0_hi_lo_lo_lo_hi_hi_13 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_13, regroupV0_hi_lo_lo_lo_hi_hi_lo_13};
  wire [63:0]        regroupV0_hi_lo_lo_lo_hi_13 = {regroupV0_hi_lo_lo_lo_hi_hi_13, regroupV0_hi_lo_lo_lo_hi_lo_13};
  wire [127:0]       regroupV0_hi_lo_lo_lo_13 = {regroupV0_hi_lo_lo_lo_hi_13, regroupV0_hi_lo_lo_lo_lo_13};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo_lo_2 = {regroupV0_hi_12[518], regroupV0_hi_12[514]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo_hi_2 = {regroupV0_hi_12[526], regroupV0_hi_12[522]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo_6 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo_hi_2, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi_lo_2 = {regroupV0_hi_12[534], regroupV0_hi_12[530]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi_hi_2 = {regroupV0_hi_12[542], regroupV0_hi_12[538]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi_6 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi_hi_2, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_10 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi_6, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo_lo_2 = {regroupV0_hi_12[550], regroupV0_hi_12[546]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo_hi_2 = {regroupV0_hi_12[558], regroupV0_hi_12[554]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo_6 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo_hi_2, regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi_lo_2 = {regroupV0_hi_12[566], regroupV0_hi_12[562]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi_hi_2 = {regroupV0_hi_12[574], regroupV0_hi_12[570]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi_6 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi_hi_2, regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_10 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi_6, regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_lo_lo_13 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_10, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_10};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo_lo_2 = {regroupV0_hi_12[582], regroupV0_hi_12[578]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo_hi_2 = {regroupV0_hi_12[590], regroupV0_hi_12[586]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo_6 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo_hi_2, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi_lo_2 = {regroupV0_hi_12[598], regroupV0_hi_12[594]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi_hi_2 = {regroupV0_hi_12[606], regroupV0_hi_12[602]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi_6 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi_hi_2, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_10 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi_6, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo_lo_2 = {regroupV0_hi_12[614], regroupV0_hi_12[610]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo_hi_2 = {regroupV0_hi_12[622], regroupV0_hi_12[618]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo_6 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo_hi_2, regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi_lo_2 = {regroupV0_hi_12[630], regroupV0_hi_12[626]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi_hi_2 = {regroupV0_hi_12[638], regroupV0_hi_12[634]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi_6 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi_hi_2, regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_10 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi_6, regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_lo_hi_13 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_10, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_10};
  wire [31:0]        regroupV0_hi_lo_lo_hi_lo_lo_13 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_13, regroupV0_hi_lo_lo_hi_lo_lo_lo_13};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo_lo_2 = {regroupV0_hi_12[646], regroupV0_hi_12[642]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo_hi_2 = {regroupV0_hi_12[654], regroupV0_hi_12[650]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo_6 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo_hi_2, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi_lo_2 = {regroupV0_hi_12[662], regroupV0_hi_12[658]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi_hi_2 = {regroupV0_hi_12[670], regroupV0_hi_12[666]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi_6 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi_hi_2, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_10 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi_6, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo_lo_2 = {regroupV0_hi_12[678], regroupV0_hi_12[674]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo_hi_2 = {regroupV0_hi_12[686], regroupV0_hi_12[682]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo_6 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo_hi_2, regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi_lo_2 = {regroupV0_hi_12[694], regroupV0_hi_12[690]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi_hi_2 = {regroupV0_hi_12[702], regroupV0_hi_12[698]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi_6 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi_hi_2, regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_10 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi_6, regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_hi_lo_13 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_10, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_10};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo_lo_2 = {regroupV0_hi_12[710], regroupV0_hi_12[706]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo_hi_2 = {regroupV0_hi_12[718], regroupV0_hi_12[714]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo_6 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo_hi_2, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi_lo_2 = {regroupV0_hi_12[726], regroupV0_hi_12[722]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi_hi_2 = {regroupV0_hi_12[734], regroupV0_hi_12[730]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi_6 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi_hi_2, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_10 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi_6, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo_lo_2 = {regroupV0_hi_12[742], regroupV0_hi_12[738]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo_hi_2 = {regroupV0_hi_12[750], regroupV0_hi_12[746]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo_6 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo_hi_2, regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi_lo_2 = {regroupV0_hi_12[758], regroupV0_hi_12[754]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi_hi_2 = {regroupV0_hi_12[766], regroupV0_hi_12[762]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi_6 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi_hi_2, regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_10 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi_6, regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_hi_hi_13 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_10, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_10};
  wire [31:0]        regroupV0_hi_lo_lo_hi_lo_hi_13 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_13, regroupV0_hi_lo_lo_hi_lo_hi_lo_13};
  wire [63:0]        regroupV0_hi_lo_lo_hi_lo_13 = {regroupV0_hi_lo_lo_hi_lo_hi_13, regroupV0_hi_lo_lo_hi_lo_lo_13};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo_lo_2 = {regroupV0_hi_12[774], regroupV0_hi_12[770]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo_hi_2 = {regroupV0_hi_12[782], regroupV0_hi_12[778]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo_6 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo_hi_2, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi_lo_2 = {regroupV0_hi_12[790], regroupV0_hi_12[786]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi_hi_2 = {regroupV0_hi_12[798], regroupV0_hi_12[794]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi_6 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi_hi_2, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_10 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi_6, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo_lo_2 = {regroupV0_hi_12[806], regroupV0_hi_12[802]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo_hi_2 = {regroupV0_hi_12[814], regroupV0_hi_12[810]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo_6 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo_hi_2, regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi_lo_2 = {regroupV0_hi_12[822], regroupV0_hi_12[818]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi_hi_2 = {regroupV0_hi_12[830], regroupV0_hi_12[826]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi_6 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi_hi_2, regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_10 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi_6, regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_lo_lo_13 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_10, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_10};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo_lo_2 = {regroupV0_hi_12[838], regroupV0_hi_12[834]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo_hi_2 = {regroupV0_hi_12[846], regroupV0_hi_12[842]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo_6 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo_hi_2, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi_lo_2 = {regroupV0_hi_12[854], regroupV0_hi_12[850]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi_hi_2 = {regroupV0_hi_12[862], regroupV0_hi_12[858]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi_6 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi_hi_2, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_10 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi_6, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo_lo_2 = {regroupV0_hi_12[870], regroupV0_hi_12[866]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo_hi_2 = {regroupV0_hi_12[878], regroupV0_hi_12[874]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo_6 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo_hi_2, regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi_lo_2 = {regroupV0_hi_12[886], regroupV0_hi_12[882]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi_hi_2 = {regroupV0_hi_12[894], regroupV0_hi_12[890]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi_6 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi_hi_2, regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_10 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi_6, regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_lo_hi_13 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_10, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_10};
  wire [31:0]        regroupV0_hi_lo_lo_hi_hi_lo_13 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_13, regroupV0_hi_lo_lo_hi_hi_lo_lo_13};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo_lo_2 = {regroupV0_hi_12[902], regroupV0_hi_12[898]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo_hi_2 = {regroupV0_hi_12[910], regroupV0_hi_12[906]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo_6 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo_hi_2, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi_lo_2 = {regroupV0_hi_12[918], regroupV0_hi_12[914]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi_hi_2 = {regroupV0_hi_12[926], regroupV0_hi_12[922]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi_6 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi_hi_2, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_10 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi_6, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo_lo_2 = {regroupV0_hi_12[934], regroupV0_hi_12[930]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo_hi_2 = {regroupV0_hi_12[942], regroupV0_hi_12[938]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo_6 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo_hi_2, regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi_lo_2 = {regroupV0_hi_12[950], regroupV0_hi_12[946]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi_hi_2 = {regroupV0_hi_12[958], regroupV0_hi_12[954]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi_6 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi_hi_2, regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_10 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi_6, regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_hi_lo_13 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_10, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_10};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo_lo_2 = {regroupV0_hi_12[966], regroupV0_hi_12[962]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo_hi_2 = {regroupV0_hi_12[974], regroupV0_hi_12[970]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo_6 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo_hi_2, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi_lo_2 = {regroupV0_hi_12[982], regroupV0_hi_12[978]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi_hi_2 = {regroupV0_hi_12[990], regroupV0_hi_12[986]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi_6 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi_hi_2, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_10 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi_6, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo_lo_2 = {regroupV0_hi_12[998], regroupV0_hi_12[994]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo_hi_2 = {regroupV0_hi_12[1006], regroupV0_hi_12[1002]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo_6 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo_hi_2, regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi_lo_2 = {regroupV0_hi_12[1014], regroupV0_hi_12[1010]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi_hi_2 = {regroupV0_hi_12[1022], regroupV0_hi_12[1018]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi_6 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi_hi_2, regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_10 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi_6, regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_hi_hi_13 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_10, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_10};
  wire [31:0]        regroupV0_hi_lo_lo_hi_hi_hi_13 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_13, regroupV0_hi_lo_lo_hi_hi_hi_lo_13};
  wire [63:0]        regroupV0_hi_lo_lo_hi_hi_13 = {regroupV0_hi_lo_lo_hi_hi_hi_13, regroupV0_hi_lo_lo_hi_hi_lo_13};
  wire [127:0]       regroupV0_hi_lo_lo_hi_13 = {regroupV0_hi_lo_lo_hi_hi_13, regroupV0_hi_lo_lo_hi_lo_13};
  wire [255:0]       regroupV0_hi_lo_lo_13 = {regroupV0_hi_lo_lo_hi_13, regroupV0_hi_lo_lo_lo_13};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo_lo_2 = {regroupV0_hi_12[1030], regroupV0_hi_12[1026]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo_hi_2 = {regroupV0_hi_12[1038], regroupV0_hi_12[1034]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo_6 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo_hi_2, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi_lo_2 = {regroupV0_hi_12[1046], regroupV0_hi_12[1042]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi_hi_2 = {regroupV0_hi_12[1054], regroupV0_hi_12[1050]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi_6 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi_hi_2, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_10 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi_6, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo_lo_2 = {regroupV0_hi_12[1062], regroupV0_hi_12[1058]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo_hi_2 = {regroupV0_hi_12[1070], regroupV0_hi_12[1066]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo_6 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo_hi_2, regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi_lo_2 = {regroupV0_hi_12[1078], regroupV0_hi_12[1074]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi_hi_2 = {regroupV0_hi_12[1086], regroupV0_hi_12[1082]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi_6 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi_hi_2, regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_10 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi_6, regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_lo_lo_13 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_10, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_10};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo_lo_2 = {regroupV0_hi_12[1094], regroupV0_hi_12[1090]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo_hi_2 = {regroupV0_hi_12[1102], regroupV0_hi_12[1098]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo_6 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo_hi_2, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi_lo_2 = {regroupV0_hi_12[1110], regroupV0_hi_12[1106]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi_hi_2 = {regroupV0_hi_12[1118], regroupV0_hi_12[1114]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi_6 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi_hi_2, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_10 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi_6, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo_lo_2 = {regroupV0_hi_12[1126], regroupV0_hi_12[1122]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo_hi_2 = {regroupV0_hi_12[1134], regroupV0_hi_12[1130]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo_6 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo_hi_2, regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi_lo_2 = {regroupV0_hi_12[1142], regroupV0_hi_12[1138]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi_hi_2 = {regroupV0_hi_12[1150], regroupV0_hi_12[1146]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi_6 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi_hi_2, regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_10 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi_6, regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_lo_hi_13 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_10, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_10};
  wire [31:0]        regroupV0_hi_lo_hi_lo_lo_lo_13 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_13, regroupV0_hi_lo_hi_lo_lo_lo_lo_13};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo_lo_2 = {regroupV0_hi_12[1158], regroupV0_hi_12[1154]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo_hi_2 = {regroupV0_hi_12[1166], regroupV0_hi_12[1162]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo_6 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo_hi_2, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi_lo_2 = {regroupV0_hi_12[1174], regroupV0_hi_12[1170]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi_hi_2 = {regroupV0_hi_12[1182], regroupV0_hi_12[1178]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi_6 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi_hi_2, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_10 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi_6, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo_lo_2 = {regroupV0_hi_12[1190], regroupV0_hi_12[1186]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo_hi_2 = {regroupV0_hi_12[1198], regroupV0_hi_12[1194]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo_6 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo_hi_2, regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi_lo_2 = {regroupV0_hi_12[1206], regroupV0_hi_12[1202]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi_hi_2 = {regroupV0_hi_12[1214], regroupV0_hi_12[1210]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi_6 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi_hi_2, regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_10 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi_6, regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_hi_lo_13 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_10, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_10};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo_lo_2 = {regroupV0_hi_12[1222], regroupV0_hi_12[1218]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo_hi_2 = {regroupV0_hi_12[1230], regroupV0_hi_12[1226]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo_6 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo_hi_2, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi_lo_2 = {regroupV0_hi_12[1238], regroupV0_hi_12[1234]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi_hi_2 = {regroupV0_hi_12[1246], regroupV0_hi_12[1242]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi_6 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi_hi_2, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_10 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi_6, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo_lo_2 = {regroupV0_hi_12[1254], regroupV0_hi_12[1250]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo_hi_2 = {regroupV0_hi_12[1262], regroupV0_hi_12[1258]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo_6 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo_hi_2, regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi_lo_2 = {regroupV0_hi_12[1270], regroupV0_hi_12[1266]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi_hi_2 = {regroupV0_hi_12[1278], regroupV0_hi_12[1274]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi_6 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi_hi_2, regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_10 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi_6, regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_hi_hi_13 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_10, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_10};
  wire [31:0]        regroupV0_hi_lo_hi_lo_lo_hi_13 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_13, regroupV0_hi_lo_hi_lo_lo_hi_lo_13};
  wire [63:0]        regroupV0_hi_lo_hi_lo_lo_13 = {regroupV0_hi_lo_hi_lo_lo_hi_13, regroupV0_hi_lo_hi_lo_lo_lo_13};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo_lo_2 = {regroupV0_hi_12[1286], regroupV0_hi_12[1282]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo_hi_2 = {regroupV0_hi_12[1294], regroupV0_hi_12[1290]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo_6 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo_hi_2, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi_lo_2 = {regroupV0_hi_12[1302], regroupV0_hi_12[1298]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi_hi_2 = {regroupV0_hi_12[1310], regroupV0_hi_12[1306]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi_6 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi_hi_2, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_10 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi_6, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo_lo_2 = {regroupV0_hi_12[1318], regroupV0_hi_12[1314]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo_hi_2 = {regroupV0_hi_12[1326], regroupV0_hi_12[1322]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo_6 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo_hi_2, regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi_lo_2 = {regroupV0_hi_12[1334], regroupV0_hi_12[1330]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi_hi_2 = {regroupV0_hi_12[1342], regroupV0_hi_12[1338]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi_6 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi_hi_2, regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_10 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi_6, regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_lo_lo_13 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_10, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_10};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo_lo_2 = {regroupV0_hi_12[1350], regroupV0_hi_12[1346]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo_hi_2 = {regroupV0_hi_12[1358], regroupV0_hi_12[1354]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo_6 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo_hi_2, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi_lo_2 = {regroupV0_hi_12[1366], regroupV0_hi_12[1362]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi_hi_2 = {regroupV0_hi_12[1374], regroupV0_hi_12[1370]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi_6 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi_hi_2, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_10 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi_6, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo_lo_2 = {regroupV0_hi_12[1382], regroupV0_hi_12[1378]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo_hi_2 = {regroupV0_hi_12[1390], regroupV0_hi_12[1386]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo_6 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo_hi_2, regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi_lo_2 = {regroupV0_hi_12[1398], regroupV0_hi_12[1394]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi_hi_2 = {regroupV0_hi_12[1406], regroupV0_hi_12[1402]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi_6 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi_hi_2, regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_10 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi_6, regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_lo_hi_13 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_10, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_10};
  wire [31:0]        regroupV0_hi_lo_hi_lo_hi_lo_13 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_13, regroupV0_hi_lo_hi_lo_hi_lo_lo_13};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo_lo_2 = {regroupV0_hi_12[1414], regroupV0_hi_12[1410]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo_hi_2 = {regroupV0_hi_12[1422], regroupV0_hi_12[1418]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo_6 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo_hi_2, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi_lo_2 = {regroupV0_hi_12[1430], regroupV0_hi_12[1426]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi_hi_2 = {regroupV0_hi_12[1438], regroupV0_hi_12[1434]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi_6 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi_hi_2, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_10 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi_6, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo_lo_2 = {regroupV0_hi_12[1446], regroupV0_hi_12[1442]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo_hi_2 = {regroupV0_hi_12[1454], regroupV0_hi_12[1450]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo_6 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo_hi_2, regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi_lo_2 = {regroupV0_hi_12[1462], regroupV0_hi_12[1458]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi_hi_2 = {regroupV0_hi_12[1470], regroupV0_hi_12[1466]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi_6 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi_hi_2, regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_10 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi_6, regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_hi_lo_13 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_10, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_10};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo_lo_2 = {regroupV0_hi_12[1478], regroupV0_hi_12[1474]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo_hi_2 = {regroupV0_hi_12[1486], regroupV0_hi_12[1482]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo_6 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo_hi_2, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi_lo_2 = {regroupV0_hi_12[1494], regroupV0_hi_12[1490]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi_hi_2 = {regroupV0_hi_12[1502], regroupV0_hi_12[1498]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi_6 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi_hi_2, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_10 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi_6, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo_lo_2 = {regroupV0_hi_12[1510], regroupV0_hi_12[1506]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo_hi_2 = {regroupV0_hi_12[1518], regroupV0_hi_12[1514]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo_6 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo_hi_2, regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi_lo_2 = {regroupV0_hi_12[1526], regroupV0_hi_12[1522]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi_hi_2 = {regroupV0_hi_12[1534], regroupV0_hi_12[1530]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi_6 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi_hi_2, regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_10 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi_6, regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_hi_hi_13 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_10, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_10};
  wire [31:0]        regroupV0_hi_lo_hi_lo_hi_hi_13 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_13, regroupV0_hi_lo_hi_lo_hi_hi_lo_13};
  wire [63:0]        regroupV0_hi_lo_hi_lo_hi_13 = {regroupV0_hi_lo_hi_lo_hi_hi_13, regroupV0_hi_lo_hi_lo_hi_lo_13};
  wire [127:0]       regroupV0_hi_lo_hi_lo_13 = {regroupV0_hi_lo_hi_lo_hi_13, regroupV0_hi_lo_hi_lo_lo_13};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo_lo_2 = {regroupV0_hi_12[1542], regroupV0_hi_12[1538]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo_hi_2 = {regroupV0_hi_12[1550], regroupV0_hi_12[1546]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo_6 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo_hi_2, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi_lo_2 = {regroupV0_hi_12[1558], regroupV0_hi_12[1554]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi_hi_2 = {regroupV0_hi_12[1566], regroupV0_hi_12[1562]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi_6 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi_hi_2, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_10 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi_6, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo_lo_2 = {regroupV0_hi_12[1574], regroupV0_hi_12[1570]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo_hi_2 = {regroupV0_hi_12[1582], regroupV0_hi_12[1578]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo_6 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo_hi_2, regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi_lo_2 = {regroupV0_hi_12[1590], regroupV0_hi_12[1586]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi_hi_2 = {regroupV0_hi_12[1598], regroupV0_hi_12[1594]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi_6 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi_hi_2, regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_10 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi_6, regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_lo_lo_13 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_10, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_10};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo_lo_2 = {regroupV0_hi_12[1606], regroupV0_hi_12[1602]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo_hi_2 = {regroupV0_hi_12[1614], regroupV0_hi_12[1610]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo_6 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo_hi_2, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi_lo_2 = {regroupV0_hi_12[1622], regroupV0_hi_12[1618]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi_hi_2 = {regroupV0_hi_12[1630], regroupV0_hi_12[1626]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi_6 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi_hi_2, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_10 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi_6, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo_lo_2 = {regroupV0_hi_12[1638], regroupV0_hi_12[1634]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo_hi_2 = {regroupV0_hi_12[1646], regroupV0_hi_12[1642]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo_6 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo_hi_2, regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi_lo_2 = {regroupV0_hi_12[1654], regroupV0_hi_12[1650]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi_hi_2 = {regroupV0_hi_12[1662], regroupV0_hi_12[1658]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi_6 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi_hi_2, regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_10 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi_6, regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_lo_hi_13 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_10, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_10};
  wire [31:0]        regroupV0_hi_lo_hi_hi_lo_lo_13 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_13, regroupV0_hi_lo_hi_hi_lo_lo_lo_13};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo_lo_2 = {regroupV0_hi_12[1670], regroupV0_hi_12[1666]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo_hi_2 = {regroupV0_hi_12[1678], regroupV0_hi_12[1674]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo_6 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo_hi_2, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi_lo_2 = {regroupV0_hi_12[1686], regroupV0_hi_12[1682]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi_hi_2 = {regroupV0_hi_12[1694], regroupV0_hi_12[1690]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi_6 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi_hi_2, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_10 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi_6, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo_lo_2 = {regroupV0_hi_12[1702], regroupV0_hi_12[1698]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo_hi_2 = {regroupV0_hi_12[1710], regroupV0_hi_12[1706]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo_6 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo_hi_2, regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi_lo_2 = {regroupV0_hi_12[1718], regroupV0_hi_12[1714]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi_hi_2 = {regroupV0_hi_12[1726], regroupV0_hi_12[1722]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi_6 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi_hi_2, regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_10 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi_6, regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_hi_lo_13 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_10, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_10};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo_lo_2 = {regroupV0_hi_12[1734], regroupV0_hi_12[1730]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo_hi_2 = {regroupV0_hi_12[1742], regroupV0_hi_12[1738]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo_6 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo_hi_2, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi_lo_2 = {regroupV0_hi_12[1750], regroupV0_hi_12[1746]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi_hi_2 = {regroupV0_hi_12[1758], regroupV0_hi_12[1754]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi_6 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi_hi_2, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_10 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi_6, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo_lo_2 = {regroupV0_hi_12[1766], regroupV0_hi_12[1762]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo_hi_2 = {regroupV0_hi_12[1774], regroupV0_hi_12[1770]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo_6 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo_hi_2, regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi_lo_2 = {regroupV0_hi_12[1782], regroupV0_hi_12[1778]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi_hi_2 = {regroupV0_hi_12[1790], regroupV0_hi_12[1786]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi_6 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi_hi_2, regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_10 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi_6, regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_hi_hi_13 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_10, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_10};
  wire [31:0]        regroupV0_hi_lo_hi_hi_lo_hi_13 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_13, regroupV0_hi_lo_hi_hi_lo_hi_lo_13};
  wire [63:0]        regroupV0_hi_lo_hi_hi_lo_13 = {regroupV0_hi_lo_hi_hi_lo_hi_13, regroupV0_hi_lo_hi_hi_lo_lo_13};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo_lo_2 = {regroupV0_hi_12[1798], regroupV0_hi_12[1794]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo_hi_2 = {regroupV0_hi_12[1806], regroupV0_hi_12[1802]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo_6 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo_hi_2, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi_lo_2 = {regroupV0_hi_12[1814], regroupV0_hi_12[1810]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi_hi_2 = {regroupV0_hi_12[1822], regroupV0_hi_12[1818]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi_6 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi_hi_2, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_10 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi_6, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo_lo_2 = {regroupV0_hi_12[1830], regroupV0_hi_12[1826]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo_hi_2 = {regroupV0_hi_12[1838], regroupV0_hi_12[1834]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo_6 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo_hi_2, regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi_lo_2 = {regroupV0_hi_12[1846], regroupV0_hi_12[1842]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi_hi_2 = {regroupV0_hi_12[1854], regroupV0_hi_12[1850]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi_6 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi_hi_2, regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_10 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi_6, regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_lo_lo_13 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_10, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_10};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo_lo_2 = {regroupV0_hi_12[1862], regroupV0_hi_12[1858]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo_hi_2 = {regroupV0_hi_12[1870], regroupV0_hi_12[1866]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo_6 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo_hi_2, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi_lo_2 = {regroupV0_hi_12[1878], regroupV0_hi_12[1874]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi_hi_2 = {regroupV0_hi_12[1886], regroupV0_hi_12[1882]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi_6 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi_hi_2, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_10 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi_6, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo_lo_2 = {regroupV0_hi_12[1894], regroupV0_hi_12[1890]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo_hi_2 = {regroupV0_hi_12[1902], regroupV0_hi_12[1898]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo_6 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo_hi_2, regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi_lo_2 = {regroupV0_hi_12[1910], regroupV0_hi_12[1906]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi_hi_2 = {regroupV0_hi_12[1918], regroupV0_hi_12[1914]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi_6 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi_hi_2, regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_10 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi_6, regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_lo_hi_13 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_10, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_10};
  wire [31:0]        regroupV0_hi_lo_hi_hi_hi_lo_13 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_13, regroupV0_hi_lo_hi_hi_hi_lo_lo_13};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo_lo_2 = {regroupV0_hi_12[1926], regroupV0_hi_12[1922]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo_hi_2 = {regroupV0_hi_12[1934], regroupV0_hi_12[1930]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo_6 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo_hi_2, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi_lo_2 = {regroupV0_hi_12[1942], regroupV0_hi_12[1938]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi_hi_2 = {regroupV0_hi_12[1950], regroupV0_hi_12[1946]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi_6 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi_hi_2, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_10 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi_6, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo_lo_2 = {regroupV0_hi_12[1958], regroupV0_hi_12[1954]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo_hi_2 = {regroupV0_hi_12[1966], regroupV0_hi_12[1962]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo_6 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo_hi_2, regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi_lo_2 = {regroupV0_hi_12[1974], regroupV0_hi_12[1970]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi_hi_2 = {regroupV0_hi_12[1982], regroupV0_hi_12[1978]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi_6 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi_hi_2, regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_10 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi_6, regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_hi_lo_13 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_10, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_10};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo_lo_2 = {regroupV0_hi_12[1990], regroupV0_hi_12[1986]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo_hi_2 = {regroupV0_hi_12[1998], regroupV0_hi_12[1994]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo_6 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo_hi_2, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi_lo_2 = {regroupV0_hi_12[2006], regroupV0_hi_12[2002]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi_hi_2 = {regroupV0_hi_12[2014], regroupV0_hi_12[2010]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi_6 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi_hi_2, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_10 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi_6, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo_lo_2 = {regroupV0_hi_12[2022], regroupV0_hi_12[2018]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo_hi_2 = {regroupV0_hi_12[2030], regroupV0_hi_12[2026]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo_6 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo_hi_2, regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi_lo_2 = {regroupV0_hi_12[2038], regroupV0_hi_12[2034]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi_hi_2 = {regroupV0_hi_12[2046], regroupV0_hi_12[2042]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi_6 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi_hi_2, regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_10 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi_6, regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_hi_hi_13 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_10, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_10};
  wire [31:0]        regroupV0_hi_lo_hi_hi_hi_hi_13 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_13, regroupV0_hi_lo_hi_hi_hi_hi_lo_13};
  wire [63:0]        regroupV0_hi_lo_hi_hi_hi_13 = {regroupV0_hi_lo_hi_hi_hi_hi_13, regroupV0_hi_lo_hi_hi_hi_lo_13};
  wire [127:0]       regroupV0_hi_lo_hi_hi_13 = {regroupV0_hi_lo_hi_hi_hi_13, regroupV0_hi_lo_hi_hi_lo_13};
  wire [255:0]       regroupV0_hi_lo_hi_13 = {regroupV0_hi_lo_hi_hi_13, regroupV0_hi_lo_hi_lo_13};
  wire [511:0]       regroupV0_hi_lo_13 = {regroupV0_hi_lo_hi_13, regroupV0_hi_lo_lo_13};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo_lo_2 = {regroupV0_hi_12[2054], regroupV0_hi_12[2050]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo_hi_2 = {regroupV0_hi_12[2062], regroupV0_hi_12[2058]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo_6 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo_hi_2, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi_lo_2 = {regroupV0_hi_12[2070], regroupV0_hi_12[2066]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi_hi_2 = {regroupV0_hi_12[2078], regroupV0_hi_12[2074]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi_6 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi_hi_2, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_10 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi_6, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo_lo_2 = {regroupV0_hi_12[2086], regroupV0_hi_12[2082]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo_hi_2 = {regroupV0_hi_12[2094], regroupV0_hi_12[2090]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo_6 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo_hi_2, regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi_lo_2 = {regroupV0_hi_12[2102], regroupV0_hi_12[2098]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi_hi_2 = {regroupV0_hi_12[2110], regroupV0_hi_12[2106]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi_6 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi_hi_2, regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_10 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi_6, regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_lo_lo_13 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_10, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_10};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo_lo_2 = {regroupV0_hi_12[2118], regroupV0_hi_12[2114]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo_hi_2 = {regroupV0_hi_12[2126], regroupV0_hi_12[2122]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo_6 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo_hi_2, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi_lo_2 = {regroupV0_hi_12[2134], regroupV0_hi_12[2130]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi_hi_2 = {regroupV0_hi_12[2142], regroupV0_hi_12[2138]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi_6 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi_hi_2, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_10 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi_6, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo_lo_2 = {regroupV0_hi_12[2150], regroupV0_hi_12[2146]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo_hi_2 = {regroupV0_hi_12[2158], regroupV0_hi_12[2154]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo_6 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo_hi_2, regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi_lo_2 = {regroupV0_hi_12[2166], regroupV0_hi_12[2162]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi_hi_2 = {regroupV0_hi_12[2174], regroupV0_hi_12[2170]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi_6 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi_hi_2, regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_10 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi_6, regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_lo_hi_13 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_10, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_10};
  wire [31:0]        regroupV0_hi_hi_lo_lo_lo_lo_13 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_13, regroupV0_hi_hi_lo_lo_lo_lo_lo_13};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo_lo_2 = {regroupV0_hi_12[2182], regroupV0_hi_12[2178]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo_hi_2 = {regroupV0_hi_12[2190], regroupV0_hi_12[2186]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo_6 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo_hi_2, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi_lo_2 = {regroupV0_hi_12[2198], regroupV0_hi_12[2194]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi_hi_2 = {regroupV0_hi_12[2206], regroupV0_hi_12[2202]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi_6 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi_hi_2, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_10 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi_6, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo_lo_2 = {regroupV0_hi_12[2214], regroupV0_hi_12[2210]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo_hi_2 = {regroupV0_hi_12[2222], regroupV0_hi_12[2218]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo_6 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo_hi_2, regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi_lo_2 = {regroupV0_hi_12[2230], regroupV0_hi_12[2226]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi_hi_2 = {regroupV0_hi_12[2238], regroupV0_hi_12[2234]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi_6 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi_hi_2, regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_10 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi_6, regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_hi_lo_13 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_10, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_10};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo_lo_2 = {regroupV0_hi_12[2246], regroupV0_hi_12[2242]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo_hi_2 = {regroupV0_hi_12[2254], regroupV0_hi_12[2250]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo_6 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo_hi_2, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi_lo_2 = {regroupV0_hi_12[2262], regroupV0_hi_12[2258]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi_hi_2 = {regroupV0_hi_12[2270], regroupV0_hi_12[2266]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi_6 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi_hi_2, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_10 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi_6, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo_lo_2 = {regroupV0_hi_12[2278], regroupV0_hi_12[2274]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo_hi_2 = {regroupV0_hi_12[2286], regroupV0_hi_12[2282]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo_6 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo_hi_2, regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi_lo_2 = {regroupV0_hi_12[2294], regroupV0_hi_12[2290]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi_hi_2 = {regroupV0_hi_12[2302], regroupV0_hi_12[2298]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi_6 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi_hi_2, regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_10 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi_6, regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_hi_hi_13 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_10, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_10};
  wire [31:0]        regroupV0_hi_hi_lo_lo_lo_hi_13 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_13, regroupV0_hi_hi_lo_lo_lo_hi_lo_13};
  wire [63:0]        regroupV0_hi_hi_lo_lo_lo_13 = {regroupV0_hi_hi_lo_lo_lo_hi_13, regroupV0_hi_hi_lo_lo_lo_lo_13};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo_lo_2 = {regroupV0_hi_12[2310], regroupV0_hi_12[2306]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo_hi_2 = {regroupV0_hi_12[2318], regroupV0_hi_12[2314]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo_6 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo_hi_2, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi_lo_2 = {regroupV0_hi_12[2326], regroupV0_hi_12[2322]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi_hi_2 = {regroupV0_hi_12[2334], regroupV0_hi_12[2330]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi_6 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi_hi_2, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_10 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi_6, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo_lo_2 = {regroupV0_hi_12[2342], regroupV0_hi_12[2338]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo_hi_2 = {regroupV0_hi_12[2350], regroupV0_hi_12[2346]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo_6 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo_hi_2, regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi_lo_2 = {regroupV0_hi_12[2358], regroupV0_hi_12[2354]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi_hi_2 = {regroupV0_hi_12[2366], regroupV0_hi_12[2362]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi_6 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi_hi_2, regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_10 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi_6, regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_lo_lo_13 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_10, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_10};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo_lo_2 = {regroupV0_hi_12[2374], regroupV0_hi_12[2370]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo_hi_2 = {regroupV0_hi_12[2382], regroupV0_hi_12[2378]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo_6 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo_hi_2, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi_lo_2 = {regroupV0_hi_12[2390], regroupV0_hi_12[2386]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi_hi_2 = {regroupV0_hi_12[2398], regroupV0_hi_12[2394]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi_6 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi_hi_2, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_10 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi_6, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo_lo_2 = {regroupV0_hi_12[2406], regroupV0_hi_12[2402]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo_hi_2 = {regroupV0_hi_12[2414], regroupV0_hi_12[2410]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo_6 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo_hi_2, regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi_lo_2 = {regroupV0_hi_12[2422], regroupV0_hi_12[2418]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi_hi_2 = {regroupV0_hi_12[2430], regroupV0_hi_12[2426]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi_6 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi_hi_2, regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_10 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi_6, regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_lo_hi_13 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_10, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_10};
  wire [31:0]        regroupV0_hi_hi_lo_lo_hi_lo_13 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_13, regroupV0_hi_hi_lo_lo_hi_lo_lo_13};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo_lo_2 = {regroupV0_hi_12[2438], regroupV0_hi_12[2434]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo_hi_2 = {regroupV0_hi_12[2446], regroupV0_hi_12[2442]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo_6 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo_hi_2, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi_lo_2 = {regroupV0_hi_12[2454], regroupV0_hi_12[2450]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi_hi_2 = {regroupV0_hi_12[2462], regroupV0_hi_12[2458]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi_6 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi_hi_2, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_10 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi_6, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo_lo_2 = {regroupV0_hi_12[2470], regroupV0_hi_12[2466]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo_hi_2 = {regroupV0_hi_12[2478], regroupV0_hi_12[2474]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo_6 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo_hi_2, regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi_lo_2 = {regroupV0_hi_12[2486], regroupV0_hi_12[2482]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi_hi_2 = {regroupV0_hi_12[2494], regroupV0_hi_12[2490]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi_6 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi_hi_2, regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_10 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi_6, regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_hi_lo_13 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_10, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_10};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo_lo_2 = {regroupV0_hi_12[2502], regroupV0_hi_12[2498]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo_hi_2 = {regroupV0_hi_12[2510], regroupV0_hi_12[2506]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo_6 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo_hi_2, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi_lo_2 = {regroupV0_hi_12[2518], regroupV0_hi_12[2514]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi_hi_2 = {regroupV0_hi_12[2526], regroupV0_hi_12[2522]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi_6 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi_hi_2, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_10 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi_6, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo_lo_2 = {regroupV0_hi_12[2534], regroupV0_hi_12[2530]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo_hi_2 = {regroupV0_hi_12[2542], regroupV0_hi_12[2538]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo_6 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo_hi_2, regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi_lo_2 = {regroupV0_hi_12[2550], regroupV0_hi_12[2546]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi_hi_2 = {regroupV0_hi_12[2558], regroupV0_hi_12[2554]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi_6 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi_hi_2, regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_10 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi_6, regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_hi_hi_13 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_10, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_10};
  wire [31:0]        regroupV0_hi_hi_lo_lo_hi_hi_13 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_13, regroupV0_hi_hi_lo_lo_hi_hi_lo_13};
  wire [63:0]        regroupV0_hi_hi_lo_lo_hi_13 = {regroupV0_hi_hi_lo_lo_hi_hi_13, regroupV0_hi_hi_lo_lo_hi_lo_13};
  wire [127:0]       regroupV0_hi_hi_lo_lo_13 = {regroupV0_hi_hi_lo_lo_hi_13, regroupV0_hi_hi_lo_lo_lo_13};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo_lo_2 = {regroupV0_hi_12[2566], regroupV0_hi_12[2562]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo_hi_2 = {regroupV0_hi_12[2574], regroupV0_hi_12[2570]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo_6 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo_hi_2, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi_lo_2 = {regroupV0_hi_12[2582], regroupV0_hi_12[2578]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi_hi_2 = {regroupV0_hi_12[2590], regroupV0_hi_12[2586]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi_6 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi_hi_2, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_10 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi_6, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo_lo_2 = {regroupV0_hi_12[2598], regroupV0_hi_12[2594]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo_hi_2 = {regroupV0_hi_12[2606], regroupV0_hi_12[2602]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo_6 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo_hi_2, regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi_lo_2 = {regroupV0_hi_12[2614], regroupV0_hi_12[2610]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi_hi_2 = {regroupV0_hi_12[2622], regroupV0_hi_12[2618]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi_6 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi_hi_2, regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_10 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi_6, regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_lo_lo_13 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_10, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_10};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo_lo_2 = {regroupV0_hi_12[2630], regroupV0_hi_12[2626]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo_hi_2 = {regroupV0_hi_12[2638], regroupV0_hi_12[2634]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo_6 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo_hi_2, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi_lo_2 = {regroupV0_hi_12[2646], regroupV0_hi_12[2642]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi_hi_2 = {regroupV0_hi_12[2654], regroupV0_hi_12[2650]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi_6 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi_hi_2, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_10 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi_6, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo_lo_2 = {regroupV0_hi_12[2662], regroupV0_hi_12[2658]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo_hi_2 = {regroupV0_hi_12[2670], regroupV0_hi_12[2666]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo_6 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo_hi_2, regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi_lo_2 = {regroupV0_hi_12[2678], regroupV0_hi_12[2674]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi_hi_2 = {regroupV0_hi_12[2686], regroupV0_hi_12[2682]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi_6 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi_hi_2, regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_10 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi_6, regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_lo_hi_13 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_10, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_10};
  wire [31:0]        regroupV0_hi_hi_lo_hi_lo_lo_13 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_13, regroupV0_hi_hi_lo_hi_lo_lo_lo_13};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo_lo_2 = {regroupV0_hi_12[2694], regroupV0_hi_12[2690]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo_hi_2 = {regroupV0_hi_12[2702], regroupV0_hi_12[2698]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo_6 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo_hi_2, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi_lo_2 = {regroupV0_hi_12[2710], regroupV0_hi_12[2706]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi_hi_2 = {regroupV0_hi_12[2718], regroupV0_hi_12[2714]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi_6 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi_hi_2, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_10 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi_6, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo_lo_2 = {regroupV0_hi_12[2726], regroupV0_hi_12[2722]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo_hi_2 = {regroupV0_hi_12[2734], regroupV0_hi_12[2730]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo_6 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo_hi_2, regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi_lo_2 = {regroupV0_hi_12[2742], regroupV0_hi_12[2738]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi_hi_2 = {regroupV0_hi_12[2750], regroupV0_hi_12[2746]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi_6 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi_hi_2, regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_10 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi_6, regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_hi_lo_13 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_10, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_10};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo_lo_2 = {regroupV0_hi_12[2758], regroupV0_hi_12[2754]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo_hi_2 = {regroupV0_hi_12[2766], regroupV0_hi_12[2762]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo_6 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo_hi_2, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi_lo_2 = {regroupV0_hi_12[2774], regroupV0_hi_12[2770]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi_hi_2 = {regroupV0_hi_12[2782], regroupV0_hi_12[2778]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi_6 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi_hi_2, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_10 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi_6, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo_lo_2 = {regroupV0_hi_12[2790], regroupV0_hi_12[2786]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo_hi_2 = {regroupV0_hi_12[2798], regroupV0_hi_12[2794]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo_6 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo_hi_2, regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi_lo_2 = {regroupV0_hi_12[2806], regroupV0_hi_12[2802]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi_hi_2 = {regroupV0_hi_12[2814], regroupV0_hi_12[2810]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi_6 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi_hi_2, regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_10 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi_6, regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_hi_hi_13 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_10, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_10};
  wire [31:0]        regroupV0_hi_hi_lo_hi_lo_hi_13 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_13, regroupV0_hi_hi_lo_hi_lo_hi_lo_13};
  wire [63:0]        regroupV0_hi_hi_lo_hi_lo_13 = {regroupV0_hi_hi_lo_hi_lo_hi_13, regroupV0_hi_hi_lo_hi_lo_lo_13};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo_lo_2 = {regroupV0_hi_12[2822], regroupV0_hi_12[2818]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo_hi_2 = {regroupV0_hi_12[2830], regroupV0_hi_12[2826]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo_6 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo_hi_2, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi_lo_2 = {regroupV0_hi_12[2838], regroupV0_hi_12[2834]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi_hi_2 = {regroupV0_hi_12[2846], regroupV0_hi_12[2842]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi_6 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi_hi_2, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_10 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi_6, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo_lo_2 = {regroupV0_hi_12[2854], regroupV0_hi_12[2850]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo_hi_2 = {regroupV0_hi_12[2862], regroupV0_hi_12[2858]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo_6 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo_hi_2, regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi_lo_2 = {regroupV0_hi_12[2870], regroupV0_hi_12[2866]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi_hi_2 = {regroupV0_hi_12[2878], regroupV0_hi_12[2874]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi_6 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi_hi_2, regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_10 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi_6, regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_lo_lo_13 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_10, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_10};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo_lo_2 = {regroupV0_hi_12[2886], regroupV0_hi_12[2882]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo_hi_2 = {regroupV0_hi_12[2894], regroupV0_hi_12[2890]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo_6 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo_hi_2, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi_lo_2 = {regroupV0_hi_12[2902], regroupV0_hi_12[2898]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi_hi_2 = {regroupV0_hi_12[2910], regroupV0_hi_12[2906]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi_6 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi_hi_2, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_10 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi_6, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo_lo_2 = {regroupV0_hi_12[2918], regroupV0_hi_12[2914]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo_hi_2 = {regroupV0_hi_12[2926], regroupV0_hi_12[2922]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo_6 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo_hi_2, regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi_lo_2 = {regroupV0_hi_12[2934], regroupV0_hi_12[2930]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi_hi_2 = {regroupV0_hi_12[2942], regroupV0_hi_12[2938]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi_6 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi_hi_2, regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_10 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi_6, regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_lo_hi_13 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_10, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_10};
  wire [31:0]        regroupV0_hi_hi_lo_hi_hi_lo_13 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_13, regroupV0_hi_hi_lo_hi_hi_lo_lo_13};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo_lo_2 = {regroupV0_hi_12[2950], regroupV0_hi_12[2946]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo_hi_2 = {regroupV0_hi_12[2958], regroupV0_hi_12[2954]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo_6 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo_hi_2, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi_lo_2 = {regroupV0_hi_12[2966], regroupV0_hi_12[2962]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi_hi_2 = {regroupV0_hi_12[2974], regroupV0_hi_12[2970]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi_6 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi_hi_2, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_10 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi_6, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo_lo_2 = {regroupV0_hi_12[2982], regroupV0_hi_12[2978]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo_hi_2 = {regroupV0_hi_12[2990], regroupV0_hi_12[2986]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo_6 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo_hi_2, regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi_lo_2 = {regroupV0_hi_12[2998], regroupV0_hi_12[2994]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi_hi_2 = {regroupV0_hi_12[3006], regroupV0_hi_12[3002]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi_6 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi_hi_2, regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_10 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi_6, regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_hi_lo_13 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_10, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_10};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo_lo_2 = {regroupV0_hi_12[3014], regroupV0_hi_12[3010]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo_hi_2 = {regroupV0_hi_12[3022], regroupV0_hi_12[3018]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo_6 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo_hi_2, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi_lo_2 = {regroupV0_hi_12[3030], regroupV0_hi_12[3026]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi_hi_2 = {regroupV0_hi_12[3038], regroupV0_hi_12[3034]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi_6 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi_hi_2, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_10 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi_6, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo_lo_2 = {regroupV0_hi_12[3046], regroupV0_hi_12[3042]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo_hi_2 = {regroupV0_hi_12[3054], regroupV0_hi_12[3050]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo_6 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo_hi_2, regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi_lo_2 = {regroupV0_hi_12[3062], regroupV0_hi_12[3058]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi_hi_2 = {regroupV0_hi_12[3070], regroupV0_hi_12[3066]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi_6 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi_hi_2, regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_10 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi_6, regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_hi_hi_13 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_10, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_10};
  wire [31:0]        regroupV0_hi_hi_lo_hi_hi_hi_13 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_13, regroupV0_hi_hi_lo_hi_hi_hi_lo_13};
  wire [63:0]        regroupV0_hi_hi_lo_hi_hi_13 = {regroupV0_hi_hi_lo_hi_hi_hi_13, regroupV0_hi_hi_lo_hi_hi_lo_13};
  wire [127:0]       regroupV0_hi_hi_lo_hi_13 = {regroupV0_hi_hi_lo_hi_hi_13, regroupV0_hi_hi_lo_hi_lo_13};
  wire [255:0]       regroupV0_hi_hi_lo_13 = {regroupV0_hi_hi_lo_hi_13, regroupV0_hi_hi_lo_lo_13};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo_lo_2 = {regroupV0_hi_12[3078], regroupV0_hi_12[3074]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo_hi_2 = {regroupV0_hi_12[3086], regroupV0_hi_12[3082]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo_6 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo_hi_2, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi_lo_2 = {regroupV0_hi_12[3094], regroupV0_hi_12[3090]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi_hi_2 = {regroupV0_hi_12[3102], regroupV0_hi_12[3098]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi_6 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi_hi_2, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_10 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi_6, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo_lo_2 = {regroupV0_hi_12[3110], regroupV0_hi_12[3106]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo_hi_2 = {regroupV0_hi_12[3118], regroupV0_hi_12[3114]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo_6 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo_hi_2, regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi_lo_2 = {regroupV0_hi_12[3126], regroupV0_hi_12[3122]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi_hi_2 = {regroupV0_hi_12[3134], regroupV0_hi_12[3130]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi_6 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi_hi_2, regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_10 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi_6, regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_lo_lo_13 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_10, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_10};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo_lo_2 = {regroupV0_hi_12[3142], regroupV0_hi_12[3138]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo_hi_2 = {regroupV0_hi_12[3150], regroupV0_hi_12[3146]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo_6 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo_hi_2, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi_lo_2 = {regroupV0_hi_12[3158], regroupV0_hi_12[3154]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi_hi_2 = {regroupV0_hi_12[3166], regroupV0_hi_12[3162]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi_6 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi_hi_2, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_10 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi_6, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo_lo_2 = {regroupV0_hi_12[3174], regroupV0_hi_12[3170]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo_hi_2 = {regroupV0_hi_12[3182], regroupV0_hi_12[3178]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo_6 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo_hi_2, regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi_lo_2 = {regroupV0_hi_12[3190], regroupV0_hi_12[3186]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi_hi_2 = {regroupV0_hi_12[3198], regroupV0_hi_12[3194]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi_6 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_10 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi_6, regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_lo_hi_13 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_10, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_10};
  wire [31:0]        regroupV0_hi_hi_hi_lo_lo_lo_13 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_13, regroupV0_hi_hi_hi_lo_lo_lo_lo_13};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo_lo_2 = {regroupV0_hi_12[3206], regroupV0_hi_12[3202]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo_hi_2 = {regroupV0_hi_12[3214], regroupV0_hi_12[3210]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo_6 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo_hi_2, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi_lo_2 = {regroupV0_hi_12[3222], regroupV0_hi_12[3218]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi_hi_2 = {regroupV0_hi_12[3230], regroupV0_hi_12[3226]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi_6 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi_hi_2, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_10 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi_6, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo_lo_2 = {regroupV0_hi_12[3238], regroupV0_hi_12[3234]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo_hi_2 = {regroupV0_hi_12[3246], regroupV0_hi_12[3242]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo_6 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo_hi_2, regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi_lo_2 = {regroupV0_hi_12[3254], regroupV0_hi_12[3250]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi_hi_2 = {regroupV0_hi_12[3262], regroupV0_hi_12[3258]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi_6 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi_hi_2, regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_10 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi_6, regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_hi_lo_13 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_10, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_10};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo_lo_2 = {regroupV0_hi_12[3270], regroupV0_hi_12[3266]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo_hi_2 = {regroupV0_hi_12[3278], regroupV0_hi_12[3274]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo_6 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo_hi_2, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi_lo_2 = {regroupV0_hi_12[3286], regroupV0_hi_12[3282]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi_hi_2 = {regroupV0_hi_12[3294], regroupV0_hi_12[3290]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi_6 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi_hi_2, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_10 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi_6, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo_lo_2 = {regroupV0_hi_12[3302], regroupV0_hi_12[3298]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo_hi_2 = {regroupV0_hi_12[3310], regroupV0_hi_12[3306]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo_6 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo_hi_2, regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi_lo_2 = {regroupV0_hi_12[3318], regroupV0_hi_12[3314]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi_hi_2 = {regroupV0_hi_12[3326], regroupV0_hi_12[3322]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi_6 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_10 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi_6, regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_hi_hi_13 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_10, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_10};
  wire [31:0]        regroupV0_hi_hi_hi_lo_lo_hi_13 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_13, regroupV0_hi_hi_hi_lo_lo_hi_lo_13};
  wire [63:0]        regroupV0_hi_hi_hi_lo_lo_13 = {regroupV0_hi_hi_hi_lo_lo_hi_13, regroupV0_hi_hi_hi_lo_lo_lo_13};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo_lo_2 = {regroupV0_hi_12[3334], regroupV0_hi_12[3330]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo_hi_2 = {regroupV0_hi_12[3342], regroupV0_hi_12[3338]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo_6 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo_hi_2, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi_lo_2 = {regroupV0_hi_12[3350], regroupV0_hi_12[3346]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi_hi_2 = {regroupV0_hi_12[3358], regroupV0_hi_12[3354]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi_6 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi_hi_2, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_10 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi_6, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo_lo_2 = {regroupV0_hi_12[3366], regroupV0_hi_12[3362]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo_hi_2 = {regroupV0_hi_12[3374], regroupV0_hi_12[3370]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo_6 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo_hi_2, regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi_lo_2 = {regroupV0_hi_12[3382], regroupV0_hi_12[3378]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi_hi_2 = {regroupV0_hi_12[3390], regroupV0_hi_12[3386]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi_6 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi_hi_2, regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_10 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi_6, regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_lo_lo_13 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_10, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_10};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo_lo_2 = {regroupV0_hi_12[3398], regroupV0_hi_12[3394]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo_hi_2 = {regroupV0_hi_12[3406], regroupV0_hi_12[3402]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo_6 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo_hi_2, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi_lo_2 = {regroupV0_hi_12[3414], regroupV0_hi_12[3410]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi_hi_2 = {regroupV0_hi_12[3422], regroupV0_hi_12[3418]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi_6 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi_hi_2, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_10 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi_6, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo_lo_2 = {regroupV0_hi_12[3430], regroupV0_hi_12[3426]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo_hi_2 = {regroupV0_hi_12[3438], regroupV0_hi_12[3434]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo_6 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo_hi_2, regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi_lo_2 = {regroupV0_hi_12[3446], regroupV0_hi_12[3442]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi_hi_2 = {regroupV0_hi_12[3454], regroupV0_hi_12[3450]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi_6 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_10 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi_6, regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_lo_hi_13 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_10, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_10};
  wire [31:0]        regroupV0_hi_hi_hi_lo_hi_lo_13 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_13, regroupV0_hi_hi_hi_lo_hi_lo_lo_13};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo_lo_2 = {regroupV0_hi_12[3462], regroupV0_hi_12[3458]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo_hi_2 = {regroupV0_hi_12[3470], regroupV0_hi_12[3466]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo_6 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo_hi_2, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi_lo_2 = {regroupV0_hi_12[3478], regroupV0_hi_12[3474]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi_hi_2 = {regroupV0_hi_12[3486], regroupV0_hi_12[3482]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi_6 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi_hi_2, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_10 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi_6, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo_lo_2 = {regroupV0_hi_12[3494], regroupV0_hi_12[3490]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo_hi_2 = {regroupV0_hi_12[3502], regroupV0_hi_12[3498]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo_6 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo_hi_2, regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi_lo_2 = {regroupV0_hi_12[3510], regroupV0_hi_12[3506]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi_hi_2 = {regroupV0_hi_12[3518], regroupV0_hi_12[3514]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi_6 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi_hi_2, regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_10 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi_6, regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_hi_lo_13 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_10, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_10};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo_lo_2 = {regroupV0_hi_12[3526], regroupV0_hi_12[3522]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo_hi_2 = {regroupV0_hi_12[3534], regroupV0_hi_12[3530]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo_6 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo_hi_2, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi_lo_2 = {regroupV0_hi_12[3542], regroupV0_hi_12[3538]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi_hi_2 = {regroupV0_hi_12[3550], regroupV0_hi_12[3546]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi_6 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi_hi_2, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_10 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi_6, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo_lo_2 = {regroupV0_hi_12[3558], regroupV0_hi_12[3554]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo_hi_2 = {regroupV0_hi_12[3566], regroupV0_hi_12[3562]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo_6 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo_hi_2, regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi_lo_2 = {regroupV0_hi_12[3574], regroupV0_hi_12[3570]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi_hi_2 = {regroupV0_hi_12[3582], regroupV0_hi_12[3578]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi_6 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_10 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi_6, regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_hi_hi_13 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_10, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_10};
  wire [31:0]        regroupV0_hi_hi_hi_lo_hi_hi_13 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_13, regroupV0_hi_hi_hi_lo_hi_hi_lo_13};
  wire [63:0]        regroupV0_hi_hi_hi_lo_hi_13 = {regroupV0_hi_hi_hi_lo_hi_hi_13, regroupV0_hi_hi_hi_lo_hi_lo_13};
  wire [127:0]       regroupV0_hi_hi_hi_lo_13 = {regroupV0_hi_hi_hi_lo_hi_13, regroupV0_hi_hi_hi_lo_lo_13};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo_lo_2 = {regroupV0_hi_12[3590], regroupV0_hi_12[3586]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo_hi_2 = {regroupV0_hi_12[3598], regroupV0_hi_12[3594]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo_6 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo_hi_2, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi_lo_2 = {regroupV0_hi_12[3606], regroupV0_hi_12[3602]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi_hi_2 = {regroupV0_hi_12[3614], regroupV0_hi_12[3610]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi_6 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi_hi_2, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_10 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi_6, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo_lo_2 = {regroupV0_hi_12[3622], regroupV0_hi_12[3618]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo_hi_2 = {regroupV0_hi_12[3630], regroupV0_hi_12[3626]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo_6 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo_hi_2, regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi_lo_2 = {regroupV0_hi_12[3638], regroupV0_hi_12[3634]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi_hi_2 = {regroupV0_hi_12[3646], regroupV0_hi_12[3642]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi_6 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi_hi_2, regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_10 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi_6, regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_lo_lo_13 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_10, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_10};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo_lo_2 = {regroupV0_hi_12[3654], regroupV0_hi_12[3650]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo_hi_2 = {regroupV0_hi_12[3662], regroupV0_hi_12[3658]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo_6 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo_hi_2, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi_lo_2 = {regroupV0_hi_12[3670], regroupV0_hi_12[3666]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi_hi_2 = {regroupV0_hi_12[3678], regroupV0_hi_12[3674]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi_6 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi_hi_2, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_10 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi_6, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo_lo_2 = {regroupV0_hi_12[3686], regroupV0_hi_12[3682]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo_hi_2 = {regroupV0_hi_12[3694], regroupV0_hi_12[3690]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo_6 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo_hi_2, regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi_lo_2 = {regroupV0_hi_12[3702], regroupV0_hi_12[3698]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi_hi_2 = {regroupV0_hi_12[3710], regroupV0_hi_12[3706]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi_6 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_10 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi_6, regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_lo_hi_13 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_10, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_10};
  wire [31:0]        regroupV0_hi_hi_hi_hi_lo_lo_13 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_13, regroupV0_hi_hi_hi_hi_lo_lo_lo_13};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo_lo_2 = {regroupV0_hi_12[3718], regroupV0_hi_12[3714]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo_hi_2 = {regroupV0_hi_12[3726], regroupV0_hi_12[3722]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo_6 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo_hi_2, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi_lo_2 = {regroupV0_hi_12[3734], regroupV0_hi_12[3730]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi_hi_2 = {regroupV0_hi_12[3742], regroupV0_hi_12[3738]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi_6 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi_hi_2, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_10 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi_6, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo_lo_2 = {regroupV0_hi_12[3750], regroupV0_hi_12[3746]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo_hi_2 = {regroupV0_hi_12[3758], regroupV0_hi_12[3754]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo_6 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo_hi_2, regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi_lo_2 = {regroupV0_hi_12[3766], regroupV0_hi_12[3762]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi_hi_2 = {regroupV0_hi_12[3774], regroupV0_hi_12[3770]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi_6 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi_hi_2, regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_10 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi_6, regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_hi_lo_13 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_10, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_10};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo_lo_2 = {regroupV0_hi_12[3782], regroupV0_hi_12[3778]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo_hi_2 = {regroupV0_hi_12[3790], regroupV0_hi_12[3786]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo_6 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo_hi_2, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi_lo_2 = {regroupV0_hi_12[3798], regroupV0_hi_12[3794]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi_hi_2 = {regroupV0_hi_12[3806], regroupV0_hi_12[3802]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi_6 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi_hi_2, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_10 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi_6, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo_lo_2 = {regroupV0_hi_12[3814], regroupV0_hi_12[3810]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo_hi_2 = {regroupV0_hi_12[3822], regroupV0_hi_12[3818]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo_6 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo_hi_2, regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi_lo_2 = {regroupV0_hi_12[3830], regroupV0_hi_12[3826]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi_hi_2 = {regroupV0_hi_12[3838], regroupV0_hi_12[3834]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi_6 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_10 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi_6, regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_hi_hi_13 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_10, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_10};
  wire [31:0]        regroupV0_hi_hi_hi_hi_lo_hi_13 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_13, regroupV0_hi_hi_hi_hi_lo_hi_lo_13};
  wire [63:0]        regroupV0_hi_hi_hi_hi_lo_13 = {regroupV0_hi_hi_hi_hi_lo_hi_13, regroupV0_hi_hi_hi_hi_lo_lo_13};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo_lo_2 = {regroupV0_hi_12[3846], regroupV0_hi_12[3842]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo_hi_2 = {regroupV0_hi_12[3854], regroupV0_hi_12[3850]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo_6 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo_hi_2, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi_lo_2 = {regroupV0_hi_12[3862], regroupV0_hi_12[3858]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi_hi_2 = {regroupV0_hi_12[3870], regroupV0_hi_12[3866]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi_6 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi_hi_2, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_10 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi_6, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo_lo_2 = {regroupV0_hi_12[3878], regroupV0_hi_12[3874]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo_hi_2 = {regroupV0_hi_12[3886], regroupV0_hi_12[3882]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo_6 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo_hi_2, regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi_lo_2 = {regroupV0_hi_12[3894], regroupV0_hi_12[3890]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi_hi_2 = {regroupV0_hi_12[3902], regroupV0_hi_12[3898]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi_6 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi_hi_2, regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_10 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi_6, regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_lo_lo_13 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_10, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_10};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo_lo_2 = {regroupV0_hi_12[3910], regroupV0_hi_12[3906]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo_hi_2 = {regroupV0_hi_12[3918], regroupV0_hi_12[3914]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo_6 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo_hi_2, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi_lo_2 = {regroupV0_hi_12[3926], regroupV0_hi_12[3922]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi_hi_2 = {regroupV0_hi_12[3934], regroupV0_hi_12[3930]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi_6 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi_hi_2, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_10 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi_6, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo_lo_2 = {regroupV0_hi_12[3942], regroupV0_hi_12[3938]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo_hi_2 = {regroupV0_hi_12[3950], regroupV0_hi_12[3946]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo_6 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo_hi_2, regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi_lo_2 = {regroupV0_hi_12[3958], regroupV0_hi_12[3954]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi_hi_2 = {regroupV0_hi_12[3966], regroupV0_hi_12[3962]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi_6 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_10 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi_6, regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_lo_hi_13 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_10, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_10};
  wire [31:0]        regroupV0_hi_hi_hi_hi_hi_lo_13 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_13, regroupV0_hi_hi_hi_hi_hi_lo_lo_13};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo_lo_2 = {regroupV0_hi_12[3974], regroupV0_hi_12[3970]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo_hi_2 = {regroupV0_hi_12[3982], regroupV0_hi_12[3978]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo_6 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo_hi_2, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi_lo_2 = {regroupV0_hi_12[3990], regroupV0_hi_12[3986]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi_hi_2 = {regroupV0_hi_12[3998], regroupV0_hi_12[3994]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi_6 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi_hi_2, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_10 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi_6, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo_lo_2 = {regroupV0_hi_12[4006], regroupV0_hi_12[4002]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo_hi_2 = {regroupV0_hi_12[4014], regroupV0_hi_12[4010]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo_6 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo_hi_2, regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi_lo_2 = {regroupV0_hi_12[4022], regroupV0_hi_12[4018]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi_hi_2 = {regroupV0_hi_12[4030], regroupV0_hi_12[4026]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi_6 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi_hi_2, regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_10 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi_6, regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_hi_lo_13 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_10, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_10};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo_lo_2 = {regroupV0_hi_12[4038], regroupV0_hi_12[4034]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo_hi_2 = {regroupV0_hi_12[4046], regroupV0_hi_12[4042]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo_6 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo_hi_2, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi_lo_2 = {regroupV0_hi_12[4054], regroupV0_hi_12[4050]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi_hi_2 = {regroupV0_hi_12[4062], regroupV0_hi_12[4058]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi_6 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi_hi_2, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_10 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi_6, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo_lo_2 = {regroupV0_hi_12[4070], regroupV0_hi_12[4066]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo_hi_2 = {regroupV0_hi_12[4078], regroupV0_hi_12[4074]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo_6 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo_hi_2, regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi_lo_2 = {regroupV0_hi_12[4086], regroupV0_hi_12[4082]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi_hi_2 = {regroupV0_hi_12[4094], regroupV0_hi_12[4090]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi_6 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_10 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi_6, regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_hi_hi_13 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_10, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_10};
  wire [31:0]        regroupV0_hi_hi_hi_hi_hi_hi_13 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_13, regroupV0_hi_hi_hi_hi_hi_hi_lo_13};
  wire [63:0]        regroupV0_hi_hi_hi_hi_hi_13 = {regroupV0_hi_hi_hi_hi_hi_hi_13, regroupV0_hi_hi_hi_hi_hi_lo_13};
  wire [127:0]       regroupV0_hi_hi_hi_hi_13 = {regroupV0_hi_hi_hi_hi_hi_13, regroupV0_hi_hi_hi_hi_lo_13};
  wire [255:0]       regroupV0_hi_hi_hi_13 = {regroupV0_hi_hi_hi_hi_13, regroupV0_hi_hi_hi_lo_13};
  wire [511:0]       regroupV0_hi_hi_13 = {regroupV0_hi_hi_hi_13, regroupV0_hi_hi_lo_13};
  wire [1023:0]      regroupV0_hi_15 = {regroupV0_hi_hi_13, regroupV0_hi_lo_13};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo_lo_3 = {regroupV0_lo_12[7], regroupV0_lo_12[3]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo_hi_3 = {regroupV0_lo_12[15], regroupV0_lo_12[11]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo_7 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi_lo_3 = {regroupV0_lo_12[23], regroupV0_lo_12[19]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi_hi_3 = {regroupV0_lo_12[31], regroupV0_lo_12[27]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi_7 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi_hi_3, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_11 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_hi_7, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo_lo_3 = {regroupV0_lo_12[39], regroupV0_lo_12[35]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo_hi_3 = {regroupV0_lo_12[47], regroupV0_lo_12[43]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo_7 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo_hi_3, regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi_lo_3 = {regroupV0_lo_12[55], regroupV0_lo_12[51]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi_hi_3 = {regroupV0_lo_12[63], regroupV0_lo_12[59]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi_7 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi_hi_3, regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_11 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_hi_7, regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_lo_lo_14 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_11, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo_lo_3 = {regroupV0_lo_12[71], regroupV0_lo_12[67]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo_hi_3 = {regroupV0_lo_12[79], regroupV0_lo_12[75]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo_7 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi_lo_3 = {regroupV0_lo_12[87], regroupV0_lo_12[83]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi_hi_3 = {regroupV0_lo_12[95], regroupV0_lo_12[91]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi_7 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi_hi_3, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_11 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_hi_7, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo_lo_3 = {regroupV0_lo_12[103], regroupV0_lo_12[99]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo_hi_3 = {regroupV0_lo_12[111], regroupV0_lo_12[107]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo_7 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo_hi_3, regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi_lo_3 = {regroupV0_lo_12[119], regroupV0_lo_12[115]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi_hi_3 = {regroupV0_lo_12[127], regroupV0_lo_12[123]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi_7 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi_hi_3, regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_11 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_hi_7, regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_lo_hi_14 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_11, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_11};
  wire [31:0]        regroupV0_lo_lo_lo_lo_lo_lo_14 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_14, regroupV0_lo_lo_lo_lo_lo_lo_lo_14};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo_lo_3 = {regroupV0_lo_12[135], regroupV0_lo_12[131]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo_hi_3 = {regroupV0_lo_12[143], regroupV0_lo_12[139]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo_7 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi_lo_3 = {regroupV0_lo_12[151], regroupV0_lo_12[147]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi_hi_3 = {regroupV0_lo_12[159], regroupV0_lo_12[155]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi_7 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi_hi_3, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_11 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_hi_7, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo_lo_3 = {regroupV0_lo_12[167], regroupV0_lo_12[163]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo_hi_3 = {regroupV0_lo_12[175], regroupV0_lo_12[171]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo_7 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo_hi_3, regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi_lo_3 = {regroupV0_lo_12[183], regroupV0_lo_12[179]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi_hi_3 = {regroupV0_lo_12[191], regroupV0_lo_12[187]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi_7 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi_hi_3, regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_11 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_hi_7, regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_hi_lo_14 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_11, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo_lo_3 = {regroupV0_lo_12[199], regroupV0_lo_12[195]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo_hi_3 = {regroupV0_lo_12[207], regroupV0_lo_12[203]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo_7 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi_lo_3 = {regroupV0_lo_12[215], regroupV0_lo_12[211]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi_hi_3 = {regroupV0_lo_12[223], regroupV0_lo_12[219]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi_7 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi_hi_3, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_11 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_hi_7, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo_lo_3 = {regroupV0_lo_12[231], regroupV0_lo_12[227]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo_hi_3 = {regroupV0_lo_12[239], regroupV0_lo_12[235]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo_7 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo_hi_3, regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi_lo_3 = {regroupV0_lo_12[247], regroupV0_lo_12[243]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi_hi_3 = {regroupV0_lo_12[255], regroupV0_lo_12[251]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi_7 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi_hi_3, regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_11 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_hi_7, regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_hi_hi_14 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_11, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_11};
  wire [31:0]        regroupV0_lo_lo_lo_lo_lo_hi_14 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_14, regroupV0_lo_lo_lo_lo_lo_hi_lo_14};
  wire [63:0]        regroupV0_lo_lo_lo_lo_lo_14 = {regroupV0_lo_lo_lo_lo_lo_hi_14, regroupV0_lo_lo_lo_lo_lo_lo_14};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo_lo_3 = {regroupV0_lo_12[263], regroupV0_lo_12[259]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo_hi_3 = {regroupV0_lo_12[271], regroupV0_lo_12[267]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo_7 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi_lo_3 = {regroupV0_lo_12[279], regroupV0_lo_12[275]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi_hi_3 = {regroupV0_lo_12[287], regroupV0_lo_12[283]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi_7 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi_hi_3, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_11 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_hi_7, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo_lo_3 = {regroupV0_lo_12[295], regroupV0_lo_12[291]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo_hi_3 = {regroupV0_lo_12[303], regroupV0_lo_12[299]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo_7 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo_hi_3, regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi_lo_3 = {regroupV0_lo_12[311], regroupV0_lo_12[307]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi_hi_3 = {regroupV0_lo_12[319], regroupV0_lo_12[315]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi_7 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi_hi_3, regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_11 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_hi_7, regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_lo_lo_14 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_11, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo_lo_3 = {regroupV0_lo_12[327], regroupV0_lo_12[323]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo_hi_3 = {regroupV0_lo_12[335], regroupV0_lo_12[331]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo_7 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi_lo_3 = {regroupV0_lo_12[343], regroupV0_lo_12[339]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi_hi_3 = {regroupV0_lo_12[351], regroupV0_lo_12[347]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi_7 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi_hi_3, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_11 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_hi_7, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo_lo_3 = {regroupV0_lo_12[359], regroupV0_lo_12[355]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo_hi_3 = {regroupV0_lo_12[367], regroupV0_lo_12[363]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo_7 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo_hi_3, regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi_lo_3 = {regroupV0_lo_12[375], regroupV0_lo_12[371]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi_hi_3 = {regroupV0_lo_12[383], regroupV0_lo_12[379]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi_7 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi_hi_3, regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_11 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_hi_7, regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_lo_hi_14 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_11, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_11};
  wire [31:0]        regroupV0_lo_lo_lo_lo_hi_lo_14 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_14, regroupV0_lo_lo_lo_lo_hi_lo_lo_14};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo_lo_3 = {regroupV0_lo_12[391], regroupV0_lo_12[387]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo_hi_3 = {regroupV0_lo_12[399], regroupV0_lo_12[395]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo_7 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi_lo_3 = {regroupV0_lo_12[407], regroupV0_lo_12[403]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi_hi_3 = {regroupV0_lo_12[415], regroupV0_lo_12[411]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi_7 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi_hi_3, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_11 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_hi_7, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo_lo_3 = {regroupV0_lo_12[423], regroupV0_lo_12[419]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo_hi_3 = {regroupV0_lo_12[431], regroupV0_lo_12[427]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo_7 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo_hi_3, regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi_lo_3 = {regroupV0_lo_12[439], regroupV0_lo_12[435]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi_hi_3 = {regroupV0_lo_12[447], regroupV0_lo_12[443]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi_7 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi_hi_3, regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_11 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_hi_7, regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_hi_lo_14 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_11, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo_lo_3 = {regroupV0_lo_12[455], regroupV0_lo_12[451]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo_hi_3 = {regroupV0_lo_12[463], regroupV0_lo_12[459]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo_7 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi_lo_3 = {regroupV0_lo_12[471], regroupV0_lo_12[467]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi_hi_3 = {regroupV0_lo_12[479], regroupV0_lo_12[475]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi_7 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi_hi_3, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_11 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_hi_7, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo_lo_3 = {regroupV0_lo_12[487], regroupV0_lo_12[483]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo_hi_3 = {regroupV0_lo_12[495], regroupV0_lo_12[491]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo_7 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo_hi_3, regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi_lo_3 = {regroupV0_lo_12[503], regroupV0_lo_12[499]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi_hi_3 = {regroupV0_lo_12[511], regroupV0_lo_12[507]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi_7 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi_hi_3, regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_11 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_hi_7, regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_hi_hi_14 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_11, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_11};
  wire [31:0]        regroupV0_lo_lo_lo_lo_hi_hi_14 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_14, regroupV0_lo_lo_lo_lo_hi_hi_lo_14};
  wire [63:0]        regroupV0_lo_lo_lo_lo_hi_14 = {regroupV0_lo_lo_lo_lo_hi_hi_14, regroupV0_lo_lo_lo_lo_hi_lo_14};
  wire [127:0]       regroupV0_lo_lo_lo_lo_14 = {regroupV0_lo_lo_lo_lo_hi_14, regroupV0_lo_lo_lo_lo_lo_14};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo_lo_3 = {regroupV0_lo_12[519], regroupV0_lo_12[515]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo_hi_3 = {regroupV0_lo_12[527], regroupV0_lo_12[523]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo_7 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi_lo_3 = {regroupV0_lo_12[535], regroupV0_lo_12[531]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi_hi_3 = {regroupV0_lo_12[543], regroupV0_lo_12[539]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi_7 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi_hi_3, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_11 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_hi_7, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo_lo_3 = {regroupV0_lo_12[551], regroupV0_lo_12[547]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo_hi_3 = {regroupV0_lo_12[559], regroupV0_lo_12[555]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo_7 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo_hi_3, regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi_lo_3 = {regroupV0_lo_12[567], regroupV0_lo_12[563]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi_hi_3 = {regroupV0_lo_12[575], regroupV0_lo_12[571]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi_7 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi_hi_3, regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_11 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_hi_7, regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_lo_lo_14 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_11, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo_lo_3 = {regroupV0_lo_12[583], regroupV0_lo_12[579]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo_hi_3 = {regroupV0_lo_12[591], regroupV0_lo_12[587]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo_7 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo_hi_3, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi_lo_3 = {regroupV0_lo_12[599], regroupV0_lo_12[595]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi_hi_3 = {regroupV0_lo_12[607], regroupV0_lo_12[603]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi_7 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi_hi_3, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_11 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_hi_7, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo_lo_3 = {regroupV0_lo_12[615], regroupV0_lo_12[611]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo_hi_3 = {regroupV0_lo_12[623], regroupV0_lo_12[619]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo_7 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo_hi_3, regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi_lo_3 = {regroupV0_lo_12[631], regroupV0_lo_12[627]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi_hi_3 = {regroupV0_lo_12[639], regroupV0_lo_12[635]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi_7 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi_hi_3, regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_11 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_hi_7, regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_lo_hi_14 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_11, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_11};
  wire [31:0]        regroupV0_lo_lo_lo_hi_lo_lo_14 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_14, regroupV0_lo_lo_lo_hi_lo_lo_lo_14};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo_lo_3 = {regroupV0_lo_12[647], regroupV0_lo_12[643]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo_hi_3 = {regroupV0_lo_12[655], regroupV0_lo_12[651]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo_7 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi_lo_3 = {regroupV0_lo_12[663], regroupV0_lo_12[659]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi_hi_3 = {regroupV0_lo_12[671], regroupV0_lo_12[667]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi_7 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi_hi_3, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_11 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_hi_7, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo_lo_3 = {regroupV0_lo_12[679], regroupV0_lo_12[675]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo_hi_3 = {regroupV0_lo_12[687], regroupV0_lo_12[683]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo_7 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo_hi_3, regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi_lo_3 = {regroupV0_lo_12[695], regroupV0_lo_12[691]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi_hi_3 = {regroupV0_lo_12[703], regroupV0_lo_12[699]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi_7 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi_hi_3, regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_11 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_hi_7, regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_hi_lo_14 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_11, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo_lo_3 = {regroupV0_lo_12[711], regroupV0_lo_12[707]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo_hi_3 = {regroupV0_lo_12[719], regroupV0_lo_12[715]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo_7 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo_hi_3, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi_lo_3 = {regroupV0_lo_12[727], regroupV0_lo_12[723]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi_hi_3 = {regroupV0_lo_12[735], regroupV0_lo_12[731]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi_7 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi_hi_3, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_11 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_hi_7, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo_lo_3 = {regroupV0_lo_12[743], regroupV0_lo_12[739]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo_hi_3 = {regroupV0_lo_12[751], regroupV0_lo_12[747]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo_7 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo_hi_3, regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi_lo_3 = {regroupV0_lo_12[759], regroupV0_lo_12[755]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi_hi_3 = {regroupV0_lo_12[767], regroupV0_lo_12[763]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi_7 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi_hi_3, regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_11 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_hi_7, regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_hi_hi_14 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_11, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_11};
  wire [31:0]        regroupV0_lo_lo_lo_hi_lo_hi_14 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_14, regroupV0_lo_lo_lo_hi_lo_hi_lo_14};
  wire [63:0]        regroupV0_lo_lo_lo_hi_lo_14 = {regroupV0_lo_lo_lo_hi_lo_hi_14, regroupV0_lo_lo_lo_hi_lo_lo_14};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo_lo_3 = {regroupV0_lo_12[775], regroupV0_lo_12[771]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo_hi_3 = {regroupV0_lo_12[783], regroupV0_lo_12[779]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo_7 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi_lo_3 = {regroupV0_lo_12[791], regroupV0_lo_12[787]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi_hi_3 = {regroupV0_lo_12[799], regroupV0_lo_12[795]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi_7 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi_hi_3, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_11 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_hi_7, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo_lo_3 = {regroupV0_lo_12[807], regroupV0_lo_12[803]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo_hi_3 = {regroupV0_lo_12[815], regroupV0_lo_12[811]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo_7 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo_hi_3, regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi_lo_3 = {regroupV0_lo_12[823], regroupV0_lo_12[819]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi_hi_3 = {regroupV0_lo_12[831], regroupV0_lo_12[827]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi_7 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi_hi_3, regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_11 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_hi_7, regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_lo_lo_14 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_11, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo_lo_3 = {regroupV0_lo_12[839], regroupV0_lo_12[835]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo_hi_3 = {regroupV0_lo_12[847], regroupV0_lo_12[843]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo_7 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo_hi_3, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi_lo_3 = {regroupV0_lo_12[855], regroupV0_lo_12[851]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi_hi_3 = {regroupV0_lo_12[863], regroupV0_lo_12[859]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi_7 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi_hi_3, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_11 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_hi_7, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo_lo_3 = {regroupV0_lo_12[871], regroupV0_lo_12[867]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo_hi_3 = {regroupV0_lo_12[879], regroupV0_lo_12[875]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo_7 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo_hi_3, regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi_lo_3 = {regroupV0_lo_12[887], regroupV0_lo_12[883]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi_hi_3 = {regroupV0_lo_12[895], regroupV0_lo_12[891]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi_7 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi_hi_3, regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_11 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_hi_7, regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_lo_hi_14 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_11, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_11};
  wire [31:0]        regroupV0_lo_lo_lo_hi_hi_lo_14 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_14, regroupV0_lo_lo_lo_hi_hi_lo_lo_14};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo_lo_3 = {regroupV0_lo_12[903], regroupV0_lo_12[899]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo_hi_3 = {regroupV0_lo_12[911], regroupV0_lo_12[907]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo_7 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi_lo_3 = {regroupV0_lo_12[919], regroupV0_lo_12[915]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi_hi_3 = {regroupV0_lo_12[927], regroupV0_lo_12[923]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi_7 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi_hi_3, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_11 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_hi_7, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo_lo_3 = {regroupV0_lo_12[935], regroupV0_lo_12[931]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo_hi_3 = {regroupV0_lo_12[943], regroupV0_lo_12[939]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo_7 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo_hi_3, regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi_lo_3 = {regroupV0_lo_12[951], regroupV0_lo_12[947]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi_hi_3 = {regroupV0_lo_12[959], regroupV0_lo_12[955]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi_7 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi_hi_3, regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_11 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_hi_7, regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_hi_lo_14 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_11, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo_lo_3 = {regroupV0_lo_12[967], regroupV0_lo_12[963]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo_hi_3 = {regroupV0_lo_12[975], regroupV0_lo_12[971]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo_7 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo_hi_3, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi_lo_3 = {regroupV0_lo_12[983], regroupV0_lo_12[979]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi_hi_3 = {regroupV0_lo_12[991], regroupV0_lo_12[987]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi_7 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi_hi_3, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_11 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_hi_7, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo_lo_3 = {regroupV0_lo_12[999], regroupV0_lo_12[995]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo_hi_3 = {regroupV0_lo_12[1007], regroupV0_lo_12[1003]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo_7 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo_hi_3, regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi_lo_3 = {regroupV0_lo_12[1015], regroupV0_lo_12[1011]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi_hi_3 = {regroupV0_lo_12[1023], regroupV0_lo_12[1019]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi_7 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi_hi_3, regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_11 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_hi_7, regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_hi_hi_14 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_11, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_11};
  wire [31:0]        regroupV0_lo_lo_lo_hi_hi_hi_14 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_14, regroupV0_lo_lo_lo_hi_hi_hi_lo_14};
  wire [63:0]        regroupV0_lo_lo_lo_hi_hi_14 = {regroupV0_lo_lo_lo_hi_hi_hi_14, regroupV0_lo_lo_lo_hi_hi_lo_14};
  wire [127:0]       regroupV0_lo_lo_lo_hi_14 = {regroupV0_lo_lo_lo_hi_hi_14, regroupV0_lo_lo_lo_hi_lo_14};
  wire [255:0]       regroupV0_lo_lo_lo_14 = {regroupV0_lo_lo_lo_hi_14, regroupV0_lo_lo_lo_lo_14};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo_lo_3 = {regroupV0_lo_12[1031], regroupV0_lo_12[1027]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo_hi_3 = {regroupV0_lo_12[1039], regroupV0_lo_12[1035]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo_7 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo_hi_3, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi_lo_3 = {regroupV0_lo_12[1047], regroupV0_lo_12[1043]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi_hi_3 = {regroupV0_lo_12[1055], regroupV0_lo_12[1051]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi_7 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi_hi_3, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_11 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_hi_7, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo_lo_3 = {regroupV0_lo_12[1063], regroupV0_lo_12[1059]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo_hi_3 = {regroupV0_lo_12[1071], regroupV0_lo_12[1067]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo_7 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo_hi_3, regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi_lo_3 = {regroupV0_lo_12[1079], regroupV0_lo_12[1075]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi_hi_3 = {regroupV0_lo_12[1087], regroupV0_lo_12[1083]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi_7 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi_hi_3, regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_11 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_hi_7, regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_lo_lo_14 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_11, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo_lo_3 = {regroupV0_lo_12[1095], regroupV0_lo_12[1091]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo_hi_3 = {regroupV0_lo_12[1103], regroupV0_lo_12[1099]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo_7 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo_hi_3, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi_lo_3 = {regroupV0_lo_12[1111], regroupV0_lo_12[1107]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi_hi_3 = {regroupV0_lo_12[1119], regroupV0_lo_12[1115]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi_7 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi_hi_3, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_11 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_hi_7, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo_lo_3 = {regroupV0_lo_12[1127], regroupV0_lo_12[1123]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo_hi_3 = {regroupV0_lo_12[1135], regroupV0_lo_12[1131]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo_7 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo_hi_3, regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi_lo_3 = {regroupV0_lo_12[1143], regroupV0_lo_12[1139]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi_hi_3 = {regroupV0_lo_12[1151], regroupV0_lo_12[1147]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi_7 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi_hi_3, regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_11 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_hi_7, regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_lo_hi_14 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_11, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_11};
  wire [31:0]        regroupV0_lo_lo_hi_lo_lo_lo_14 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_14, regroupV0_lo_lo_hi_lo_lo_lo_lo_14};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo_lo_3 = {regroupV0_lo_12[1159], regroupV0_lo_12[1155]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo_hi_3 = {regroupV0_lo_12[1167], regroupV0_lo_12[1163]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo_7 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo_hi_3, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi_lo_3 = {regroupV0_lo_12[1175], regroupV0_lo_12[1171]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi_hi_3 = {regroupV0_lo_12[1183], regroupV0_lo_12[1179]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi_7 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi_hi_3, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_11 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_hi_7, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo_lo_3 = {regroupV0_lo_12[1191], regroupV0_lo_12[1187]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo_hi_3 = {regroupV0_lo_12[1199], regroupV0_lo_12[1195]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo_7 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo_hi_3, regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi_lo_3 = {regroupV0_lo_12[1207], regroupV0_lo_12[1203]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi_hi_3 = {regroupV0_lo_12[1215], regroupV0_lo_12[1211]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi_7 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi_hi_3, regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_11 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_hi_7, regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_hi_lo_14 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_11, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo_lo_3 = {regroupV0_lo_12[1223], regroupV0_lo_12[1219]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo_hi_3 = {regroupV0_lo_12[1231], regroupV0_lo_12[1227]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo_7 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo_hi_3, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi_lo_3 = {regroupV0_lo_12[1239], regroupV0_lo_12[1235]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi_hi_3 = {regroupV0_lo_12[1247], regroupV0_lo_12[1243]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi_7 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi_hi_3, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_11 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_hi_7, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo_lo_3 = {regroupV0_lo_12[1255], regroupV0_lo_12[1251]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo_hi_3 = {regroupV0_lo_12[1263], regroupV0_lo_12[1259]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo_7 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo_hi_3, regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi_lo_3 = {regroupV0_lo_12[1271], regroupV0_lo_12[1267]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi_hi_3 = {regroupV0_lo_12[1279], regroupV0_lo_12[1275]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi_7 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi_hi_3, regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_11 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_hi_7, regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_hi_hi_14 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_11, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_11};
  wire [31:0]        regroupV0_lo_lo_hi_lo_lo_hi_14 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_14, regroupV0_lo_lo_hi_lo_lo_hi_lo_14};
  wire [63:0]        regroupV0_lo_lo_hi_lo_lo_14 = {regroupV0_lo_lo_hi_lo_lo_hi_14, regroupV0_lo_lo_hi_lo_lo_lo_14};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo_lo_3 = {regroupV0_lo_12[1287], regroupV0_lo_12[1283]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo_hi_3 = {regroupV0_lo_12[1295], regroupV0_lo_12[1291]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo_7 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo_hi_3, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi_lo_3 = {regroupV0_lo_12[1303], regroupV0_lo_12[1299]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi_hi_3 = {regroupV0_lo_12[1311], regroupV0_lo_12[1307]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi_7 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi_hi_3, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_11 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_hi_7, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo_lo_3 = {regroupV0_lo_12[1319], regroupV0_lo_12[1315]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo_hi_3 = {regroupV0_lo_12[1327], regroupV0_lo_12[1323]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo_7 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo_hi_3, regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi_lo_3 = {regroupV0_lo_12[1335], regroupV0_lo_12[1331]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi_hi_3 = {regroupV0_lo_12[1343], regroupV0_lo_12[1339]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi_7 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi_hi_3, regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_11 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_hi_7, regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_lo_lo_14 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_11, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo_lo_3 = {regroupV0_lo_12[1351], regroupV0_lo_12[1347]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo_hi_3 = {regroupV0_lo_12[1359], regroupV0_lo_12[1355]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo_7 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo_hi_3, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi_lo_3 = {regroupV0_lo_12[1367], regroupV0_lo_12[1363]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi_hi_3 = {regroupV0_lo_12[1375], regroupV0_lo_12[1371]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi_7 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi_hi_3, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_11 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_hi_7, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo_lo_3 = {regroupV0_lo_12[1383], regroupV0_lo_12[1379]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo_hi_3 = {regroupV0_lo_12[1391], regroupV0_lo_12[1387]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo_7 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo_hi_3, regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi_lo_3 = {regroupV0_lo_12[1399], regroupV0_lo_12[1395]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi_hi_3 = {regroupV0_lo_12[1407], regroupV0_lo_12[1403]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi_7 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi_hi_3, regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_11 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_hi_7, regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_lo_hi_14 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_11, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_11};
  wire [31:0]        regroupV0_lo_lo_hi_lo_hi_lo_14 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_14, regroupV0_lo_lo_hi_lo_hi_lo_lo_14};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo_lo_3 = {regroupV0_lo_12[1415], regroupV0_lo_12[1411]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo_hi_3 = {regroupV0_lo_12[1423], regroupV0_lo_12[1419]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo_7 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo_hi_3, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi_lo_3 = {regroupV0_lo_12[1431], regroupV0_lo_12[1427]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi_hi_3 = {regroupV0_lo_12[1439], regroupV0_lo_12[1435]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi_7 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi_hi_3, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_11 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_hi_7, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo_lo_3 = {regroupV0_lo_12[1447], regroupV0_lo_12[1443]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo_hi_3 = {regroupV0_lo_12[1455], regroupV0_lo_12[1451]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo_7 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo_hi_3, regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi_lo_3 = {regroupV0_lo_12[1463], regroupV0_lo_12[1459]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi_hi_3 = {regroupV0_lo_12[1471], regroupV0_lo_12[1467]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi_7 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi_hi_3, regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_11 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_hi_7, regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_hi_lo_14 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_11, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo_lo_3 = {regroupV0_lo_12[1479], regroupV0_lo_12[1475]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo_hi_3 = {regroupV0_lo_12[1487], regroupV0_lo_12[1483]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo_7 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo_hi_3, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi_lo_3 = {regroupV0_lo_12[1495], regroupV0_lo_12[1491]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi_hi_3 = {regroupV0_lo_12[1503], regroupV0_lo_12[1499]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi_7 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi_hi_3, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_11 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_hi_7, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo_lo_3 = {regroupV0_lo_12[1511], regroupV0_lo_12[1507]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo_hi_3 = {regroupV0_lo_12[1519], regroupV0_lo_12[1515]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo_7 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo_hi_3, regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi_lo_3 = {regroupV0_lo_12[1527], regroupV0_lo_12[1523]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi_hi_3 = {regroupV0_lo_12[1535], regroupV0_lo_12[1531]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi_7 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi_hi_3, regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_11 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_hi_7, regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_hi_hi_14 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_11, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_11};
  wire [31:0]        regroupV0_lo_lo_hi_lo_hi_hi_14 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_14, regroupV0_lo_lo_hi_lo_hi_hi_lo_14};
  wire [63:0]        regroupV0_lo_lo_hi_lo_hi_14 = {regroupV0_lo_lo_hi_lo_hi_hi_14, regroupV0_lo_lo_hi_lo_hi_lo_14};
  wire [127:0]       regroupV0_lo_lo_hi_lo_14 = {regroupV0_lo_lo_hi_lo_hi_14, regroupV0_lo_lo_hi_lo_lo_14};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo_lo_3 = {regroupV0_lo_12[1543], regroupV0_lo_12[1539]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo_hi_3 = {regroupV0_lo_12[1551], regroupV0_lo_12[1547]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo_7 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo_hi_3, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi_lo_3 = {regroupV0_lo_12[1559], regroupV0_lo_12[1555]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi_hi_3 = {regroupV0_lo_12[1567], regroupV0_lo_12[1563]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi_7 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi_hi_3, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_11 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_hi_7, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo_lo_3 = {regroupV0_lo_12[1575], regroupV0_lo_12[1571]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo_hi_3 = {regroupV0_lo_12[1583], regroupV0_lo_12[1579]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo_7 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo_hi_3, regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi_lo_3 = {regroupV0_lo_12[1591], regroupV0_lo_12[1587]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi_hi_3 = {regroupV0_lo_12[1599], regroupV0_lo_12[1595]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi_7 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi_hi_3, regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_11 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_hi_7, regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_lo_lo_14 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_11, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo_lo_3 = {regroupV0_lo_12[1607], regroupV0_lo_12[1603]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo_hi_3 = {regroupV0_lo_12[1615], regroupV0_lo_12[1611]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo_7 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo_hi_3, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi_lo_3 = {regroupV0_lo_12[1623], regroupV0_lo_12[1619]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi_hi_3 = {regroupV0_lo_12[1631], regroupV0_lo_12[1627]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi_7 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi_hi_3, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_11 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_hi_7, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo_lo_3 = {regroupV0_lo_12[1639], regroupV0_lo_12[1635]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo_hi_3 = {regroupV0_lo_12[1647], regroupV0_lo_12[1643]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo_7 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo_hi_3, regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi_lo_3 = {regroupV0_lo_12[1655], regroupV0_lo_12[1651]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi_hi_3 = {regroupV0_lo_12[1663], regroupV0_lo_12[1659]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi_7 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi_hi_3, regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_11 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_hi_7, regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_lo_hi_14 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_11, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_11};
  wire [31:0]        regroupV0_lo_lo_hi_hi_lo_lo_14 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_14, regroupV0_lo_lo_hi_hi_lo_lo_lo_14};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo_lo_3 = {regroupV0_lo_12[1671], regroupV0_lo_12[1667]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo_hi_3 = {regroupV0_lo_12[1679], regroupV0_lo_12[1675]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo_7 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo_hi_3, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi_lo_3 = {regroupV0_lo_12[1687], regroupV0_lo_12[1683]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi_hi_3 = {regroupV0_lo_12[1695], regroupV0_lo_12[1691]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi_7 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi_hi_3, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_11 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_hi_7, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo_lo_3 = {regroupV0_lo_12[1703], regroupV0_lo_12[1699]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo_hi_3 = {regroupV0_lo_12[1711], regroupV0_lo_12[1707]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo_7 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo_hi_3, regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi_lo_3 = {regroupV0_lo_12[1719], regroupV0_lo_12[1715]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi_hi_3 = {regroupV0_lo_12[1727], regroupV0_lo_12[1723]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi_7 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi_hi_3, regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_11 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_hi_7, regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_hi_lo_14 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_11, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo_lo_3 = {regroupV0_lo_12[1735], regroupV0_lo_12[1731]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo_hi_3 = {regroupV0_lo_12[1743], regroupV0_lo_12[1739]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo_7 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo_hi_3, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi_lo_3 = {regroupV0_lo_12[1751], regroupV0_lo_12[1747]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi_hi_3 = {regroupV0_lo_12[1759], regroupV0_lo_12[1755]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi_7 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi_hi_3, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_11 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_hi_7, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo_lo_3 = {regroupV0_lo_12[1767], regroupV0_lo_12[1763]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo_hi_3 = {regroupV0_lo_12[1775], regroupV0_lo_12[1771]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo_7 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo_hi_3, regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi_lo_3 = {regroupV0_lo_12[1783], regroupV0_lo_12[1779]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi_hi_3 = {regroupV0_lo_12[1791], regroupV0_lo_12[1787]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi_7 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi_hi_3, regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_11 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_hi_7, regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_hi_hi_14 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_11, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_11};
  wire [31:0]        regroupV0_lo_lo_hi_hi_lo_hi_14 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_14, regroupV0_lo_lo_hi_hi_lo_hi_lo_14};
  wire [63:0]        regroupV0_lo_lo_hi_hi_lo_14 = {regroupV0_lo_lo_hi_hi_lo_hi_14, regroupV0_lo_lo_hi_hi_lo_lo_14};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo_lo_3 = {regroupV0_lo_12[1799], regroupV0_lo_12[1795]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo_hi_3 = {regroupV0_lo_12[1807], regroupV0_lo_12[1803]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo_7 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo_hi_3, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi_lo_3 = {regroupV0_lo_12[1815], regroupV0_lo_12[1811]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi_hi_3 = {regroupV0_lo_12[1823], regroupV0_lo_12[1819]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi_7 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi_hi_3, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_11 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_hi_7, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo_lo_3 = {regroupV0_lo_12[1831], regroupV0_lo_12[1827]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo_hi_3 = {regroupV0_lo_12[1839], regroupV0_lo_12[1835]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo_7 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo_hi_3, regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi_lo_3 = {regroupV0_lo_12[1847], regroupV0_lo_12[1843]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi_hi_3 = {regroupV0_lo_12[1855], regroupV0_lo_12[1851]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi_7 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi_hi_3, regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_11 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_hi_7, regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_lo_lo_14 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_11, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo_lo_3 = {regroupV0_lo_12[1863], regroupV0_lo_12[1859]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo_hi_3 = {regroupV0_lo_12[1871], regroupV0_lo_12[1867]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo_7 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo_hi_3, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi_lo_3 = {regroupV0_lo_12[1879], regroupV0_lo_12[1875]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi_hi_3 = {regroupV0_lo_12[1887], regroupV0_lo_12[1883]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi_7 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi_hi_3, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_11 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_hi_7, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo_lo_3 = {regroupV0_lo_12[1895], regroupV0_lo_12[1891]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo_hi_3 = {regroupV0_lo_12[1903], regroupV0_lo_12[1899]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo_7 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo_hi_3, regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi_lo_3 = {regroupV0_lo_12[1911], regroupV0_lo_12[1907]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi_hi_3 = {regroupV0_lo_12[1919], regroupV0_lo_12[1915]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi_7 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi_hi_3, regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_11 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_hi_7, regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_lo_hi_14 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_11, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_11};
  wire [31:0]        regroupV0_lo_lo_hi_hi_hi_lo_14 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_14, regroupV0_lo_lo_hi_hi_hi_lo_lo_14};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo_lo_3 = {regroupV0_lo_12[1927], regroupV0_lo_12[1923]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo_hi_3 = {regroupV0_lo_12[1935], regroupV0_lo_12[1931]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo_7 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo_hi_3, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi_lo_3 = {regroupV0_lo_12[1943], regroupV0_lo_12[1939]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi_hi_3 = {regroupV0_lo_12[1951], regroupV0_lo_12[1947]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi_7 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi_hi_3, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_11 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_hi_7, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo_lo_3 = {regroupV0_lo_12[1959], regroupV0_lo_12[1955]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo_hi_3 = {regroupV0_lo_12[1967], regroupV0_lo_12[1963]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo_7 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo_hi_3, regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi_lo_3 = {regroupV0_lo_12[1975], regroupV0_lo_12[1971]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi_hi_3 = {regroupV0_lo_12[1983], regroupV0_lo_12[1979]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi_7 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi_hi_3, regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_11 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_hi_7, regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_hi_lo_14 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_11, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo_lo_3 = {regroupV0_lo_12[1991], regroupV0_lo_12[1987]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo_hi_3 = {regroupV0_lo_12[1999], regroupV0_lo_12[1995]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo_7 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo_hi_3, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi_lo_3 = {regroupV0_lo_12[2007], regroupV0_lo_12[2003]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi_hi_3 = {regroupV0_lo_12[2015], regroupV0_lo_12[2011]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi_7 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi_hi_3, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_11 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_hi_7, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo_lo_3 = {regroupV0_lo_12[2023], regroupV0_lo_12[2019]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo_hi_3 = {regroupV0_lo_12[2031], regroupV0_lo_12[2027]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo_7 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo_hi_3, regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi_lo_3 = {regroupV0_lo_12[2039], regroupV0_lo_12[2035]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi_hi_3 = {regroupV0_lo_12[2047], regroupV0_lo_12[2043]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi_7 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi_hi_3, regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_11 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_hi_7, regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_hi_hi_14 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_11, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_11};
  wire [31:0]        regroupV0_lo_lo_hi_hi_hi_hi_14 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_14, regroupV0_lo_lo_hi_hi_hi_hi_lo_14};
  wire [63:0]        regroupV0_lo_lo_hi_hi_hi_14 = {regroupV0_lo_lo_hi_hi_hi_hi_14, regroupV0_lo_lo_hi_hi_hi_lo_14};
  wire [127:0]       regroupV0_lo_lo_hi_hi_14 = {regroupV0_lo_lo_hi_hi_hi_14, regroupV0_lo_lo_hi_hi_lo_14};
  wire [255:0]       regroupV0_lo_lo_hi_14 = {regroupV0_lo_lo_hi_hi_14, regroupV0_lo_lo_hi_lo_14};
  wire [511:0]       regroupV0_lo_lo_14 = {regroupV0_lo_lo_hi_14, regroupV0_lo_lo_lo_14};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo_lo_3 = {regroupV0_lo_12[2055], regroupV0_lo_12[2051]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo_hi_3 = {regroupV0_lo_12[2063], regroupV0_lo_12[2059]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo_7 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo_hi_3, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi_lo_3 = {regroupV0_lo_12[2071], regroupV0_lo_12[2067]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi_hi_3 = {regroupV0_lo_12[2079], regroupV0_lo_12[2075]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi_7 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi_hi_3, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_11 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_hi_7, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo_lo_3 = {regroupV0_lo_12[2087], regroupV0_lo_12[2083]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo_hi_3 = {regroupV0_lo_12[2095], regroupV0_lo_12[2091]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo_7 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo_hi_3, regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi_lo_3 = {regroupV0_lo_12[2103], regroupV0_lo_12[2099]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi_hi_3 = {regroupV0_lo_12[2111], regroupV0_lo_12[2107]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi_7 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi_hi_3, regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_11 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_hi_7, regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_lo_lo_14 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_11, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo_lo_3 = {regroupV0_lo_12[2119], regroupV0_lo_12[2115]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo_hi_3 = {regroupV0_lo_12[2127], regroupV0_lo_12[2123]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo_7 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo_hi_3, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi_lo_3 = {regroupV0_lo_12[2135], regroupV0_lo_12[2131]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi_hi_3 = {regroupV0_lo_12[2143], regroupV0_lo_12[2139]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi_7 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi_hi_3, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_11 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_hi_7, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo_lo_3 = {regroupV0_lo_12[2151], regroupV0_lo_12[2147]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo_hi_3 = {regroupV0_lo_12[2159], regroupV0_lo_12[2155]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo_7 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo_hi_3, regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi_lo_3 = {regroupV0_lo_12[2167], regroupV0_lo_12[2163]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi_hi_3 = {regroupV0_lo_12[2175], regroupV0_lo_12[2171]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi_7 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi_hi_3, regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_11 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_hi_7, regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_lo_hi_14 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_11, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_11};
  wire [31:0]        regroupV0_lo_hi_lo_lo_lo_lo_14 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_14, regroupV0_lo_hi_lo_lo_lo_lo_lo_14};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo_lo_3 = {regroupV0_lo_12[2183], regroupV0_lo_12[2179]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo_hi_3 = {regroupV0_lo_12[2191], regroupV0_lo_12[2187]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo_7 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo_hi_3, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi_lo_3 = {regroupV0_lo_12[2199], regroupV0_lo_12[2195]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi_hi_3 = {regroupV0_lo_12[2207], regroupV0_lo_12[2203]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi_7 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi_hi_3, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_11 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_hi_7, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo_lo_3 = {regroupV0_lo_12[2215], regroupV0_lo_12[2211]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo_hi_3 = {regroupV0_lo_12[2223], regroupV0_lo_12[2219]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo_7 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo_hi_3, regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi_lo_3 = {regroupV0_lo_12[2231], regroupV0_lo_12[2227]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi_hi_3 = {regroupV0_lo_12[2239], regroupV0_lo_12[2235]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi_7 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi_hi_3, regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_11 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_hi_7, regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_hi_lo_14 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_11, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo_lo_3 = {regroupV0_lo_12[2247], regroupV0_lo_12[2243]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo_hi_3 = {regroupV0_lo_12[2255], regroupV0_lo_12[2251]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo_7 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo_hi_3, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi_lo_3 = {regroupV0_lo_12[2263], regroupV0_lo_12[2259]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi_hi_3 = {regroupV0_lo_12[2271], regroupV0_lo_12[2267]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi_7 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi_hi_3, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_11 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_hi_7, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo_lo_3 = {regroupV0_lo_12[2279], regroupV0_lo_12[2275]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo_hi_3 = {regroupV0_lo_12[2287], regroupV0_lo_12[2283]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo_7 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo_hi_3, regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi_lo_3 = {regroupV0_lo_12[2295], regroupV0_lo_12[2291]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi_hi_3 = {regroupV0_lo_12[2303], regroupV0_lo_12[2299]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi_7 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi_hi_3, regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_11 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_hi_7, regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_hi_hi_14 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_11, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_11};
  wire [31:0]        regroupV0_lo_hi_lo_lo_lo_hi_14 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_14, regroupV0_lo_hi_lo_lo_lo_hi_lo_14};
  wire [63:0]        regroupV0_lo_hi_lo_lo_lo_14 = {regroupV0_lo_hi_lo_lo_lo_hi_14, regroupV0_lo_hi_lo_lo_lo_lo_14};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo_lo_3 = {regroupV0_lo_12[2311], regroupV0_lo_12[2307]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo_hi_3 = {regroupV0_lo_12[2319], regroupV0_lo_12[2315]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo_7 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo_hi_3, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi_lo_3 = {regroupV0_lo_12[2327], regroupV0_lo_12[2323]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi_hi_3 = {regroupV0_lo_12[2335], regroupV0_lo_12[2331]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi_7 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi_hi_3, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_11 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_hi_7, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo_lo_3 = {regroupV0_lo_12[2343], regroupV0_lo_12[2339]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo_hi_3 = {regroupV0_lo_12[2351], regroupV0_lo_12[2347]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo_7 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo_hi_3, regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi_lo_3 = {regroupV0_lo_12[2359], regroupV0_lo_12[2355]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi_hi_3 = {regroupV0_lo_12[2367], regroupV0_lo_12[2363]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi_7 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi_hi_3, regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_11 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_hi_7, regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_lo_lo_14 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_11, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo_lo_3 = {regroupV0_lo_12[2375], regroupV0_lo_12[2371]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo_hi_3 = {regroupV0_lo_12[2383], regroupV0_lo_12[2379]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo_7 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo_hi_3, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi_lo_3 = {regroupV0_lo_12[2391], regroupV0_lo_12[2387]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi_hi_3 = {regroupV0_lo_12[2399], regroupV0_lo_12[2395]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi_7 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi_hi_3, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_11 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_hi_7, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo_lo_3 = {regroupV0_lo_12[2407], regroupV0_lo_12[2403]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo_hi_3 = {regroupV0_lo_12[2415], regroupV0_lo_12[2411]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo_7 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo_hi_3, regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi_lo_3 = {regroupV0_lo_12[2423], regroupV0_lo_12[2419]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi_hi_3 = {regroupV0_lo_12[2431], regroupV0_lo_12[2427]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi_7 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi_hi_3, regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_11 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_hi_7, regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_lo_hi_14 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_11, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_11};
  wire [31:0]        regroupV0_lo_hi_lo_lo_hi_lo_14 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_14, regroupV0_lo_hi_lo_lo_hi_lo_lo_14};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo_lo_3 = {regroupV0_lo_12[2439], regroupV0_lo_12[2435]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo_hi_3 = {regroupV0_lo_12[2447], regroupV0_lo_12[2443]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo_7 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo_hi_3, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi_lo_3 = {regroupV0_lo_12[2455], regroupV0_lo_12[2451]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi_hi_3 = {regroupV0_lo_12[2463], regroupV0_lo_12[2459]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi_7 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi_hi_3, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_11 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_hi_7, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo_lo_3 = {regroupV0_lo_12[2471], regroupV0_lo_12[2467]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo_hi_3 = {regroupV0_lo_12[2479], regroupV0_lo_12[2475]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo_7 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo_hi_3, regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi_lo_3 = {regroupV0_lo_12[2487], regroupV0_lo_12[2483]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi_hi_3 = {regroupV0_lo_12[2495], regroupV0_lo_12[2491]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi_7 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi_hi_3, regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_11 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_hi_7, regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_hi_lo_14 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_11, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo_lo_3 = {regroupV0_lo_12[2503], regroupV0_lo_12[2499]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo_hi_3 = {regroupV0_lo_12[2511], regroupV0_lo_12[2507]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo_7 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo_hi_3, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi_lo_3 = {regroupV0_lo_12[2519], regroupV0_lo_12[2515]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi_hi_3 = {regroupV0_lo_12[2527], regroupV0_lo_12[2523]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi_7 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi_hi_3, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_11 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_hi_7, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo_lo_3 = {regroupV0_lo_12[2535], regroupV0_lo_12[2531]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo_hi_3 = {regroupV0_lo_12[2543], regroupV0_lo_12[2539]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo_7 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo_hi_3, regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi_lo_3 = {regroupV0_lo_12[2551], regroupV0_lo_12[2547]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi_hi_3 = {regroupV0_lo_12[2559], regroupV0_lo_12[2555]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi_7 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi_hi_3, regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_11 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_hi_7, regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_hi_hi_14 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_11, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_11};
  wire [31:0]        regroupV0_lo_hi_lo_lo_hi_hi_14 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_14, regroupV0_lo_hi_lo_lo_hi_hi_lo_14};
  wire [63:0]        regroupV0_lo_hi_lo_lo_hi_14 = {regroupV0_lo_hi_lo_lo_hi_hi_14, regroupV0_lo_hi_lo_lo_hi_lo_14};
  wire [127:0]       regroupV0_lo_hi_lo_lo_14 = {regroupV0_lo_hi_lo_lo_hi_14, regroupV0_lo_hi_lo_lo_lo_14};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo_lo_3 = {regroupV0_lo_12[2567], regroupV0_lo_12[2563]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo_hi_3 = {regroupV0_lo_12[2575], regroupV0_lo_12[2571]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo_7 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo_hi_3, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi_lo_3 = {regroupV0_lo_12[2583], regroupV0_lo_12[2579]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi_hi_3 = {regroupV0_lo_12[2591], regroupV0_lo_12[2587]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi_7 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi_hi_3, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_11 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_hi_7, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo_lo_3 = {regroupV0_lo_12[2599], regroupV0_lo_12[2595]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo_hi_3 = {regroupV0_lo_12[2607], regroupV0_lo_12[2603]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo_7 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo_hi_3, regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi_lo_3 = {regroupV0_lo_12[2615], regroupV0_lo_12[2611]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi_hi_3 = {regroupV0_lo_12[2623], regroupV0_lo_12[2619]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi_7 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi_hi_3, regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_11 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_hi_7, regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_lo_lo_14 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_11, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo_lo_3 = {regroupV0_lo_12[2631], regroupV0_lo_12[2627]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo_hi_3 = {regroupV0_lo_12[2639], regroupV0_lo_12[2635]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo_7 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo_hi_3, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi_lo_3 = {regroupV0_lo_12[2647], regroupV0_lo_12[2643]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi_hi_3 = {regroupV0_lo_12[2655], regroupV0_lo_12[2651]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi_7 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi_hi_3, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_11 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_hi_7, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo_lo_3 = {regroupV0_lo_12[2663], regroupV0_lo_12[2659]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo_hi_3 = {regroupV0_lo_12[2671], regroupV0_lo_12[2667]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo_7 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo_hi_3, regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi_lo_3 = {regroupV0_lo_12[2679], regroupV0_lo_12[2675]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi_hi_3 = {regroupV0_lo_12[2687], regroupV0_lo_12[2683]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi_7 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi_hi_3, regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_11 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_hi_7, regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_lo_hi_14 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_11, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_11};
  wire [31:0]        regroupV0_lo_hi_lo_hi_lo_lo_14 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_14, regroupV0_lo_hi_lo_hi_lo_lo_lo_14};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo_lo_3 = {regroupV0_lo_12[2695], regroupV0_lo_12[2691]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo_hi_3 = {regroupV0_lo_12[2703], regroupV0_lo_12[2699]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo_7 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo_hi_3, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi_lo_3 = {regroupV0_lo_12[2711], regroupV0_lo_12[2707]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi_hi_3 = {regroupV0_lo_12[2719], regroupV0_lo_12[2715]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi_7 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi_hi_3, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_11 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_hi_7, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo_lo_3 = {regroupV0_lo_12[2727], regroupV0_lo_12[2723]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo_hi_3 = {regroupV0_lo_12[2735], regroupV0_lo_12[2731]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo_7 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo_hi_3, regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi_lo_3 = {regroupV0_lo_12[2743], regroupV0_lo_12[2739]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi_hi_3 = {regroupV0_lo_12[2751], regroupV0_lo_12[2747]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi_7 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi_hi_3, regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_11 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_hi_7, regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_hi_lo_14 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_11, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo_lo_3 = {regroupV0_lo_12[2759], regroupV0_lo_12[2755]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo_hi_3 = {regroupV0_lo_12[2767], regroupV0_lo_12[2763]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo_7 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo_hi_3, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi_lo_3 = {regroupV0_lo_12[2775], regroupV0_lo_12[2771]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi_hi_3 = {regroupV0_lo_12[2783], regroupV0_lo_12[2779]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi_7 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi_hi_3, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_11 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_hi_7, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo_lo_3 = {regroupV0_lo_12[2791], regroupV0_lo_12[2787]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo_hi_3 = {regroupV0_lo_12[2799], regroupV0_lo_12[2795]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo_7 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo_hi_3, regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi_lo_3 = {regroupV0_lo_12[2807], regroupV0_lo_12[2803]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi_hi_3 = {regroupV0_lo_12[2815], regroupV0_lo_12[2811]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi_7 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi_hi_3, regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_11 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_hi_7, regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_hi_hi_14 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_11, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_11};
  wire [31:0]        regroupV0_lo_hi_lo_hi_lo_hi_14 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_14, regroupV0_lo_hi_lo_hi_lo_hi_lo_14};
  wire [63:0]        regroupV0_lo_hi_lo_hi_lo_14 = {regroupV0_lo_hi_lo_hi_lo_hi_14, regroupV0_lo_hi_lo_hi_lo_lo_14};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo_lo_3 = {regroupV0_lo_12[2823], regroupV0_lo_12[2819]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo_hi_3 = {regroupV0_lo_12[2831], regroupV0_lo_12[2827]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo_7 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo_hi_3, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi_lo_3 = {regroupV0_lo_12[2839], regroupV0_lo_12[2835]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi_hi_3 = {regroupV0_lo_12[2847], regroupV0_lo_12[2843]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi_7 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi_hi_3, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_11 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_hi_7, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo_lo_3 = {regroupV0_lo_12[2855], regroupV0_lo_12[2851]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo_hi_3 = {regroupV0_lo_12[2863], regroupV0_lo_12[2859]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo_7 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo_hi_3, regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi_lo_3 = {regroupV0_lo_12[2871], regroupV0_lo_12[2867]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi_hi_3 = {regroupV0_lo_12[2879], regroupV0_lo_12[2875]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi_7 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi_hi_3, regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_11 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_hi_7, regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_lo_lo_14 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_11, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo_lo_3 = {regroupV0_lo_12[2887], regroupV0_lo_12[2883]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo_hi_3 = {regroupV0_lo_12[2895], regroupV0_lo_12[2891]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo_7 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo_hi_3, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi_lo_3 = {regroupV0_lo_12[2903], regroupV0_lo_12[2899]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi_hi_3 = {regroupV0_lo_12[2911], regroupV0_lo_12[2907]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi_7 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi_hi_3, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_11 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_hi_7, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo_lo_3 = {regroupV0_lo_12[2919], regroupV0_lo_12[2915]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo_hi_3 = {regroupV0_lo_12[2927], regroupV0_lo_12[2923]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo_7 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo_hi_3, regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi_lo_3 = {regroupV0_lo_12[2935], regroupV0_lo_12[2931]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi_hi_3 = {regroupV0_lo_12[2943], regroupV0_lo_12[2939]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi_7 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi_hi_3, regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_11 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_hi_7, regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_lo_hi_14 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_11, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_11};
  wire [31:0]        regroupV0_lo_hi_lo_hi_hi_lo_14 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_14, regroupV0_lo_hi_lo_hi_hi_lo_lo_14};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo_lo_3 = {regroupV0_lo_12[2951], regroupV0_lo_12[2947]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo_hi_3 = {regroupV0_lo_12[2959], regroupV0_lo_12[2955]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo_7 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo_hi_3, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi_lo_3 = {regroupV0_lo_12[2967], regroupV0_lo_12[2963]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi_hi_3 = {regroupV0_lo_12[2975], regroupV0_lo_12[2971]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi_7 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi_hi_3, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_11 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_hi_7, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo_lo_3 = {regroupV0_lo_12[2983], regroupV0_lo_12[2979]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo_hi_3 = {regroupV0_lo_12[2991], regroupV0_lo_12[2987]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo_7 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo_hi_3, regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi_lo_3 = {regroupV0_lo_12[2999], regroupV0_lo_12[2995]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi_hi_3 = {regroupV0_lo_12[3007], regroupV0_lo_12[3003]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi_7 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi_hi_3, regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_11 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_hi_7, regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_hi_lo_14 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_11, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo_lo_3 = {regroupV0_lo_12[3015], regroupV0_lo_12[3011]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo_hi_3 = {regroupV0_lo_12[3023], regroupV0_lo_12[3019]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo_7 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo_hi_3, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi_lo_3 = {regroupV0_lo_12[3031], regroupV0_lo_12[3027]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi_hi_3 = {regroupV0_lo_12[3039], regroupV0_lo_12[3035]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi_7 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi_hi_3, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_11 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_hi_7, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo_lo_3 = {regroupV0_lo_12[3047], regroupV0_lo_12[3043]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo_hi_3 = {regroupV0_lo_12[3055], regroupV0_lo_12[3051]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo_7 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo_hi_3, regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi_lo_3 = {regroupV0_lo_12[3063], regroupV0_lo_12[3059]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi_hi_3 = {regroupV0_lo_12[3071], regroupV0_lo_12[3067]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi_7 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi_hi_3, regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_11 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_hi_7, regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_hi_hi_14 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_11, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_11};
  wire [31:0]        regroupV0_lo_hi_lo_hi_hi_hi_14 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_14, regroupV0_lo_hi_lo_hi_hi_hi_lo_14};
  wire [63:0]        regroupV0_lo_hi_lo_hi_hi_14 = {regroupV0_lo_hi_lo_hi_hi_hi_14, regroupV0_lo_hi_lo_hi_hi_lo_14};
  wire [127:0]       regroupV0_lo_hi_lo_hi_14 = {regroupV0_lo_hi_lo_hi_hi_14, regroupV0_lo_hi_lo_hi_lo_14};
  wire [255:0]       regroupV0_lo_hi_lo_14 = {regroupV0_lo_hi_lo_hi_14, regroupV0_lo_hi_lo_lo_14};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo_lo_3 = {regroupV0_lo_12[3079], regroupV0_lo_12[3075]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo_hi_3 = {regroupV0_lo_12[3087], regroupV0_lo_12[3083]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo_7 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo_hi_3, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi_lo_3 = {regroupV0_lo_12[3095], regroupV0_lo_12[3091]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi_hi_3 = {regroupV0_lo_12[3103], regroupV0_lo_12[3099]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi_7 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi_hi_3, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_11 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_hi_7, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo_lo_3 = {regroupV0_lo_12[3111], regroupV0_lo_12[3107]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo_hi_3 = {regroupV0_lo_12[3119], regroupV0_lo_12[3115]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo_7 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo_hi_3, regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi_lo_3 = {regroupV0_lo_12[3127], regroupV0_lo_12[3123]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi_hi_3 = {regroupV0_lo_12[3135], regroupV0_lo_12[3131]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi_7 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi_hi_3, regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_11 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_hi_7, regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_lo_lo_14 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_11, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo_lo_3 = {regroupV0_lo_12[3143], regroupV0_lo_12[3139]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo_hi_3 = {regroupV0_lo_12[3151], regroupV0_lo_12[3147]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo_7 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo_hi_3, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi_lo_3 = {regroupV0_lo_12[3159], regroupV0_lo_12[3155]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi_hi_3 = {regroupV0_lo_12[3167], regroupV0_lo_12[3163]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi_7 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi_hi_3, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_11 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_hi_7, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo_lo_3 = {regroupV0_lo_12[3175], regroupV0_lo_12[3171]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo_hi_3 = {regroupV0_lo_12[3183], regroupV0_lo_12[3179]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo_7 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo_hi_3, regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi_lo_3 = {regroupV0_lo_12[3191], regroupV0_lo_12[3187]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi_hi_3 = {regroupV0_lo_12[3199], regroupV0_lo_12[3195]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi_7 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi_hi_3, regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_11 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_hi_7, regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_lo_hi_14 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_11, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_11};
  wire [31:0]        regroupV0_lo_hi_hi_lo_lo_lo_14 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_14, regroupV0_lo_hi_hi_lo_lo_lo_lo_14};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo_lo_3 = {regroupV0_lo_12[3207], regroupV0_lo_12[3203]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo_hi_3 = {regroupV0_lo_12[3215], regroupV0_lo_12[3211]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo_7 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo_hi_3, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi_lo_3 = {regroupV0_lo_12[3223], regroupV0_lo_12[3219]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi_hi_3 = {regroupV0_lo_12[3231], regroupV0_lo_12[3227]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi_7 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi_hi_3, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_11 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_hi_7, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo_lo_3 = {regroupV0_lo_12[3239], regroupV0_lo_12[3235]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo_hi_3 = {regroupV0_lo_12[3247], regroupV0_lo_12[3243]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo_7 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo_hi_3, regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi_lo_3 = {regroupV0_lo_12[3255], regroupV0_lo_12[3251]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi_hi_3 = {regroupV0_lo_12[3263], regroupV0_lo_12[3259]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi_7 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi_hi_3, regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_11 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_hi_7, regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_hi_lo_14 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_11, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo_lo_3 = {regroupV0_lo_12[3271], regroupV0_lo_12[3267]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo_hi_3 = {regroupV0_lo_12[3279], regroupV0_lo_12[3275]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo_7 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo_hi_3, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi_lo_3 = {regroupV0_lo_12[3287], regroupV0_lo_12[3283]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi_hi_3 = {regroupV0_lo_12[3295], regroupV0_lo_12[3291]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi_7 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi_hi_3, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_11 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_hi_7, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo_lo_3 = {regroupV0_lo_12[3303], regroupV0_lo_12[3299]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo_hi_3 = {regroupV0_lo_12[3311], regroupV0_lo_12[3307]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo_7 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo_hi_3, regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi_lo_3 = {regroupV0_lo_12[3319], regroupV0_lo_12[3315]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi_hi_3 = {regroupV0_lo_12[3327], regroupV0_lo_12[3323]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi_7 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi_hi_3, regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_11 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_hi_7, regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_hi_hi_14 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_11, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_11};
  wire [31:0]        regroupV0_lo_hi_hi_lo_lo_hi_14 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_14, regroupV0_lo_hi_hi_lo_lo_hi_lo_14};
  wire [63:0]        regroupV0_lo_hi_hi_lo_lo_14 = {regroupV0_lo_hi_hi_lo_lo_hi_14, regroupV0_lo_hi_hi_lo_lo_lo_14};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo_lo_3 = {regroupV0_lo_12[3335], regroupV0_lo_12[3331]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo_hi_3 = {regroupV0_lo_12[3343], regroupV0_lo_12[3339]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo_7 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo_hi_3, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi_lo_3 = {regroupV0_lo_12[3351], regroupV0_lo_12[3347]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi_hi_3 = {regroupV0_lo_12[3359], regroupV0_lo_12[3355]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi_7 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi_hi_3, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_11 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_hi_7, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo_lo_3 = {regroupV0_lo_12[3367], regroupV0_lo_12[3363]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo_hi_3 = {regroupV0_lo_12[3375], regroupV0_lo_12[3371]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo_7 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo_hi_3, regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi_lo_3 = {regroupV0_lo_12[3383], regroupV0_lo_12[3379]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi_hi_3 = {regroupV0_lo_12[3391], regroupV0_lo_12[3387]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi_7 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi_hi_3, regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_11 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_hi_7, regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_lo_lo_14 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_11, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo_lo_3 = {regroupV0_lo_12[3399], regroupV0_lo_12[3395]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo_hi_3 = {regroupV0_lo_12[3407], regroupV0_lo_12[3403]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo_7 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo_hi_3, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi_lo_3 = {regroupV0_lo_12[3415], regroupV0_lo_12[3411]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi_hi_3 = {regroupV0_lo_12[3423], regroupV0_lo_12[3419]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi_7 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi_hi_3, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_11 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_hi_7, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo_lo_3 = {regroupV0_lo_12[3431], regroupV0_lo_12[3427]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo_hi_3 = {regroupV0_lo_12[3439], regroupV0_lo_12[3435]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo_7 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo_hi_3, regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi_lo_3 = {regroupV0_lo_12[3447], regroupV0_lo_12[3443]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi_hi_3 = {regroupV0_lo_12[3455], regroupV0_lo_12[3451]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi_7 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi_hi_3, regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_11 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_hi_7, regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_lo_hi_14 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_11, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_11};
  wire [31:0]        regroupV0_lo_hi_hi_lo_hi_lo_14 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_14, regroupV0_lo_hi_hi_lo_hi_lo_lo_14};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo_lo_3 = {regroupV0_lo_12[3463], regroupV0_lo_12[3459]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo_hi_3 = {regroupV0_lo_12[3471], regroupV0_lo_12[3467]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo_7 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo_hi_3, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi_lo_3 = {regroupV0_lo_12[3479], regroupV0_lo_12[3475]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi_hi_3 = {regroupV0_lo_12[3487], regroupV0_lo_12[3483]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi_7 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi_hi_3, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_11 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_hi_7, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo_lo_3 = {regroupV0_lo_12[3495], regroupV0_lo_12[3491]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo_hi_3 = {regroupV0_lo_12[3503], regroupV0_lo_12[3499]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo_7 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo_hi_3, regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi_lo_3 = {regroupV0_lo_12[3511], regroupV0_lo_12[3507]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi_hi_3 = {regroupV0_lo_12[3519], regroupV0_lo_12[3515]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi_7 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi_hi_3, regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_11 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_hi_7, regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_hi_lo_14 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_11, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo_lo_3 = {regroupV0_lo_12[3527], regroupV0_lo_12[3523]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo_hi_3 = {regroupV0_lo_12[3535], regroupV0_lo_12[3531]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo_7 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo_hi_3, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi_lo_3 = {regroupV0_lo_12[3543], regroupV0_lo_12[3539]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi_hi_3 = {regroupV0_lo_12[3551], regroupV0_lo_12[3547]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi_7 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi_hi_3, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_11 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_hi_7, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo_lo_3 = {regroupV0_lo_12[3559], regroupV0_lo_12[3555]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo_hi_3 = {regroupV0_lo_12[3567], regroupV0_lo_12[3563]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo_7 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo_hi_3, regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi_lo_3 = {regroupV0_lo_12[3575], regroupV0_lo_12[3571]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi_hi_3 = {regroupV0_lo_12[3583], regroupV0_lo_12[3579]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi_7 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi_hi_3, regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_11 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_hi_7, regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_hi_hi_14 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_11, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_11};
  wire [31:0]        regroupV0_lo_hi_hi_lo_hi_hi_14 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_14, regroupV0_lo_hi_hi_lo_hi_hi_lo_14};
  wire [63:0]        regroupV0_lo_hi_hi_lo_hi_14 = {regroupV0_lo_hi_hi_lo_hi_hi_14, regroupV0_lo_hi_hi_lo_hi_lo_14};
  wire [127:0]       regroupV0_lo_hi_hi_lo_14 = {regroupV0_lo_hi_hi_lo_hi_14, regroupV0_lo_hi_hi_lo_lo_14};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo_lo_3 = {regroupV0_lo_12[3591], regroupV0_lo_12[3587]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo_hi_3 = {regroupV0_lo_12[3599], regroupV0_lo_12[3595]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo_7 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo_hi_3, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi_lo_3 = {regroupV0_lo_12[3607], regroupV0_lo_12[3603]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi_hi_3 = {regroupV0_lo_12[3615], regroupV0_lo_12[3611]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi_7 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi_hi_3, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_11 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_hi_7, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo_lo_3 = {regroupV0_lo_12[3623], regroupV0_lo_12[3619]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo_hi_3 = {regroupV0_lo_12[3631], regroupV0_lo_12[3627]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo_7 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo_hi_3, regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi_lo_3 = {regroupV0_lo_12[3639], regroupV0_lo_12[3635]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi_hi_3 = {regroupV0_lo_12[3647], regroupV0_lo_12[3643]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi_7 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi_hi_3, regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_11 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_hi_7, regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_lo_lo_14 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_11, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo_lo_3 = {regroupV0_lo_12[3655], regroupV0_lo_12[3651]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo_hi_3 = {regroupV0_lo_12[3663], regroupV0_lo_12[3659]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo_7 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo_hi_3, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi_lo_3 = {regroupV0_lo_12[3671], regroupV0_lo_12[3667]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi_hi_3 = {regroupV0_lo_12[3679], regroupV0_lo_12[3675]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi_7 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi_hi_3, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_11 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_hi_7, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo_lo_3 = {regroupV0_lo_12[3687], regroupV0_lo_12[3683]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo_hi_3 = {regroupV0_lo_12[3695], regroupV0_lo_12[3691]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo_7 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo_hi_3, regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi_lo_3 = {regroupV0_lo_12[3703], regroupV0_lo_12[3699]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi_hi_3 = {regroupV0_lo_12[3711], regroupV0_lo_12[3707]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi_7 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi_hi_3, regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_11 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_hi_7, regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_lo_hi_14 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_11, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_11};
  wire [31:0]        regroupV0_lo_hi_hi_hi_lo_lo_14 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_14, regroupV0_lo_hi_hi_hi_lo_lo_lo_14};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo_lo_3 = {regroupV0_lo_12[3719], regroupV0_lo_12[3715]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo_hi_3 = {regroupV0_lo_12[3727], regroupV0_lo_12[3723]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo_7 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo_hi_3, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi_lo_3 = {regroupV0_lo_12[3735], regroupV0_lo_12[3731]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi_hi_3 = {regroupV0_lo_12[3743], regroupV0_lo_12[3739]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi_7 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi_hi_3, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_11 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_hi_7, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo_lo_3 = {regroupV0_lo_12[3751], regroupV0_lo_12[3747]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo_hi_3 = {regroupV0_lo_12[3759], regroupV0_lo_12[3755]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo_7 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo_hi_3, regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi_lo_3 = {regroupV0_lo_12[3767], regroupV0_lo_12[3763]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi_hi_3 = {regroupV0_lo_12[3775], regroupV0_lo_12[3771]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi_7 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi_hi_3, regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_11 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_hi_7, regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_hi_lo_14 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_11, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo_lo_3 = {regroupV0_lo_12[3783], regroupV0_lo_12[3779]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo_hi_3 = {regroupV0_lo_12[3791], regroupV0_lo_12[3787]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo_7 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo_hi_3, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi_lo_3 = {regroupV0_lo_12[3799], regroupV0_lo_12[3795]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi_hi_3 = {regroupV0_lo_12[3807], regroupV0_lo_12[3803]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi_7 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi_hi_3, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_11 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_hi_7, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo_lo_3 = {regroupV0_lo_12[3815], regroupV0_lo_12[3811]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo_hi_3 = {regroupV0_lo_12[3823], regroupV0_lo_12[3819]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo_7 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo_hi_3, regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi_lo_3 = {regroupV0_lo_12[3831], regroupV0_lo_12[3827]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi_hi_3 = {regroupV0_lo_12[3839], regroupV0_lo_12[3835]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi_7 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi_hi_3, regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_11 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_hi_7, regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_hi_hi_14 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_11, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_11};
  wire [31:0]        regroupV0_lo_hi_hi_hi_lo_hi_14 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_14, regroupV0_lo_hi_hi_hi_lo_hi_lo_14};
  wire [63:0]        regroupV0_lo_hi_hi_hi_lo_14 = {regroupV0_lo_hi_hi_hi_lo_hi_14, regroupV0_lo_hi_hi_hi_lo_lo_14};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo_lo_3 = {regroupV0_lo_12[3847], regroupV0_lo_12[3843]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo_hi_3 = {regroupV0_lo_12[3855], regroupV0_lo_12[3851]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo_7 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo_hi_3, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi_lo_3 = {regroupV0_lo_12[3863], regroupV0_lo_12[3859]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi_hi_3 = {regroupV0_lo_12[3871], regroupV0_lo_12[3867]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi_7 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi_hi_3, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_11 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_hi_7, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo_lo_3 = {regroupV0_lo_12[3879], regroupV0_lo_12[3875]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo_hi_3 = {regroupV0_lo_12[3887], regroupV0_lo_12[3883]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo_7 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo_hi_3, regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi_lo_3 = {regroupV0_lo_12[3895], regroupV0_lo_12[3891]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi_hi_3 = {regroupV0_lo_12[3903], regroupV0_lo_12[3899]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi_7 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi_hi_3, regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_11 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_hi_7, regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_lo_lo_14 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_11, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo_lo_3 = {regroupV0_lo_12[3911], regroupV0_lo_12[3907]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo_hi_3 = {regroupV0_lo_12[3919], regroupV0_lo_12[3915]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo_7 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo_hi_3, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi_lo_3 = {regroupV0_lo_12[3927], regroupV0_lo_12[3923]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi_hi_3 = {regroupV0_lo_12[3935], regroupV0_lo_12[3931]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi_7 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi_hi_3, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_11 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_hi_7, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo_lo_3 = {regroupV0_lo_12[3943], regroupV0_lo_12[3939]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo_hi_3 = {regroupV0_lo_12[3951], regroupV0_lo_12[3947]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo_7 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo_hi_3, regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi_lo_3 = {regroupV0_lo_12[3959], regroupV0_lo_12[3955]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi_hi_3 = {regroupV0_lo_12[3967], regroupV0_lo_12[3963]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi_7 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi_hi_3, regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_11 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_hi_7, regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_lo_hi_14 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_11, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_11};
  wire [31:0]        regroupV0_lo_hi_hi_hi_hi_lo_14 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_14, regroupV0_lo_hi_hi_hi_hi_lo_lo_14};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo_lo_3 = {regroupV0_lo_12[3975], regroupV0_lo_12[3971]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo_hi_3 = {regroupV0_lo_12[3983], regroupV0_lo_12[3979]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo_7 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo_hi_3, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi_lo_3 = {regroupV0_lo_12[3991], regroupV0_lo_12[3987]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi_hi_3 = {regroupV0_lo_12[3999], regroupV0_lo_12[3995]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi_7 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi_hi_3, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_11 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_hi_7, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo_lo_3 = {regroupV0_lo_12[4007], regroupV0_lo_12[4003]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo_hi_3 = {regroupV0_lo_12[4015], regroupV0_lo_12[4011]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo_7 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo_hi_3, regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi_lo_3 = {regroupV0_lo_12[4023], regroupV0_lo_12[4019]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi_hi_3 = {regroupV0_lo_12[4031], regroupV0_lo_12[4027]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi_7 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi_hi_3, regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_11 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_hi_7, regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_hi_lo_14 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_11, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo_lo_3 = {regroupV0_lo_12[4039], regroupV0_lo_12[4035]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo_hi_3 = {regroupV0_lo_12[4047], regroupV0_lo_12[4043]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo_7 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo_hi_3, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi_lo_3 = {regroupV0_lo_12[4055], regroupV0_lo_12[4051]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi_hi_3 = {regroupV0_lo_12[4063], regroupV0_lo_12[4059]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi_7 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi_hi_3, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_11 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_hi_7, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo_lo_3 = {regroupV0_lo_12[4071], regroupV0_lo_12[4067]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo_hi_3 = {regroupV0_lo_12[4079], regroupV0_lo_12[4075]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo_7 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo_hi_3, regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi_lo_3 = {regroupV0_lo_12[4087], regroupV0_lo_12[4083]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi_hi_3 = {regroupV0_lo_12[4095], regroupV0_lo_12[4091]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi_7 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi_hi_3, regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_11 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_hi_7, regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_hi_hi_14 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_11, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_11};
  wire [31:0]        regroupV0_lo_hi_hi_hi_hi_hi_14 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_14, regroupV0_lo_hi_hi_hi_hi_hi_lo_14};
  wire [63:0]        regroupV0_lo_hi_hi_hi_hi_14 = {regroupV0_lo_hi_hi_hi_hi_hi_14, regroupV0_lo_hi_hi_hi_hi_lo_14};
  wire [127:0]       regroupV0_lo_hi_hi_hi_14 = {regroupV0_lo_hi_hi_hi_hi_14, regroupV0_lo_hi_hi_hi_lo_14};
  wire [255:0]       regroupV0_lo_hi_hi_14 = {regroupV0_lo_hi_hi_hi_14, regroupV0_lo_hi_hi_lo_14};
  wire [511:0]       regroupV0_lo_hi_14 = {regroupV0_lo_hi_hi_14, regroupV0_lo_hi_lo_14};
  wire [1023:0]      regroupV0_lo_16 = {regroupV0_lo_hi_14, regroupV0_lo_lo_14};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo_lo_3 = {regroupV0_hi_12[7], regroupV0_hi_12[3]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo_hi_3 = {regroupV0_hi_12[15], regroupV0_hi_12[11]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo_7 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi_lo_3 = {regroupV0_hi_12[23], regroupV0_hi_12[19]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi_hi_3 = {regroupV0_hi_12[31], regroupV0_hi_12[27]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi_7 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi_hi_3, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_11 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_hi_7, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo_lo_3 = {regroupV0_hi_12[39], regroupV0_hi_12[35]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo_hi_3 = {regroupV0_hi_12[47], regroupV0_hi_12[43]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo_7 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo_hi_3, regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi_lo_3 = {regroupV0_hi_12[55], regroupV0_hi_12[51]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi_hi_3 = {regroupV0_hi_12[63], regroupV0_hi_12[59]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi_7 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi_hi_3, regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_11 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_hi_7, regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_lo_lo_14 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_11, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo_lo_3 = {regroupV0_hi_12[71], regroupV0_hi_12[67]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo_hi_3 = {regroupV0_hi_12[79], regroupV0_hi_12[75]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo_7 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi_lo_3 = {regroupV0_hi_12[87], regroupV0_hi_12[83]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi_hi_3 = {regroupV0_hi_12[95], regroupV0_hi_12[91]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi_7 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi_hi_3, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_11 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_hi_7, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo_lo_3 = {regroupV0_hi_12[103], regroupV0_hi_12[99]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo_hi_3 = {regroupV0_hi_12[111], regroupV0_hi_12[107]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo_7 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo_hi_3, regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi_lo_3 = {regroupV0_hi_12[119], regroupV0_hi_12[115]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi_hi_3 = {regroupV0_hi_12[127], regroupV0_hi_12[123]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi_7 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi_hi_3, regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_11 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_hi_7, regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_lo_hi_14 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_11, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_11};
  wire [31:0]        regroupV0_hi_lo_lo_lo_lo_lo_14 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_14, regroupV0_hi_lo_lo_lo_lo_lo_lo_14};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo_lo_3 = {regroupV0_hi_12[135], regroupV0_hi_12[131]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo_hi_3 = {regroupV0_hi_12[143], regroupV0_hi_12[139]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo_7 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi_lo_3 = {regroupV0_hi_12[151], regroupV0_hi_12[147]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi_hi_3 = {regroupV0_hi_12[159], regroupV0_hi_12[155]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi_7 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi_hi_3, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_11 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_hi_7, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo_lo_3 = {regroupV0_hi_12[167], regroupV0_hi_12[163]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo_hi_3 = {regroupV0_hi_12[175], regroupV0_hi_12[171]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo_7 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo_hi_3, regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi_lo_3 = {regroupV0_hi_12[183], regroupV0_hi_12[179]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi_hi_3 = {regroupV0_hi_12[191], regroupV0_hi_12[187]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi_7 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi_hi_3, regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_11 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_hi_7, regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_hi_lo_14 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_11, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo_lo_3 = {regroupV0_hi_12[199], regroupV0_hi_12[195]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo_hi_3 = {regroupV0_hi_12[207], regroupV0_hi_12[203]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo_7 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi_lo_3 = {regroupV0_hi_12[215], regroupV0_hi_12[211]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi_hi_3 = {regroupV0_hi_12[223], regroupV0_hi_12[219]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi_7 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi_hi_3, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_11 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_hi_7, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo_lo_3 = {regroupV0_hi_12[231], regroupV0_hi_12[227]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo_hi_3 = {regroupV0_hi_12[239], regroupV0_hi_12[235]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo_7 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo_hi_3, regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi_lo_3 = {regroupV0_hi_12[247], regroupV0_hi_12[243]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi_hi_3 = {regroupV0_hi_12[255], regroupV0_hi_12[251]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi_7 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi_hi_3, regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_11 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_hi_7, regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_hi_hi_14 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_11, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_11};
  wire [31:0]        regroupV0_hi_lo_lo_lo_lo_hi_14 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_14, regroupV0_hi_lo_lo_lo_lo_hi_lo_14};
  wire [63:0]        regroupV0_hi_lo_lo_lo_lo_14 = {regroupV0_hi_lo_lo_lo_lo_hi_14, regroupV0_hi_lo_lo_lo_lo_lo_14};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo_lo_3 = {regroupV0_hi_12[263], regroupV0_hi_12[259]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo_hi_3 = {regroupV0_hi_12[271], regroupV0_hi_12[267]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo_7 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi_lo_3 = {regroupV0_hi_12[279], regroupV0_hi_12[275]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi_hi_3 = {regroupV0_hi_12[287], regroupV0_hi_12[283]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi_7 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi_hi_3, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_11 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_hi_7, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo_lo_3 = {regroupV0_hi_12[295], regroupV0_hi_12[291]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo_hi_3 = {regroupV0_hi_12[303], regroupV0_hi_12[299]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo_7 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo_hi_3, regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi_lo_3 = {regroupV0_hi_12[311], regroupV0_hi_12[307]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi_hi_3 = {regroupV0_hi_12[319], regroupV0_hi_12[315]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi_7 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi_hi_3, regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_11 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_hi_7, regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_lo_lo_14 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_11, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo_lo_3 = {regroupV0_hi_12[327], regroupV0_hi_12[323]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo_hi_3 = {regroupV0_hi_12[335], regroupV0_hi_12[331]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo_7 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi_lo_3 = {regroupV0_hi_12[343], regroupV0_hi_12[339]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi_hi_3 = {regroupV0_hi_12[351], regroupV0_hi_12[347]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi_7 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi_hi_3, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_11 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_hi_7, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo_lo_3 = {regroupV0_hi_12[359], regroupV0_hi_12[355]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo_hi_3 = {regroupV0_hi_12[367], regroupV0_hi_12[363]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo_7 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo_hi_3, regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi_lo_3 = {regroupV0_hi_12[375], regroupV0_hi_12[371]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi_hi_3 = {regroupV0_hi_12[383], regroupV0_hi_12[379]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi_7 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi_hi_3, regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_11 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_hi_7, regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_lo_hi_14 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_11, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_11};
  wire [31:0]        regroupV0_hi_lo_lo_lo_hi_lo_14 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_14, regroupV0_hi_lo_lo_lo_hi_lo_lo_14};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo_lo_3 = {regroupV0_hi_12[391], regroupV0_hi_12[387]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo_hi_3 = {regroupV0_hi_12[399], regroupV0_hi_12[395]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo_7 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi_lo_3 = {regroupV0_hi_12[407], regroupV0_hi_12[403]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi_hi_3 = {regroupV0_hi_12[415], regroupV0_hi_12[411]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi_7 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi_hi_3, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_11 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_hi_7, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo_lo_3 = {regroupV0_hi_12[423], regroupV0_hi_12[419]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo_hi_3 = {regroupV0_hi_12[431], regroupV0_hi_12[427]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo_7 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo_hi_3, regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi_lo_3 = {regroupV0_hi_12[439], regroupV0_hi_12[435]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi_hi_3 = {regroupV0_hi_12[447], regroupV0_hi_12[443]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi_7 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi_hi_3, regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_11 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_hi_7, regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_hi_lo_14 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_11, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo_lo_3 = {regroupV0_hi_12[455], regroupV0_hi_12[451]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo_hi_3 = {regroupV0_hi_12[463], regroupV0_hi_12[459]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo_7 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi_lo_3 = {regroupV0_hi_12[471], regroupV0_hi_12[467]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi_hi_3 = {regroupV0_hi_12[479], regroupV0_hi_12[475]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi_7 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi_hi_3, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_11 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_hi_7, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo_lo_3 = {regroupV0_hi_12[487], regroupV0_hi_12[483]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo_hi_3 = {regroupV0_hi_12[495], regroupV0_hi_12[491]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo_7 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo_hi_3, regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi_lo_3 = {regroupV0_hi_12[503], regroupV0_hi_12[499]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi_hi_3 = {regroupV0_hi_12[511], regroupV0_hi_12[507]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi_7 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi_hi_3, regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_11 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_hi_7, regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_hi_hi_14 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_11, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_11};
  wire [31:0]        regroupV0_hi_lo_lo_lo_hi_hi_14 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_14, regroupV0_hi_lo_lo_lo_hi_hi_lo_14};
  wire [63:0]        regroupV0_hi_lo_lo_lo_hi_14 = {regroupV0_hi_lo_lo_lo_hi_hi_14, regroupV0_hi_lo_lo_lo_hi_lo_14};
  wire [127:0]       regroupV0_hi_lo_lo_lo_14 = {regroupV0_hi_lo_lo_lo_hi_14, regroupV0_hi_lo_lo_lo_lo_14};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo_lo_3 = {regroupV0_hi_12[519], regroupV0_hi_12[515]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo_hi_3 = {regroupV0_hi_12[527], regroupV0_hi_12[523]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo_7 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo_hi_3, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi_lo_3 = {regroupV0_hi_12[535], regroupV0_hi_12[531]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi_hi_3 = {regroupV0_hi_12[543], regroupV0_hi_12[539]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi_7 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi_hi_3, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_11 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_hi_7, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo_lo_3 = {regroupV0_hi_12[551], regroupV0_hi_12[547]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo_hi_3 = {regroupV0_hi_12[559], regroupV0_hi_12[555]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo_7 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo_hi_3, regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi_lo_3 = {regroupV0_hi_12[567], regroupV0_hi_12[563]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi_hi_3 = {regroupV0_hi_12[575], regroupV0_hi_12[571]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi_7 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi_hi_3, regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_11 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_hi_7, regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_lo_lo_14 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_11, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo_lo_3 = {regroupV0_hi_12[583], regroupV0_hi_12[579]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo_hi_3 = {regroupV0_hi_12[591], regroupV0_hi_12[587]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo_7 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo_hi_3, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi_lo_3 = {regroupV0_hi_12[599], regroupV0_hi_12[595]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi_hi_3 = {regroupV0_hi_12[607], regroupV0_hi_12[603]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi_7 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi_hi_3, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_11 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_hi_7, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo_lo_3 = {regroupV0_hi_12[615], regroupV0_hi_12[611]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo_hi_3 = {regroupV0_hi_12[623], regroupV0_hi_12[619]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo_7 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo_hi_3, regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi_lo_3 = {regroupV0_hi_12[631], regroupV0_hi_12[627]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi_hi_3 = {regroupV0_hi_12[639], regroupV0_hi_12[635]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi_7 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi_hi_3, regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_11 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_hi_7, regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_lo_hi_14 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_11, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_11};
  wire [31:0]        regroupV0_hi_lo_lo_hi_lo_lo_14 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_14, regroupV0_hi_lo_lo_hi_lo_lo_lo_14};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo_lo_3 = {regroupV0_hi_12[647], regroupV0_hi_12[643]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo_hi_3 = {regroupV0_hi_12[655], regroupV0_hi_12[651]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo_7 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo_hi_3, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi_lo_3 = {regroupV0_hi_12[663], regroupV0_hi_12[659]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi_hi_3 = {regroupV0_hi_12[671], regroupV0_hi_12[667]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi_7 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi_hi_3, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_11 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_hi_7, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo_lo_3 = {regroupV0_hi_12[679], regroupV0_hi_12[675]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo_hi_3 = {regroupV0_hi_12[687], regroupV0_hi_12[683]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo_7 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo_hi_3, regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi_lo_3 = {regroupV0_hi_12[695], regroupV0_hi_12[691]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi_hi_3 = {regroupV0_hi_12[703], regroupV0_hi_12[699]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi_7 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi_hi_3, regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_11 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_hi_7, regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_hi_lo_14 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_11, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo_lo_3 = {regroupV0_hi_12[711], regroupV0_hi_12[707]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo_hi_3 = {regroupV0_hi_12[719], regroupV0_hi_12[715]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo_7 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo_hi_3, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi_lo_3 = {regroupV0_hi_12[727], regroupV0_hi_12[723]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi_hi_3 = {regroupV0_hi_12[735], regroupV0_hi_12[731]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi_7 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi_hi_3, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_11 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_hi_7, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo_lo_3 = {regroupV0_hi_12[743], regroupV0_hi_12[739]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo_hi_3 = {regroupV0_hi_12[751], regroupV0_hi_12[747]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo_7 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo_hi_3, regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi_lo_3 = {regroupV0_hi_12[759], regroupV0_hi_12[755]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi_hi_3 = {regroupV0_hi_12[767], regroupV0_hi_12[763]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi_7 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi_hi_3, regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_11 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_hi_7, regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_hi_hi_14 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_11, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_11};
  wire [31:0]        regroupV0_hi_lo_lo_hi_lo_hi_14 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_14, regroupV0_hi_lo_lo_hi_lo_hi_lo_14};
  wire [63:0]        regroupV0_hi_lo_lo_hi_lo_14 = {regroupV0_hi_lo_lo_hi_lo_hi_14, regroupV0_hi_lo_lo_hi_lo_lo_14};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo_lo_3 = {regroupV0_hi_12[775], regroupV0_hi_12[771]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo_hi_3 = {regroupV0_hi_12[783], regroupV0_hi_12[779]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo_7 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo_hi_3, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi_lo_3 = {regroupV0_hi_12[791], regroupV0_hi_12[787]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi_hi_3 = {regroupV0_hi_12[799], regroupV0_hi_12[795]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi_7 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi_hi_3, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_11 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_hi_7, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo_lo_3 = {regroupV0_hi_12[807], regroupV0_hi_12[803]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo_hi_3 = {regroupV0_hi_12[815], regroupV0_hi_12[811]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo_7 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo_hi_3, regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi_lo_3 = {regroupV0_hi_12[823], regroupV0_hi_12[819]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi_hi_3 = {regroupV0_hi_12[831], regroupV0_hi_12[827]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi_7 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi_hi_3, regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_11 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_hi_7, regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_lo_lo_14 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_11, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo_lo_3 = {regroupV0_hi_12[839], regroupV0_hi_12[835]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo_hi_3 = {regroupV0_hi_12[847], regroupV0_hi_12[843]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo_7 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo_hi_3, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi_lo_3 = {regroupV0_hi_12[855], regroupV0_hi_12[851]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi_hi_3 = {regroupV0_hi_12[863], regroupV0_hi_12[859]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi_7 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi_hi_3, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_11 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_hi_7, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo_lo_3 = {regroupV0_hi_12[871], regroupV0_hi_12[867]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo_hi_3 = {regroupV0_hi_12[879], regroupV0_hi_12[875]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo_7 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo_hi_3, regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi_lo_3 = {regroupV0_hi_12[887], regroupV0_hi_12[883]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi_hi_3 = {regroupV0_hi_12[895], regroupV0_hi_12[891]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi_7 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi_hi_3, regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_11 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_hi_7, regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_lo_hi_14 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_11, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_11};
  wire [31:0]        regroupV0_hi_lo_lo_hi_hi_lo_14 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_14, regroupV0_hi_lo_lo_hi_hi_lo_lo_14};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo_lo_3 = {regroupV0_hi_12[903], regroupV0_hi_12[899]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo_hi_3 = {regroupV0_hi_12[911], regroupV0_hi_12[907]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo_7 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo_hi_3, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi_lo_3 = {regroupV0_hi_12[919], regroupV0_hi_12[915]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi_hi_3 = {regroupV0_hi_12[927], regroupV0_hi_12[923]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi_7 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi_hi_3, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_11 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_hi_7, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo_lo_3 = {regroupV0_hi_12[935], regroupV0_hi_12[931]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo_hi_3 = {regroupV0_hi_12[943], regroupV0_hi_12[939]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo_7 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo_hi_3, regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi_lo_3 = {regroupV0_hi_12[951], regroupV0_hi_12[947]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi_hi_3 = {regroupV0_hi_12[959], regroupV0_hi_12[955]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi_7 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi_hi_3, regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_11 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_hi_7, regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_hi_lo_14 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_11, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo_lo_3 = {regroupV0_hi_12[967], regroupV0_hi_12[963]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo_hi_3 = {regroupV0_hi_12[975], regroupV0_hi_12[971]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo_7 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo_hi_3, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi_lo_3 = {regroupV0_hi_12[983], regroupV0_hi_12[979]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi_hi_3 = {regroupV0_hi_12[991], regroupV0_hi_12[987]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi_7 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi_hi_3, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_11 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_hi_7, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo_lo_3 = {regroupV0_hi_12[999], regroupV0_hi_12[995]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo_hi_3 = {regroupV0_hi_12[1007], regroupV0_hi_12[1003]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo_7 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo_hi_3, regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi_lo_3 = {regroupV0_hi_12[1015], regroupV0_hi_12[1011]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi_hi_3 = {regroupV0_hi_12[1023], regroupV0_hi_12[1019]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi_7 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi_hi_3, regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_11 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_hi_7, regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_hi_hi_14 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_11, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_11};
  wire [31:0]        regroupV0_hi_lo_lo_hi_hi_hi_14 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_14, regroupV0_hi_lo_lo_hi_hi_hi_lo_14};
  wire [63:0]        regroupV0_hi_lo_lo_hi_hi_14 = {regroupV0_hi_lo_lo_hi_hi_hi_14, regroupV0_hi_lo_lo_hi_hi_lo_14};
  wire [127:0]       regroupV0_hi_lo_lo_hi_14 = {regroupV0_hi_lo_lo_hi_hi_14, regroupV0_hi_lo_lo_hi_lo_14};
  wire [255:0]       regroupV0_hi_lo_lo_14 = {regroupV0_hi_lo_lo_hi_14, regroupV0_hi_lo_lo_lo_14};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo_lo_3 = {regroupV0_hi_12[1031], regroupV0_hi_12[1027]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo_hi_3 = {regroupV0_hi_12[1039], regroupV0_hi_12[1035]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo_7 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo_hi_3, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi_lo_3 = {regroupV0_hi_12[1047], regroupV0_hi_12[1043]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi_hi_3 = {regroupV0_hi_12[1055], regroupV0_hi_12[1051]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi_7 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi_hi_3, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_11 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_hi_7, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo_lo_3 = {regroupV0_hi_12[1063], regroupV0_hi_12[1059]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo_hi_3 = {regroupV0_hi_12[1071], regroupV0_hi_12[1067]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo_7 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo_hi_3, regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi_lo_3 = {regroupV0_hi_12[1079], regroupV0_hi_12[1075]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi_hi_3 = {regroupV0_hi_12[1087], regroupV0_hi_12[1083]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi_7 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi_hi_3, regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_11 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_hi_7, regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_lo_lo_14 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_11, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo_lo_3 = {regroupV0_hi_12[1095], regroupV0_hi_12[1091]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo_hi_3 = {regroupV0_hi_12[1103], regroupV0_hi_12[1099]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo_7 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo_hi_3, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi_lo_3 = {regroupV0_hi_12[1111], regroupV0_hi_12[1107]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi_hi_3 = {regroupV0_hi_12[1119], regroupV0_hi_12[1115]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi_7 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi_hi_3, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_11 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_hi_7, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo_lo_3 = {regroupV0_hi_12[1127], regroupV0_hi_12[1123]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo_hi_3 = {regroupV0_hi_12[1135], regroupV0_hi_12[1131]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo_7 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo_hi_3, regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi_lo_3 = {regroupV0_hi_12[1143], regroupV0_hi_12[1139]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi_hi_3 = {regroupV0_hi_12[1151], regroupV0_hi_12[1147]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi_7 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi_hi_3, regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_11 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_hi_7, regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_lo_hi_14 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_11, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_11};
  wire [31:0]        regroupV0_hi_lo_hi_lo_lo_lo_14 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_14, regroupV0_hi_lo_hi_lo_lo_lo_lo_14};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo_lo_3 = {regroupV0_hi_12[1159], regroupV0_hi_12[1155]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo_hi_3 = {regroupV0_hi_12[1167], regroupV0_hi_12[1163]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo_7 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo_hi_3, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi_lo_3 = {regroupV0_hi_12[1175], regroupV0_hi_12[1171]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi_hi_3 = {regroupV0_hi_12[1183], regroupV0_hi_12[1179]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi_7 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi_hi_3, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_11 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_hi_7, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo_lo_3 = {regroupV0_hi_12[1191], regroupV0_hi_12[1187]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo_hi_3 = {regroupV0_hi_12[1199], regroupV0_hi_12[1195]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo_7 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo_hi_3, regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi_lo_3 = {regroupV0_hi_12[1207], regroupV0_hi_12[1203]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi_hi_3 = {regroupV0_hi_12[1215], regroupV0_hi_12[1211]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi_7 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi_hi_3, regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_11 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_hi_7, regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_hi_lo_14 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_11, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo_lo_3 = {regroupV0_hi_12[1223], regroupV0_hi_12[1219]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo_hi_3 = {regroupV0_hi_12[1231], regroupV0_hi_12[1227]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo_7 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo_hi_3, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi_lo_3 = {regroupV0_hi_12[1239], regroupV0_hi_12[1235]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi_hi_3 = {regroupV0_hi_12[1247], regroupV0_hi_12[1243]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi_7 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi_hi_3, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_11 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_hi_7, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo_lo_3 = {regroupV0_hi_12[1255], regroupV0_hi_12[1251]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo_hi_3 = {regroupV0_hi_12[1263], regroupV0_hi_12[1259]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo_7 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo_hi_3, regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi_lo_3 = {regroupV0_hi_12[1271], regroupV0_hi_12[1267]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi_hi_3 = {regroupV0_hi_12[1279], regroupV0_hi_12[1275]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi_7 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi_hi_3, regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_11 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_hi_7, regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_hi_hi_14 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_11, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_11};
  wire [31:0]        regroupV0_hi_lo_hi_lo_lo_hi_14 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_14, regroupV0_hi_lo_hi_lo_lo_hi_lo_14};
  wire [63:0]        regroupV0_hi_lo_hi_lo_lo_14 = {regroupV0_hi_lo_hi_lo_lo_hi_14, regroupV0_hi_lo_hi_lo_lo_lo_14};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo_lo_3 = {regroupV0_hi_12[1287], regroupV0_hi_12[1283]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo_hi_3 = {regroupV0_hi_12[1295], regroupV0_hi_12[1291]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo_7 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo_hi_3, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi_lo_3 = {regroupV0_hi_12[1303], regroupV0_hi_12[1299]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi_hi_3 = {regroupV0_hi_12[1311], regroupV0_hi_12[1307]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi_7 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi_hi_3, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_11 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_hi_7, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo_lo_3 = {regroupV0_hi_12[1319], regroupV0_hi_12[1315]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo_hi_3 = {regroupV0_hi_12[1327], regroupV0_hi_12[1323]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo_7 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo_hi_3, regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi_lo_3 = {regroupV0_hi_12[1335], regroupV0_hi_12[1331]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi_hi_3 = {regroupV0_hi_12[1343], regroupV0_hi_12[1339]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi_7 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi_hi_3, regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_11 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_hi_7, regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_lo_lo_14 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_11, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo_lo_3 = {regroupV0_hi_12[1351], regroupV0_hi_12[1347]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo_hi_3 = {regroupV0_hi_12[1359], regroupV0_hi_12[1355]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo_7 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo_hi_3, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi_lo_3 = {regroupV0_hi_12[1367], regroupV0_hi_12[1363]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi_hi_3 = {regroupV0_hi_12[1375], regroupV0_hi_12[1371]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi_7 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi_hi_3, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_11 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_hi_7, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo_lo_3 = {regroupV0_hi_12[1383], regroupV0_hi_12[1379]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo_hi_3 = {regroupV0_hi_12[1391], regroupV0_hi_12[1387]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo_7 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo_hi_3, regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi_lo_3 = {regroupV0_hi_12[1399], regroupV0_hi_12[1395]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi_hi_3 = {regroupV0_hi_12[1407], regroupV0_hi_12[1403]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi_7 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi_hi_3, regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_11 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_hi_7, regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_lo_hi_14 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_11, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_11};
  wire [31:0]        regroupV0_hi_lo_hi_lo_hi_lo_14 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_14, regroupV0_hi_lo_hi_lo_hi_lo_lo_14};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo_lo_3 = {regroupV0_hi_12[1415], regroupV0_hi_12[1411]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo_hi_3 = {regroupV0_hi_12[1423], regroupV0_hi_12[1419]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo_7 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo_hi_3, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi_lo_3 = {regroupV0_hi_12[1431], regroupV0_hi_12[1427]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi_hi_3 = {regroupV0_hi_12[1439], regroupV0_hi_12[1435]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi_7 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi_hi_3, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_11 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_hi_7, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo_lo_3 = {regroupV0_hi_12[1447], regroupV0_hi_12[1443]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo_hi_3 = {regroupV0_hi_12[1455], regroupV0_hi_12[1451]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo_7 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo_hi_3, regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi_lo_3 = {regroupV0_hi_12[1463], regroupV0_hi_12[1459]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi_hi_3 = {regroupV0_hi_12[1471], regroupV0_hi_12[1467]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi_7 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi_hi_3, regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_11 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_hi_7, regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_hi_lo_14 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_11, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo_lo_3 = {regroupV0_hi_12[1479], regroupV0_hi_12[1475]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo_hi_3 = {regroupV0_hi_12[1487], regroupV0_hi_12[1483]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo_7 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo_hi_3, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi_lo_3 = {regroupV0_hi_12[1495], regroupV0_hi_12[1491]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi_hi_3 = {regroupV0_hi_12[1503], regroupV0_hi_12[1499]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi_7 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi_hi_3, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_11 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_hi_7, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo_lo_3 = {regroupV0_hi_12[1511], regroupV0_hi_12[1507]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo_hi_3 = {regroupV0_hi_12[1519], regroupV0_hi_12[1515]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo_7 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo_hi_3, regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi_lo_3 = {regroupV0_hi_12[1527], regroupV0_hi_12[1523]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi_hi_3 = {regroupV0_hi_12[1535], regroupV0_hi_12[1531]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi_7 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi_hi_3, regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_11 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_hi_7, regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_hi_hi_14 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_11, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_11};
  wire [31:0]        regroupV0_hi_lo_hi_lo_hi_hi_14 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_14, regroupV0_hi_lo_hi_lo_hi_hi_lo_14};
  wire [63:0]        regroupV0_hi_lo_hi_lo_hi_14 = {regroupV0_hi_lo_hi_lo_hi_hi_14, regroupV0_hi_lo_hi_lo_hi_lo_14};
  wire [127:0]       regroupV0_hi_lo_hi_lo_14 = {regroupV0_hi_lo_hi_lo_hi_14, regroupV0_hi_lo_hi_lo_lo_14};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo_lo_3 = {regroupV0_hi_12[1543], regroupV0_hi_12[1539]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo_hi_3 = {regroupV0_hi_12[1551], regroupV0_hi_12[1547]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo_7 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo_hi_3, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi_lo_3 = {regroupV0_hi_12[1559], regroupV0_hi_12[1555]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi_hi_3 = {regroupV0_hi_12[1567], regroupV0_hi_12[1563]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi_7 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi_hi_3, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_11 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_hi_7, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo_lo_3 = {regroupV0_hi_12[1575], regroupV0_hi_12[1571]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo_hi_3 = {regroupV0_hi_12[1583], regroupV0_hi_12[1579]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo_7 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo_hi_3, regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi_lo_3 = {regroupV0_hi_12[1591], regroupV0_hi_12[1587]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi_hi_3 = {regroupV0_hi_12[1599], regroupV0_hi_12[1595]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi_7 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi_hi_3, regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_11 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_hi_7, regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_lo_lo_14 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_11, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo_lo_3 = {regroupV0_hi_12[1607], regroupV0_hi_12[1603]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo_hi_3 = {regroupV0_hi_12[1615], regroupV0_hi_12[1611]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo_7 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo_hi_3, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi_lo_3 = {regroupV0_hi_12[1623], regroupV0_hi_12[1619]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi_hi_3 = {regroupV0_hi_12[1631], regroupV0_hi_12[1627]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi_7 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi_hi_3, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_11 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_hi_7, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo_lo_3 = {regroupV0_hi_12[1639], regroupV0_hi_12[1635]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo_hi_3 = {regroupV0_hi_12[1647], regroupV0_hi_12[1643]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo_7 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo_hi_3, regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi_lo_3 = {regroupV0_hi_12[1655], regroupV0_hi_12[1651]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi_hi_3 = {regroupV0_hi_12[1663], regroupV0_hi_12[1659]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi_7 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi_hi_3, regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_11 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_hi_7, regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_lo_hi_14 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_11, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_11};
  wire [31:0]        regroupV0_hi_lo_hi_hi_lo_lo_14 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_14, regroupV0_hi_lo_hi_hi_lo_lo_lo_14};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo_lo_3 = {regroupV0_hi_12[1671], regroupV0_hi_12[1667]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo_hi_3 = {regroupV0_hi_12[1679], regroupV0_hi_12[1675]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo_7 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo_hi_3, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi_lo_3 = {regroupV0_hi_12[1687], regroupV0_hi_12[1683]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi_hi_3 = {regroupV0_hi_12[1695], regroupV0_hi_12[1691]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi_7 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi_hi_3, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_11 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_hi_7, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo_lo_3 = {regroupV0_hi_12[1703], regroupV0_hi_12[1699]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo_hi_3 = {regroupV0_hi_12[1711], regroupV0_hi_12[1707]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo_7 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo_hi_3, regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi_lo_3 = {regroupV0_hi_12[1719], regroupV0_hi_12[1715]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi_hi_3 = {regroupV0_hi_12[1727], regroupV0_hi_12[1723]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi_7 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi_hi_3, regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_11 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_hi_7, regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_hi_lo_14 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_11, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo_lo_3 = {regroupV0_hi_12[1735], regroupV0_hi_12[1731]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo_hi_3 = {regroupV0_hi_12[1743], regroupV0_hi_12[1739]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo_7 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo_hi_3, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi_lo_3 = {regroupV0_hi_12[1751], regroupV0_hi_12[1747]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi_hi_3 = {regroupV0_hi_12[1759], regroupV0_hi_12[1755]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi_7 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi_hi_3, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_11 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_hi_7, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo_lo_3 = {regroupV0_hi_12[1767], regroupV0_hi_12[1763]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo_hi_3 = {regroupV0_hi_12[1775], regroupV0_hi_12[1771]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo_7 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo_hi_3, regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi_lo_3 = {regroupV0_hi_12[1783], regroupV0_hi_12[1779]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi_hi_3 = {regroupV0_hi_12[1791], regroupV0_hi_12[1787]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi_7 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi_hi_3, regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_11 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_hi_7, regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_hi_hi_14 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_11, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_11};
  wire [31:0]        regroupV0_hi_lo_hi_hi_lo_hi_14 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_14, regroupV0_hi_lo_hi_hi_lo_hi_lo_14};
  wire [63:0]        regroupV0_hi_lo_hi_hi_lo_14 = {regroupV0_hi_lo_hi_hi_lo_hi_14, regroupV0_hi_lo_hi_hi_lo_lo_14};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo_lo_3 = {regroupV0_hi_12[1799], regroupV0_hi_12[1795]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo_hi_3 = {regroupV0_hi_12[1807], regroupV0_hi_12[1803]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo_7 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo_hi_3, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi_lo_3 = {regroupV0_hi_12[1815], regroupV0_hi_12[1811]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi_hi_3 = {regroupV0_hi_12[1823], regroupV0_hi_12[1819]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi_7 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi_hi_3, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_11 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_hi_7, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo_lo_3 = {regroupV0_hi_12[1831], regroupV0_hi_12[1827]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo_hi_3 = {regroupV0_hi_12[1839], regroupV0_hi_12[1835]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo_7 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo_hi_3, regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi_lo_3 = {regroupV0_hi_12[1847], regroupV0_hi_12[1843]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi_hi_3 = {regroupV0_hi_12[1855], regroupV0_hi_12[1851]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi_7 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi_hi_3, regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_11 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_hi_7, regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_lo_lo_14 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_11, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo_lo_3 = {regroupV0_hi_12[1863], regroupV0_hi_12[1859]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo_hi_3 = {regroupV0_hi_12[1871], regroupV0_hi_12[1867]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo_7 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo_hi_3, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi_lo_3 = {regroupV0_hi_12[1879], regroupV0_hi_12[1875]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi_hi_3 = {regroupV0_hi_12[1887], regroupV0_hi_12[1883]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi_7 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi_hi_3, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_11 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_hi_7, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo_lo_3 = {regroupV0_hi_12[1895], regroupV0_hi_12[1891]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo_hi_3 = {regroupV0_hi_12[1903], regroupV0_hi_12[1899]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo_7 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo_hi_3, regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi_lo_3 = {regroupV0_hi_12[1911], regroupV0_hi_12[1907]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi_hi_3 = {regroupV0_hi_12[1919], regroupV0_hi_12[1915]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi_7 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi_hi_3, regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_11 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_hi_7, regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_lo_hi_14 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_11, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_11};
  wire [31:0]        regroupV0_hi_lo_hi_hi_hi_lo_14 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_14, regroupV0_hi_lo_hi_hi_hi_lo_lo_14};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo_lo_3 = {regroupV0_hi_12[1927], regroupV0_hi_12[1923]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo_hi_3 = {regroupV0_hi_12[1935], regroupV0_hi_12[1931]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo_7 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo_hi_3, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi_lo_3 = {regroupV0_hi_12[1943], regroupV0_hi_12[1939]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi_hi_3 = {regroupV0_hi_12[1951], regroupV0_hi_12[1947]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi_7 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi_hi_3, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_11 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_hi_7, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo_lo_3 = {regroupV0_hi_12[1959], regroupV0_hi_12[1955]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo_hi_3 = {regroupV0_hi_12[1967], regroupV0_hi_12[1963]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo_7 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo_hi_3, regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi_lo_3 = {regroupV0_hi_12[1975], regroupV0_hi_12[1971]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi_hi_3 = {regroupV0_hi_12[1983], regroupV0_hi_12[1979]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi_7 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi_hi_3, regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_11 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_hi_7, regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_hi_lo_14 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_11, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo_lo_3 = {regroupV0_hi_12[1991], regroupV0_hi_12[1987]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo_hi_3 = {regroupV0_hi_12[1999], regroupV0_hi_12[1995]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo_7 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo_hi_3, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi_lo_3 = {regroupV0_hi_12[2007], regroupV0_hi_12[2003]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi_hi_3 = {regroupV0_hi_12[2015], regroupV0_hi_12[2011]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi_7 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi_hi_3, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_11 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_hi_7, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo_lo_3 = {regroupV0_hi_12[2023], regroupV0_hi_12[2019]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo_hi_3 = {regroupV0_hi_12[2031], regroupV0_hi_12[2027]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo_7 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo_hi_3, regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi_lo_3 = {regroupV0_hi_12[2039], regroupV0_hi_12[2035]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi_hi_3 = {regroupV0_hi_12[2047], regroupV0_hi_12[2043]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi_7 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi_hi_3, regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_11 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_hi_7, regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_hi_hi_14 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_11, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_11};
  wire [31:0]        regroupV0_hi_lo_hi_hi_hi_hi_14 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_14, regroupV0_hi_lo_hi_hi_hi_hi_lo_14};
  wire [63:0]        regroupV0_hi_lo_hi_hi_hi_14 = {regroupV0_hi_lo_hi_hi_hi_hi_14, regroupV0_hi_lo_hi_hi_hi_lo_14};
  wire [127:0]       regroupV0_hi_lo_hi_hi_14 = {regroupV0_hi_lo_hi_hi_hi_14, regroupV0_hi_lo_hi_hi_lo_14};
  wire [255:0]       regroupV0_hi_lo_hi_14 = {regroupV0_hi_lo_hi_hi_14, regroupV0_hi_lo_hi_lo_14};
  wire [511:0]       regroupV0_hi_lo_14 = {regroupV0_hi_lo_hi_14, regroupV0_hi_lo_lo_14};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo_lo_3 = {regroupV0_hi_12[2055], regroupV0_hi_12[2051]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo_hi_3 = {regroupV0_hi_12[2063], regroupV0_hi_12[2059]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo_7 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo_hi_3, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi_lo_3 = {regroupV0_hi_12[2071], regroupV0_hi_12[2067]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi_hi_3 = {regroupV0_hi_12[2079], regroupV0_hi_12[2075]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi_7 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi_hi_3, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_11 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_hi_7, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo_lo_3 = {regroupV0_hi_12[2087], regroupV0_hi_12[2083]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo_hi_3 = {regroupV0_hi_12[2095], regroupV0_hi_12[2091]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo_7 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo_hi_3, regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi_lo_3 = {regroupV0_hi_12[2103], regroupV0_hi_12[2099]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi_hi_3 = {regroupV0_hi_12[2111], regroupV0_hi_12[2107]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi_7 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi_hi_3, regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_11 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_hi_7, regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_lo_lo_14 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_11, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo_lo_3 = {regroupV0_hi_12[2119], regroupV0_hi_12[2115]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo_hi_3 = {regroupV0_hi_12[2127], regroupV0_hi_12[2123]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo_7 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo_hi_3, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi_lo_3 = {regroupV0_hi_12[2135], regroupV0_hi_12[2131]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi_hi_3 = {regroupV0_hi_12[2143], regroupV0_hi_12[2139]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi_7 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi_hi_3, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_11 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_hi_7, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo_lo_3 = {regroupV0_hi_12[2151], regroupV0_hi_12[2147]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo_hi_3 = {regroupV0_hi_12[2159], regroupV0_hi_12[2155]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo_7 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo_hi_3, regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi_lo_3 = {regroupV0_hi_12[2167], regroupV0_hi_12[2163]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi_hi_3 = {regroupV0_hi_12[2175], regroupV0_hi_12[2171]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi_7 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi_hi_3, regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_11 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_hi_7, regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_lo_hi_14 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_11, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_11};
  wire [31:0]        regroupV0_hi_hi_lo_lo_lo_lo_14 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_14, regroupV0_hi_hi_lo_lo_lo_lo_lo_14};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo_lo_3 = {regroupV0_hi_12[2183], regroupV0_hi_12[2179]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo_hi_3 = {regroupV0_hi_12[2191], regroupV0_hi_12[2187]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo_7 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo_hi_3, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi_lo_3 = {regroupV0_hi_12[2199], regroupV0_hi_12[2195]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi_hi_3 = {regroupV0_hi_12[2207], regroupV0_hi_12[2203]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi_7 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi_hi_3, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_11 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_hi_7, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo_lo_3 = {regroupV0_hi_12[2215], regroupV0_hi_12[2211]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo_hi_3 = {regroupV0_hi_12[2223], regroupV0_hi_12[2219]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo_7 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo_hi_3, regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi_lo_3 = {regroupV0_hi_12[2231], regroupV0_hi_12[2227]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi_hi_3 = {regroupV0_hi_12[2239], regroupV0_hi_12[2235]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi_7 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi_hi_3, regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_11 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_hi_7, regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_hi_lo_14 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_11, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo_lo_3 = {regroupV0_hi_12[2247], regroupV0_hi_12[2243]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo_hi_3 = {regroupV0_hi_12[2255], regroupV0_hi_12[2251]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo_7 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo_hi_3, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi_lo_3 = {regroupV0_hi_12[2263], regroupV0_hi_12[2259]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi_hi_3 = {regroupV0_hi_12[2271], regroupV0_hi_12[2267]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi_7 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi_hi_3, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_11 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_hi_7, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo_lo_3 = {regroupV0_hi_12[2279], regroupV0_hi_12[2275]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo_hi_3 = {regroupV0_hi_12[2287], regroupV0_hi_12[2283]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo_7 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo_hi_3, regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi_lo_3 = {regroupV0_hi_12[2295], regroupV0_hi_12[2291]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi_hi_3 = {regroupV0_hi_12[2303], regroupV0_hi_12[2299]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi_7 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi_hi_3, regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_11 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_hi_7, regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_hi_hi_14 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_11, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_11};
  wire [31:0]        regroupV0_hi_hi_lo_lo_lo_hi_14 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_14, regroupV0_hi_hi_lo_lo_lo_hi_lo_14};
  wire [63:0]        regroupV0_hi_hi_lo_lo_lo_14 = {regroupV0_hi_hi_lo_lo_lo_hi_14, regroupV0_hi_hi_lo_lo_lo_lo_14};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo_lo_3 = {regroupV0_hi_12[2311], regroupV0_hi_12[2307]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo_hi_3 = {regroupV0_hi_12[2319], regroupV0_hi_12[2315]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo_7 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo_hi_3, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi_lo_3 = {regroupV0_hi_12[2327], regroupV0_hi_12[2323]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi_hi_3 = {regroupV0_hi_12[2335], regroupV0_hi_12[2331]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi_7 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi_hi_3, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_11 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_hi_7, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo_lo_3 = {regroupV0_hi_12[2343], regroupV0_hi_12[2339]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo_hi_3 = {regroupV0_hi_12[2351], regroupV0_hi_12[2347]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo_7 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo_hi_3, regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi_lo_3 = {regroupV0_hi_12[2359], regroupV0_hi_12[2355]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi_hi_3 = {regroupV0_hi_12[2367], regroupV0_hi_12[2363]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi_7 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi_hi_3, regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_11 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_hi_7, regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_lo_lo_14 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_11, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo_lo_3 = {regroupV0_hi_12[2375], regroupV0_hi_12[2371]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo_hi_3 = {regroupV0_hi_12[2383], regroupV0_hi_12[2379]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo_7 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo_hi_3, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi_lo_3 = {regroupV0_hi_12[2391], regroupV0_hi_12[2387]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi_hi_3 = {regroupV0_hi_12[2399], regroupV0_hi_12[2395]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi_7 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi_hi_3, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_11 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_hi_7, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo_lo_3 = {regroupV0_hi_12[2407], regroupV0_hi_12[2403]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo_hi_3 = {regroupV0_hi_12[2415], regroupV0_hi_12[2411]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo_7 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo_hi_3, regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi_lo_3 = {regroupV0_hi_12[2423], regroupV0_hi_12[2419]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi_hi_3 = {regroupV0_hi_12[2431], regroupV0_hi_12[2427]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi_7 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi_hi_3, regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_11 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_hi_7, regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_lo_hi_14 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_11, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_11};
  wire [31:0]        regroupV0_hi_hi_lo_lo_hi_lo_14 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_14, regroupV0_hi_hi_lo_lo_hi_lo_lo_14};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo_lo_3 = {regroupV0_hi_12[2439], regroupV0_hi_12[2435]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo_hi_3 = {regroupV0_hi_12[2447], regroupV0_hi_12[2443]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo_7 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo_hi_3, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi_lo_3 = {regroupV0_hi_12[2455], regroupV0_hi_12[2451]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi_hi_3 = {regroupV0_hi_12[2463], regroupV0_hi_12[2459]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi_7 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi_hi_3, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_11 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_hi_7, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo_lo_3 = {regroupV0_hi_12[2471], regroupV0_hi_12[2467]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo_hi_3 = {regroupV0_hi_12[2479], regroupV0_hi_12[2475]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo_7 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo_hi_3, regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi_lo_3 = {regroupV0_hi_12[2487], regroupV0_hi_12[2483]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi_hi_3 = {regroupV0_hi_12[2495], regroupV0_hi_12[2491]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi_7 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi_hi_3, regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_11 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_hi_7, regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_hi_lo_14 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_11, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo_lo_3 = {regroupV0_hi_12[2503], regroupV0_hi_12[2499]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo_hi_3 = {regroupV0_hi_12[2511], regroupV0_hi_12[2507]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo_7 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo_hi_3, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi_lo_3 = {regroupV0_hi_12[2519], regroupV0_hi_12[2515]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi_hi_3 = {regroupV0_hi_12[2527], regroupV0_hi_12[2523]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi_7 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi_hi_3, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_11 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_hi_7, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo_lo_3 = {regroupV0_hi_12[2535], regroupV0_hi_12[2531]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo_hi_3 = {regroupV0_hi_12[2543], regroupV0_hi_12[2539]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo_7 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo_hi_3, regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi_lo_3 = {regroupV0_hi_12[2551], regroupV0_hi_12[2547]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi_hi_3 = {regroupV0_hi_12[2559], regroupV0_hi_12[2555]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi_7 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi_hi_3, regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_11 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_hi_7, regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_hi_hi_14 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_11, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_11};
  wire [31:0]        regroupV0_hi_hi_lo_lo_hi_hi_14 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_14, regroupV0_hi_hi_lo_lo_hi_hi_lo_14};
  wire [63:0]        regroupV0_hi_hi_lo_lo_hi_14 = {regroupV0_hi_hi_lo_lo_hi_hi_14, regroupV0_hi_hi_lo_lo_hi_lo_14};
  wire [127:0]       regroupV0_hi_hi_lo_lo_14 = {regroupV0_hi_hi_lo_lo_hi_14, regroupV0_hi_hi_lo_lo_lo_14};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo_lo_3 = {regroupV0_hi_12[2567], regroupV0_hi_12[2563]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo_hi_3 = {regroupV0_hi_12[2575], regroupV0_hi_12[2571]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo_7 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo_hi_3, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi_lo_3 = {regroupV0_hi_12[2583], regroupV0_hi_12[2579]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi_hi_3 = {regroupV0_hi_12[2591], regroupV0_hi_12[2587]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi_7 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi_hi_3, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_11 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_hi_7, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo_lo_3 = {regroupV0_hi_12[2599], regroupV0_hi_12[2595]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo_hi_3 = {regroupV0_hi_12[2607], regroupV0_hi_12[2603]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo_7 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo_hi_3, regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi_lo_3 = {regroupV0_hi_12[2615], regroupV0_hi_12[2611]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi_hi_3 = {regroupV0_hi_12[2623], regroupV0_hi_12[2619]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi_7 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi_hi_3, regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_11 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_hi_7, regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_lo_lo_14 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_11, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo_lo_3 = {regroupV0_hi_12[2631], regroupV0_hi_12[2627]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo_hi_3 = {regroupV0_hi_12[2639], regroupV0_hi_12[2635]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo_7 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo_hi_3, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi_lo_3 = {regroupV0_hi_12[2647], regroupV0_hi_12[2643]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi_hi_3 = {regroupV0_hi_12[2655], regroupV0_hi_12[2651]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi_7 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi_hi_3, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_11 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_hi_7, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo_lo_3 = {regroupV0_hi_12[2663], regroupV0_hi_12[2659]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo_hi_3 = {regroupV0_hi_12[2671], regroupV0_hi_12[2667]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo_7 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo_hi_3, regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi_lo_3 = {regroupV0_hi_12[2679], regroupV0_hi_12[2675]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi_hi_3 = {regroupV0_hi_12[2687], regroupV0_hi_12[2683]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi_7 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi_hi_3, regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_11 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_hi_7, regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_lo_hi_14 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_11, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_11};
  wire [31:0]        regroupV0_hi_hi_lo_hi_lo_lo_14 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_14, regroupV0_hi_hi_lo_hi_lo_lo_lo_14};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo_lo_3 = {regroupV0_hi_12[2695], regroupV0_hi_12[2691]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo_hi_3 = {regroupV0_hi_12[2703], regroupV0_hi_12[2699]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo_7 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo_hi_3, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi_lo_3 = {regroupV0_hi_12[2711], regroupV0_hi_12[2707]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi_hi_3 = {regroupV0_hi_12[2719], regroupV0_hi_12[2715]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi_7 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi_hi_3, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_11 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_hi_7, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo_lo_3 = {regroupV0_hi_12[2727], regroupV0_hi_12[2723]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo_hi_3 = {regroupV0_hi_12[2735], regroupV0_hi_12[2731]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo_7 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo_hi_3, regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi_lo_3 = {regroupV0_hi_12[2743], regroupV0_hi_12[2739]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi_hi_3 = {regroupV0_hi_12[2751], regroupV0_hi_12[2747]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi_7 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi_hi_3, regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_11 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_hi_7, regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_hi_lo_14 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_11, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo_lo_3 = {regroupV0_hi_12[2759], regroupV0_hi_12[2755]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo_hi_3 = {regroupV0_hi_12[2767], regroupV0_hi_12[2763]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo_7 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo_hi_3, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi_lo_3 = {regroupV0_hi_12[2775], regroupV0_hi_12[2771]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi_hi_3 = {regroupV0_hi_12[2783], regroupV0_hi_12[2779]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi_7 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi_hi_3, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_11 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_hi_7, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo_lo_3 = {regroupV0_hi_12[2791], regroupV0_hi_12[2787]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo_hi_3 = {regroupV0_hi_12[2799], regroupV0_hi_12[2795]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo_7 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo_hi_3, regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi_lo_3 = {regroupV0_hi_12[2807], regroupV0_hi_12[2803]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi_hi_3 = {regroupV0_hi_12[2815], regroupV0_hi_12[2811]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi_7 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi_hi_3, regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_11 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_hi_7, regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_hi_hi_14 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_11, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_11};
  wire [31:0]        regroupV0_hi_hi_lo_hi_lo_hi_14 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_14, regroupV0_hi_hi_lo_hi_lo_hi_lo_14};
  wire [63:0]        regroupV0_hi_hi_lo_hi_lo_14 = {regroupV0_hi_hi_lo_hi_lo_hi_14, regroupV0_hi_hi_lo_hi_lo_lo_14};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo_lo_3 = {regroupV0_hi_12[2823], regroupV0_hi_12[2819]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo_hi_3 = {regroupV0_hi_12[2831], regroupV0_hi_12[2827]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo_7 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo_hi_3, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi_lo_3 = {regroupV0_hi_12[2839], regroupV0_hi_12[2835]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi_hi_3 = {regroupV0_hi_12[2847], regroupV0_hi_12[2843]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi_7 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi_hi_3, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_11 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_hi_7, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo_lo_3 = {regroupV0_hi_12[2855], regroupV0_hi_12[2851]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo_hi_3 = {regroupV0_hi_12[2863], regroupV0_hi_12[2859]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo_7 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo_hi_3, regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi_lo_3 = {regroupV0_hi_12[2871], regroupV0_hi_12[2867]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi_hi_3 = {regroupV0_hi_12[2879], regroupV0_hi_12[2875]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi_7 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi_hi_3, regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_11 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_hi_7, regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_lo_lo_14 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_11, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo_lo_3 = {regroupV0_hi_12[2887], regroupV0_hi_12[2883]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo_hi_3 = {regroupV0_hi_12[2895], regroupV0_hi_12[2891]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo_7 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo_hi_3, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi_lo_3 = {regroupV0_hi_12[2903], regroupV0_hi_12[2899]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi_hi_3 = {regroupV0_hi_12[2911], regroupV0_hi_12[2907]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi_7 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi_hi_3, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_11 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_hi_7, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo_lo_3 = {regroupV0_hi_12[2919], regroupV0_hi_12[2915]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo_hi_3 = {regroupV0_hi_12[2927], regroupV0_hi_12[2923]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo_7 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo_hi_3, regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi_lo_3 = {regroupV0_hi_12[2935], regroupV0_hi_12[2931]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi_hi_3 = {regroupV0_hi_12[2943], regroupV0_hi_12[2939]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi_7 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi_hi_3, regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_11 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_hi_7, regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_lo_hi_14 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_11, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_11};
  wire [31:0]        regroupV0_hi_hi_lo_hi_hi_lo_14 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_14, regroupV0_hi_hi_lo_hi_hi_lo_lo_14};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo_lo_3 = {regroupV0_hi_12[2951], regroupV0_hi_12[2947]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo_hi_3 = {regroupV0_hi_12[2959], regroupV0_hi_12[2955]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo_7 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo_hi_3, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi_lo_3 = {regroupV0_hi_12[2967], regroupV0_hi_12[2963]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi_hi_3 = {regroupV0_hi_12[2975], regroupV0_hi_12[2971]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi_7 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi_hi_3, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_11 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_hi_7, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo_lo_3 = {regroupV0_hi_12[2983], regroupV0_hi_12[2979]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo_hi_3 = {regroupV0_hi_12[2991], regroupV0_hi_12[2987]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo_7 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo_hi_3, regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi_lo_3 = {regroupV0_hi_12[2999], regroupV0_hi_12[2995]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi_hi_3 = {regroupV0_hi_12[3007], regroupV0_hi_12[3003]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi_7 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi_hi_3, regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_11 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_hi_7, regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_hi_lo_14 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_11, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo_lo_3 = {regroupV0_hi_12[3015], regroupV0_hi_12[3011]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo_hi_3 = {regroupV0_hi_12[3023], regroupV0_hi_12[3019]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo_7 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo_hi_3, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi_lo_3 = {regroupV0_hi_12[3031], regroupV0_hi_12[3027]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi_hi_3 = {regroupV0_hi_12[3039], regroupV0_hi_12[3035]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi_7 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi_hi_3, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_11 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_hi_7, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo_lo_3 = {regroupV0_hi_12[3047], regroupV0_hi_12[3043]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo_hi_3 = {regroupV0_hi_12[3055], regroupV0_hi_12[3051]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo_7 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo_hi_3, regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi_lo_3 = {regroupV0_hi_12[3063], regroupV0_hi_12[3059]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi_hi_3 = {regroupV0_hi_12[3071], regroupV0_hi_12[3067]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi_7 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi_hi_3, regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_11 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_hi_7, regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_hi_hi_14 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_11, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_11};
  wire [31:0]        regroupV0_hi_hi_lo_hi_hi_hi_14 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_14, regroupV0_hi_hi_lo_hi_hi_hi_lo_14};
  wire [63:0]        regroupV0_hi_hi_lo_hi_hi_14 = {regroupV0_hi_hi_lo_hi_hi_hi_14, regroupV0_hi_hi_lo_hi_hi_lo_14};
  wire [127:0]       regroupV0_hi_hi_lo_hi_14 = {regroupV0_hi_hi_lo_hi_hi_14, regroupV0_hi_hi_lo_hi_lo_14};
  wire [255:0]       regroupV0_hi_hi_lo_14 = {regroupV0_hi_hi_lo_hi_14, regroupV0_hi_hi_lo_lo_14};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo_lo_3 = {regroupV0_hi_12[3079], regroupV0_hi_12[3075]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo_hi_3 = {regroupV0_hi_12[3087], regroupV0_hi_12[3083]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo_7 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo_hi_3, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi_lo_3 = {regroupV0_hi_12[3095], regroupV0_hi_12[3091]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi_hi_3 = {regroupV0_hi_12[3103], regroupV0_hi_12[3099]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi_7 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi_hi_3, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_11 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_hi_7, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo_lo_3 = {regroupV0_hi_12[3111], regroupV0_hi_12[3107]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo_hi_3 = {regroupV0_hi_12[3119], regroupV0_hi_12[3115]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo_7 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo_hi_3, regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi_lo_3 = {regroupV0_hi_12[3127], regroupV0_hi_12[3123]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi_hi_3 = {regroupV0_hi_12[3135], regroupV0_hi_12[3131]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi_7 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi_hi_3, regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_11 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_hi_7, regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_lo_lo_14 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_11, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo_lo_3 = {regroupV0_hi_12[3143], regroupV0_hi_12[3139]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo_hi_3 = {regroupV0_hi_12[3151], regroupV0_hi_12[3147]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo_7 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo_hi_3, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi_lo_3 = {regroupV0_hi_12[3159], regroupV0_hi_12[3155]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi_hi_3 = {regroupV0_hi_12[3167], regroupV0_hi_12[3163]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi_7 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi_hi_3, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_11 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_hi_7, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo_lo_3 = {regroupV0_hi_12[3175], regroupV0_hi_12[3171]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo_hi_3 = {regroupV0_hi_12[3183], regroupV0_hi_12[3179]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo_7 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo_hi_3, regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi_lo_3 = {regroupV0_hi_12[3191], regroupV0_hi_12[3187]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi_hi_3 = {regroupV0_hi_12[3199], regroupV0_hi_12[3195]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi_7 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_11 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_hi_7, regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_lo_hi_14 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_11, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_11};
  wire [31:0]        regroupV0_hi_hi_hi_lo_lo_lo_14 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_14, regroupV0_hi_hi_hi_lo_lo_lo_lo_14};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo_lo_3 = {regroupV0_hi_12[3207], regroupV0_hi_12[3203]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo_hi_3 = {regroupV0_hi_12[3215], regroupV0_hi_12[3211]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo_7 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo_hi_3, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi_lo_3 = {regroupV0_hi_12[3223], regroupV0_hi_12[3219]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi_hi_3 = {regroupV0_hi_12[3231], regroupV0_hi_12[3227]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi_7 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi_hi_3, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_11 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_hi_7, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo_lo_3 = {regroupV0_hi_12[3239], regroupV0_hi_12[3235]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo_hi_3 = {regroupV0_hi_12[3247], regroupV0_hi_12[3243]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo_7 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo_hi_3, regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi_lo_3 = {regroupV0_hi_12[3255], regroupV0_hi_12[3251]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi_hi_3 = {regroupV0_hi_12[3263], regroupV0_hi_12[3259]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi_7 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi_hi_3, regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_11 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_hi_7, regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_hi_lo_14 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_11, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo_lo_3 = {regroupV0_hi_12[3271], regroupV0_hi_12[3267]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo_hi_3 = {regroupV0_hi_12[3279], regroupV0_hi_12[3275]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo_7 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo_hi_3, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi_lo_3 = {regroupV0_hi_12[3287], regroupV0_hi_12[3283]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi_hi_3 = {regroupV0_hi_12[3295], regroupV0_hi_12[3291]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi_7 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi_hi_3, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_11 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_hi_7, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo_lo_3 = {regroupV0_hi_12[3303], regroupV0_hi_12[3299]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo_hi_3 = {regroupV0_hi_12[3311], regroupV0_hi_12[3307]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo_7 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo_hi_3, regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi_lo_3 = {regroupV0_hi_12[3319], regroupV0_hi_12[3315]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi_hi_3 = {regroupV0_hi_12[3327], regroupV0_hi_12[3323]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi_7 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_11 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_hi_7, regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_hi_hi_14 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_11, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_11};
  wire [31:0]        regroupV0_hi_hi_hi_lo_lo_hi_14 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_14, regroupV0_hi_hi_hi_lo_lo_hi_lo_14};
  wire [63:0]        regroupV0_hi_hi_hi_lo_lo_14 = {regroupV0_hi_hi_hi_lo_lo_hi_14, regroupV0_hi_hi_hi_lo_lo_lo_14};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo_lo_3 = {regroupV0_hi_12[3335], regroupV0_hi_12[3331]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo_hi_3 = {regroupV0_hi_12[3343], regroupV0_hi_12[3339]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo_7 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo_hi_3, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi_lo_3 = {regroupV0_hi_12[3351], regroupV0_hi_12[3347]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi_hi_3 = {regroupV0_hi_12[3359], regroupV0_hi_12[3355]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi_7 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi_hi_3, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_11 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_hi_7, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo_lo_3 = {regroupV0_hi_12[3367], regroupV0_hi_12[3363]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo_hi_3 = {regroupV0_hi_12[3375], regroupV0_hi_12[3371]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo_7 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo_hi_3, regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi_lo_3 = {regroupV0_hi_12[3383], regroupV0_hi_12[3379]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi_hi_3 = {regroupV0_hi_12[3391], regroupV0_hi_12[3387]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi_7 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi_hi_3, regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_11 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_hi_7, regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_lo_lo_14 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_11, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo_lo_3 = {regroupV0_hi_12[3399], regroupV0_hi_12[3395]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo_hi_3 = {regroupV0_hi_12[3407], regroupV0_hi_12[3403]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo_7 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo_hi_3, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi_lo_3 = {regroupV0_hi_12[3415], regroupV0_hi_12[3411]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi_hi_3 = {regroupV0_hi_12[3423], regroupV0_hi_12[3419]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi_7 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi_hi_3, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_11 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_hi_7, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo_lo_3 = {regroupV0_hi_12[3431], regroupV0_hi_12[3427]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo_hi_3 = {regroupV0_hi_12[3439], regroupV0_hi_12[3435]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo_7 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo_hi_3, regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi_lo_3 = {regroupV0_hi_12[3447], regroupV0_hi_12[3443]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi_hi_3 = {regroupV0_hi_12[3455], regroupV0_hi_12[3451]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi_7 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_11 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_hi_7, regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_lo_hi_14 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_11, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_11};
  wire [31:0]        regroupV0_hi_hi_hi_lo_hi_lo_14 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_14, regroupV0_hi_hi_hi_lo_hi_lo_lo_14};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo_lo_3 = {regroupV0_hi_12[3463], regroupV0_hi_12[3459]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo_hi_3 = {regroupV0_hi_12[3471], regroupV0_hi_12[3467]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo_7 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo_hi_3, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi_lo_3 = {regroupV0_hi_12[3479], regroupV0_hi_12[3475]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi_hi_3 = {regroupV0_hi_12[3487], regroupV0_hi_12[3483]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi_7 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi_hi_3, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_11 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_hi_7, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo_lo_3 = {regroupV0_hi_12[3495], regroupV0_hi_12[3491]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo_hi_3 = {regroupV0_hi_12[3503], regroupV0_hi_12[3499]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo_7 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo_hi_3, regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi_lo_3 = {regroupV0_hi_12[3511], regroupV0_hi_12[3507]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi_hi_3 = {regroupV0_hi_12[3519], regroupV0_hi_12[3515]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi_7 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi_hi_3, regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_11 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_hi_7, regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_hi_lo_14 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_11, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo_lo_3 = {regroupV0_hi_12[3527], regroupV0_hi_12[3523]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo_hi_3 = {regroupV0_hi_12[3535], regroupV0_hi_12[3531]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo_7 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo_hi_3, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi_lo_3 = {regroupV0_hi_12[3543], regroupV0_hi_12[3539]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi_hi_3 = {regroupV0_hi_12[3551], regroupV0_hi_12[3547]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi_7 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi_hi_3, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_11 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_hi_7, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo_lo_3 = {regroupV0_hi_12[3559], regroupV0_hi_12[3555]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo_hi_3 = {regroupV0_hi_12[3567], regroupV0_hi_12[3563]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo_7 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo_hi_3, regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi_lo_3 = {regroupV0_hi_12[3575], regroupV0_hi_12[3571]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi_hi_3 = {regroupV0_hi_12[3583], regroupV0_hi_12[3579]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi_7 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_11 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_hi_7, regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_hi_hi_14 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_11, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_11};
  wire [31:0]        regroupV0_hi_hi_hi_lo_hi_hi_14 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_14, regroupV0_hi_hi_hi_lo_hi_hi_lo_14};
  wire [63:0]        regroupV0_hi_hi_hi_lo_hi_14 = {regroupV0_hi_hi_hi_lo_hi_hi_14, regroupV0_hi_hi_hi_lo_hi_lo_14};
  wire [127:0]       regroupV0_hi_hi_hi_lo_14 = {regroupV0_hi_hi_hi_lo_hi_14, regroupV0_hi_hi_hi_lo_lo_14};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo_lo_3 = {regroupV0_hi_12[3591], regroupV0_hi_12[3587]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo_hi_3 = {regroupV0_hi_12[3599], regroupV0_hi_12[3595]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo_7 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo_hi_3, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi_lo_3 = {regroupV0_hi_12[3607], regroupV0_hi_12[3603]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi_hi_3 = {regroupV0_hi_12[3615], regroupV0_hi_12[3611]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi_7 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi_hi_3, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_11 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_hi_7, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo_lo_3 = {regroupV0_hi_12[3623], regroupV0_hi_12[3619]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo_hi_3 = {regroupV0_hi_12[3631], regroupV0_hi_12[3627]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo_7 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo_hi_3, regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi_lo_3 = {regroupV0_hi_12[3639], regroupV0_hi_12[3635]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi_hi_3 = {regroupV0_hi_12[3647], regroupV0_hi_12[3643]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi_7 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi_hi_3, regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_11 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_hi_7, regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_lo_lo_14 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_11, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo_lo_3 = {regroupV0_hi_12[3655], regroupV0_hi_12[3651]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo_hi_3 = {regroupV0_hi_12[3663], regroupV0_hi_12[3659]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo_7 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo_hi_3, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi_lo_3 = {regroupV0_hi_12[3671], regroupV0_hi_12[3667]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi_hi_3 = {regroupV0_hi_12[3679], regroupV0_hi_12[3675]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi_7 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi_hi_3, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_11 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_hi_7, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo_lo_3 = {regroupV0_hi_12[3687], regroupV0_hi_12[3683]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo_hi_3 = {regroupV0_hi_12[3695], regroupV0_hi_12[3691]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo_7 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo_hi_3, regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi_lo_3 = {regroupV0_hi_12[3703], regroupV0_hi_12[3699]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi_hi_3 = {regroupV0_hi_12[3711], regroupV0_hi_12[3707]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi_7 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_11 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_hi_7, regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_lo_hi_14 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_11, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_11};
  wire [31:0]        regroupV0_hi_hi_hi_hi_lo_lo_14 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_14, regroupV0_hi_hi_hi_hi_lo_lo_lo_14};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo_lo_3 = {regroupV0_hi_12[3719], regroupV0_hi_12[3715]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo_hi_3 = {regroupV0_hi_12[3727], regroupV0_hi_12[3723]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo_7 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo_hi_3, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi_lo_3 = {regroupV0_hi_12[3735], regroupV0_hi_12[3731]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi_hi_3 = {regroupV0_hi_12[3743], regroupV0_hi_12[3739]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi_7 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi_hi_3, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_11 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_hi_7, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo_lo_3 = {regroupV0_hi_12[3751], regroupV0_hi_12[3747]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo_hi_3 = {regroupV0_hi_12[3759], regroupV0_hi_12[3755]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo_7 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo_hi_3, regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi_lo_3 = {regroupV0_hi_12[3767], regroupV0_hi_12[3763]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi_hi_3 = {regroupV0_hi_12[3775], regroupV0_hi_12[3771]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi_7 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi_hi_3, regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_11 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_hi_7, regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_hi_lo_14 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_11, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo_lo_3 = {regroupV0_hi_12[3783], regroupV0_hi_12[3779]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo_hi_3 = {regroupV0_hi_12[3791], regroupV0_hi_12[3787]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo_7 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo_hi_3, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi_lo_3 = {regroupV0_hi_12[3799], regroupV0_hi_12[3795]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi_hi_3 = {regroupV0_hi_12[3807], regroupV0_hi_12[3803]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi_7 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi_hi_3, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_11 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_hi_7, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo_lo_3 = {regroupV0_hi_12[3815], regroupV0_hi_12[3811]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo_hi_3 = {regroupV0_hi_12[3823], regroupV0_hi_12[3819]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo_7 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo_hi_3, regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi_lo_3 = {regroupV0_hi_12[3831], regroupV0_hi_12[3827]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi_hi_3 = {regroupV0_hi_12[3839], regroupV0_hi_12[3835]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi_7 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_11 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_hi_7, regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_hi_hi_14 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_11, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_11};
  wire [31:0]        regroupV0_hi_hi_hi_hi_lo_hi_14 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_14, regroupV0_hi_hi_hi_hi_lo_hi_lo_14};
  wire [63:0]        regroupV0_hi_hi_hi_hi_lo_14 = {regroupV0_hi_hi_hi_hi_lo_hi_14, regroupV0_hi_hi_hi_hi_lo_lo_14};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo_lo_3 = {regroupV0_hi_12[3847], regroupV0_hi_12[3843]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo_hi_3 = {regroupV0_hi_12[3855], regroupV0_hi_12[3851]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo_7 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo_hi_3, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi_lo_3 = {regroupV0_hi_12[3863], regroupV0_hi_12[3859]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi_hi_3 = {regroupV0_hi_12[3871], regroupV0_hi_12[3867]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi_7 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi_hi_3, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_11 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_hi_7, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo_lo_3 = {regroupV0_hi_12[3879], regroupV0_hi_12[3875]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo_hi_3 = {regroupV0_hi_12[3887], regroupV0_hi_12[3883]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo_7 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo_hi_3, regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi_lo_3 = {regroupV0_hi_12[3895], regroupV0_hi_12[3891]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi_hi_3 = {regroupV0_hi_12[3903], regroupV0_hi_12[3899]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi_7 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi_hi_3, regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_11 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_hi_7, regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_lo_lo_14 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_11, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo_lo_3 = {regroupV0_hi_12[3911], regroupV0_hi_12[3907]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo_hi_3 = {regroupV0_hi_12[3919], regroupV0_hi_12[3915]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo_7 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo_hi_3, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi_lo_3 = {regroupV0_hi_12[3927], regroupV0_hi_12[3923]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi_hi_3 = {regroupV0_hi_12[3935], regroupV0_hi_12[3931]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi_7 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi_hi_3, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_11 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_hi_7, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo_lo_3 = {regroupV0_hi_12[3943], regroupV0_hi_12[3939]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo_hi_3 = {regroupV0_hi_12[3951], regroupV0_hi_12[3947]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo_7 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo_hi_3, regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi_lo_3 = {regroupV0_hi_12[3959], regroupV0_hi_12[3955]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi_hi_3 = {regroupV0_hi_12[3967], regroupV0_hi_12[3963]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi_7 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_11 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_hi_7, regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_lo_hi_14 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_11, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_11};
  wire [31:0]        regroupV0_hi_hi_hi_hi_hi_lo_14 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_14, regroupV0_hi_hi_hi_hi_hi_lo_lo_14};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo_lo_3 = {regroupV0_hi_12[3975], regroupV0_hi_12[3971]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo_hi_3 = {regroupV0_hi_12[3983], regroupV0_hi_12[3979]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo_7 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo_hi_3, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi_lo_3 = {regroupV0_hi_12[3991], regroupV0_hi_12[3987]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi_hi_3 = {regroupV0_hi_12[3999], regroupV0_hi_12[3995]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi_7 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi_hi_3, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_11 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_hi_7, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo_lo_3 = {regroupV0_hi_12[4007], regroupV0_hi_12[4003]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo_hi_3 = {regroupV0_hi_12[4015], regroupV0_hi_12[4011]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo_7 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo_hi_3, regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi_lo_3 = {regroupV0_hi_12[4023], regroupV0_hi_12[4019]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi_hi_3 = {regroupV0_hi_12[4031], regroupV0_hi_12[4027]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi_7 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi_hi_3, regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_11 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_hi_7, regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_hi_lo_14 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_11, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo_lo_3 = {regroupV0_hi_12[4039], regroupV0_hi_12[4035]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo_hi_3 = {regroupV0_hi_12[4047], regroupV0_hi_12[4043]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo_7 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo_hi_3, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi_lo_3 = {regroupV0_hi_12[4055], regroupV0_hi_12[4051]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi_hi_3 = {regroupV0_hi_12[4063], regroupV0_hi_12[4059]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi_7 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi_hi_3, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_11 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_hi_7, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo_lo_3 = {regroupV0_hi_12[4071], regroupV0_hi_12[4067]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo_hi_3 = {regroupV0_hi_12[4079], regroupV0_hi_12[4075]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo_7 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo_hi_3, regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi_lo_3 = {regroupV0_hi_12[4087], regroupV0_hi_12[4083]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi_hi_3 = {regroupV0_hi_12[4095], regroupV0_hi_12[4091]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi_7 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_11 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_hi_7, regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_hi_hi_14 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_11, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_11};
  wire [31:0]        regroupV0_hi_hi_hi_hi_hi_hi_14 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_14, regroupV0_hi_hi_hi_hi_hi_hi_lo_14};
  wire [63:0]        regroupV0_hi_hi_hi_hi_hi_14 = {regroupV0_hi_hi_hi_hi_hi_hi_14, regroupV0_hi_hi_hi_hi_hi_lo_14};
  wire [127:0]       regroupV0_hi_hi_hi_hi_14 = {regroupV0_hi_hi_hi_hi_hi_14, regroupV0_hi_hi_hi_hi_lo_14};
  wire [255:0]       regroupV0_hi_hi_hi_14 = {regroupV0_hi_hi_hi_hi_14, regroupV0_hi_hi_hi_lo_14};
  wire [511:0]       regroupV0_hi_hi_14 = {regroupV0_hi_hi_hi_14, regroupV0_hi_hi_lo_14};
  wire [1023:0]      regroupV0_hi_16 = {regroupV0_hi_hi_14, regroupV0_hi_lo_14};
  wire [4095:0]      regroupV0_lo_17 = {regroupV0_hi_14, regroupV0_lo_14, regroupV0_hi_13, regroupV0_lo_13};
  wire [4095:0]      regroupV0_hi_17 = {regroupV0_hi_16, regroupV0_lo_16, regroupV0_hi_15, regroupV0_lo_15};
  wire [8191:0]      regroupV0_2 = {regroupV0_hi_17, regroupV0_lo_17};
  wire [3:0]         _v0SelectBySew_T = 4'h1 << laneMaskSewSelect_0;
  wire [2047:0]      v0SelectBySew = (_v0SelectBySew_T[0] ? regroupV0_0[2047:0] : 2048'h0) | (_v0SelectBySew_T[1] ? regroupV0_1[2047:0] : 2048'h0) | (_v0SelectBySew_T[2] ? regroupV0_2[2047:0] : 2048'h0);
  wire [63:0][31:0]  _GEN_127 =
    {{v0SelectBySew[2047:2016]},
     {v0SelectBySew[2015:1984]},
     {v0SelectBySew[1983:1952]},
     {v0SelectBySew[1951:1920]},
     {v0SelectBySew[1919:1888]},
     {v0SelectBySew[1887:1856]},
     {v0SelectBySew[1855:1824]},
     {v0SelectBySew[1823:1792]},
     {v0SelectBySew[1791:1760]},
     {v0SelectBySew[1759:1728]},
     {v0SelectBySew[1727:1696]},
     {v0SelectBySew[1695:1664]},
     {v0SelectBySew[1663:1632]},
     {v0SelectBySew[1631:1600]},
     {v0SelectBySew[1599:1568]},
     {v0SelectBySew[1567:1536]},
     {v0SelectBySew[1535:1504]},
     {v0SelectBySew[1503:1472]},
     {v0SelectBySew[1471:1440]},
     {v0SelectBySew[1439:1408]},
     {v0SelectBySew[1407:1376]},
     {v0SelectBySew[1375:1344]},
     {v0SelectBySew[1343:1312]},
     {v0SelectBySew[1311:1280]},
     {v0SelectBySew[1279:1248]},
     {v0SelectBySew[1247:1216]},
     {v0SelectBySew[1215:1184]},
     {v0SelectBySew[1183:1152]},
     {v0SelectBySew[1151:1120]},
     {v0SelectBySew[1119:1088]},
     {v0SelectBySew[1087:1056]},
     {v0SelectBySew[1055:1024]},
     {v0SelectBySew[1023:992]},
     {v0SelectBySew[991:960]},
     {v0SelectBySew[959:928]},
     {v0SelectBySew[927:896]},
     {v0SelectBySew[895:864]},
     {v0SelectBySew[863:832]},
     {v0SelectBySew[831:800]},
     {v0SelectBySew[799:768]},
     {v0SelectBySew[767:736]},
     {v0SelectBySew[735:704]},
     {v0SelectBySew[703:672]},
     {v0SelectBySew[671:640]},
     {v0SelectBySew[639:608]},
     {v0SelectBySew[607:576]},
     {v0SelectBySew[575:544]},
     {v0SelectBySew[543:512]},
     {v0SelectBySew[511:480]},
     {v0SelectBySew[479:448]},
     {v0SelectBySew[447:416]},
     {v0SelectBySew[415:384]},
     {v0SelectBySew[383:352]},
     {v0SelectBySew[351:320]},
     {v0SelectBySew[319:288]},
     {v0SelectBySew[287:256]},
     {v0SelectBySew[255:224]},
     {v0SelectBySew[223:192]},
     {v0SelectBySew[191:160]},
     {v0SelectBySew[159:128]},
     {v0SelectBySew[127:96]},
     {v0SelectBySew[95:64]},
     {v0SelectBySew[63:32]},
     {v0SelectBySew[31:0]}};
  wire [3:0]         _v0SelectBySew_T_9 = 4'h1 << laneMaskSewSelect_1;
  wire [2047:0]      v0SelectBySew_1 = (_v0SelectBySew_T_9[0] ? regroupV0_0[4095:2048] : 2048'h0) | (_v0SelectBySew_T_9[1] ? regroupV0_1[4095:2048] : 2048'h0) | (_v0SelectBySew_T_9[2] ? regroupV0_2[4095:2048] : 2048'h0);
  wire [63:0][31:0]  _GEN_128 =
    {{v0SelectBySew_1[2047:2016]},
     {v0SelectBySew_1[2015:1984]},
     {v0SelectBySew_1[1983:1952]},
     {v0SelectBySew_1[1951:1920]},
     {v0SelectBySew_1[1919:1888]},
     {v0SelectBySew_1[1887:1856]},
     {v0SelectBySew_1[1855:1824]},
     {v0SelectBySew_1[1823:1792]},
     {v0SelectBySew_1[1791:1760]},
     {v0SelectBySew_1[1759:1728]},
     {v0SelectBySew_1[1727:1696]},
     {v0SelectBySew_1[1695:1664]},
     {v0SelectBySew_1[1663:1632]},
     {v0SelectBySew_1[1631:1600]},
     {v0SelectBySew_1[1599:1568]},
     {v0SelectBySew_1[1567:1536]},
     {v0SelectBySew_1[1535:1504]},
     {v0SelectBySew_1[1503:1472]},
     {v0SelectBySew_1[1471:1440]},
     {v0SelectBySew_1[1439:1408]},
     {v0SelectBySew_1[1407:1376]},
     {v0SelectBySew_1[1375:1344]},
     {v0SelectBySew_1[1343:1312]},
     {v0SelectBySew_1[1311:1280]},
     {v0SelectBySew_1[1279:1248]},
     {v0SelectBySew_1[1247:1216]},
     {v0SelectBySew_1[1215:1184]},
     {v0SelectBySew_1[1183:1152]},
     {v0SelectBySew_1[1151:1120]},
     {v0SelectBySew_1[1119:1088]},
     {v0SelectBySew_1[1087:1056]},
     {v0SelectBySew_1[1055:1024]},
     {v0SelectBySew_1[1023:992]},
     {v0SelectBySew_1[991:960]},
     {v0SelectBySew_1[959:928]},
     {v0SelectBySew_1[927:896]},
     {v0SelectBySew_1[895:864]},
     {v0SelectBySew_1[863:832]},
     {v0SelectBySew_1[831:800]},
     {v0SelectBySew_1[799:768]},
     {v0SelectBySew_1[767:736]},
     {v0SelectBySew_1[735:704]},
     {v0SelectBySew_1[703:672]},
     {v0SelectBySew_1[671:640]},
     {v0SelectBySew_1[639:608]},
     {v0SelectBySew_1[607:576]},
     {v0SelectBySew_1[575:544]},
     {v0SelectBySew_1[543:512]},
     {v0SelectBySew_1[511:480]},
     {v0SelectBySew_1[479:448]},
     {v0SelectBySew_1[447:416]},
     {v0SelectBySew_1[415:384]},
     {v0SelectBySew_1[383:352]},
     {v0SelectBySew_1[351:320]},
     {v0SelectBySew_1[319:288]},
     {v0SelectBySew_1[287:256]},
     {v0SelectBySew_1[255:224]},
     {v0SelectBySew_1[223:192]},
     {v0SelectBySew_1[191:160]},
     {v0SelectBySew_1[159:128]},
     {v0SelectBySew_1[127:96]},
     {v0SelectBySew_1[95:64]},
     {v0SelectBySew_1[63:32]},
     {v0SelectBySew_1[31:0]}};
  wire [3:0]         _v0SelectBySew_T_18 = 4'h1 << laneMaskSewSelect_2;
  wire [2047:0]      v0SelectBySew_2 = (_v0SelectBySew_T_18[0] ? regroupV0_0[6143:4096] : 2048'h0) | (_v0SelectBySew_T_18[1] ? regroupV0_1[6143:4096] : 2048'h0) | (_v0SelectBySew_T_18[2] ? regroupV0_2[6143:4096] : 2048'h0);
  wire [63:0][31:0]  _GEN_129 =
    {{v0SelectBySew_2[2047:2016]},
     {v0SelectBySew_2[2015:1984]},
     {v0SelectBySew_2[1983:1952]},
     {v0SelectBySew_2[1951:1920]},
     {v0SelectBySew_2[1919:1888]},
     {v0SelectBySew_2[1887:1856]},
     {v0SelectBySew_2[1855:1824]},
     {v0SelectBySew_2[1823:1792]},
     {v0SelectBySew_2[1791:1760]},
     {v0SelectBySew_2[1759:1728]},
     {v0SelectBySew_2[1727:1696]},
     {v0SelectBySew_2[1695:1664]},
     {v0SelectBySew_2[1663:1632]},
     {v0SelectBySew_2[1631:1600]},
     {v0SelectBySew_2[1599:1568]},
     {v0SelectBySew_2[1567:1536]},
     {v0SelectBySew_2[1535:1504]},
     {v0SelectBySew_2[1503:1472]},
     {v0SelectBySew_2[1471:1440]},
     {v0SelectBySew_2[1439:1408]},
     {v0SelectBySew_2[1407:1376]},
     {v0SelectBySew_2[1375:1344]},
     {v0SelectBySew_2[1343:1312]},
     {v0SelectBySew_2[1311:1280]},
     {v0SelectBySew_2[1279:1248]},
     {v0SelectBySew_2[1247:1216]},
     {v0SelectBySew_2[1215:1184]},
     {v0SelectBySew_2[1183:1152]},
     {v0SelectBySew_2[1151:1120]},
     {v0SelectBySew_2[1119:1088]},
     {v0SelectBySew_2[1087:1056]},
     {v0SelectBySew_2[1055:1024]},
     {v0SelectBySew_2[1023:992]},
     {v0SelectBySew_2[991:960]},
     {v0SelectBySew_2[959:928]},
     {v0SelectBySew_2[927:896]},
     {v0SelectBySew_2[895:864]},
     {v0SelectBySew_2[863:832]},
     {v0SelectBySew_2[831:800]},
     {v0SelectBySew_2[799:768]},
     {v0SelectBySew_2[767:736]},
     {v0SelectBySew_2[735:704]},
     {v0SelectBySew_2[703:672]},
     {v0SelectBySew_2[671:640]},
     {v0SelectBySew_2[639:608]},
     {v0SelectBySew_2[607:576]},
     {v0SelectBySew_2[575:544]},
     {v0SelectBySew_2[543:512]},
     {v0SelectBySew_2[511:480]},
     {v0SelectBySew_2[479:448]},
     {v0SelectBySew_2[447:416]},
     {v0SelectBySew_2[415:384]},
     {v0SelectBySew_2[383:352]},
     {v0SelectBySew_2[351:320]},
     {v0SelectBySew_2[319:288]},
     {v0SelectBySew_2[287:256]},
     {v0SelectBySew_2[255:224]},
     {v0SelectBySew_2[223:192]},
     {v0SelectBySew_2[191:160]},
     {v0SelectBySew_2[159:128]},
     {v0SelectBySew_2[127:96]},
     {v0SelectBySew_2[95:64]},
     {v0SelectBySew_2[63:32]},
     {v0SelectBySew_2[31:0]}};
  wire [3:0]         _v0SelectBySew_T_27 = 4'h1 << laneMaskSewSelect_3;
  wire [2047:0]      v0SelectBySew_3 = (_v0SelectBySew_T_27[0] ? regroupV0_0[8191:6144] : 2048'h0) | (_v0SelectBySew_T_27[1] ? regroupV0_1[8191:6144] : 2048'h0) | (_v0SelectBySew_T_27[2] ? regroupV0_2[8191:6144] : 2048'h0);
  wire [63:0][31:0]  _GEN_130 =
    {{v0SelectBySew_3[2047:2016]},
     {v0SelectBySew_3[2015:1984]},
     {v0SelectBySew_3[1983:1952]},
     {v0SelectBySew_3[1951:1920]},
     {v0SelectBySew_3[1919:1888]},
     {v0SelectBySew_3[1887:1856]},
     {v0SelectBySew_3[1855:1824]},
     {v0SelectBySew_3[1823:1792]},
     {v0SelectBySew_3[1791:1760]},
     {v0SelectBySew_3[1759:1728]},
     {v0SelectBySew_3[1727:1696]},
     {v0SelectBySew_3[1695:1664]},
     {v0SelectBySew_3[1663:1632]},
     {v0SelectBySew_3[1631:1600]},
     {v0SelectBySew_3[1599:1568]},
     {v0SelectBySew_3[1567:1536]},
     {v0SelectBySew_3[1535:1504]},
     {v0SelectBySew_3[1503:1472]},
     {v0SelectBySew_3[1471:1440]},
     {v0SelectBySew_3[1439:1408]},
     {v0SelectBySew_3[1407:1376]},
     {v0SelectBySew_3[1375:1344]},
     {v0SelectBySew_3[1343:1312]},
     {v0SelectBySew_3[1311:1280]},
     {v0SelectBySew_3[1279:1248]},
     {v0SelectBySew_3[1247:1216]},
     {v0SelectBySew_3[1215:1184]},
     {v0SelectBySew_3[1183:1152]},
     {v0SelectBySew_3[1151:1120]},
     {v0SelectBySew_3[1119:1088]},
     {v0SelectBySew_3[1087:1056]},
     {v0SelectBySew_3[1055:1024]},
     {v0SelectBySew_3[1023:992]},
     {v0SelectBySew_3[991:960]},
     {v0SelectBySew_3[959:928]},
     {v0SelectBySew_3[927:896]},
     {v0SelectBySew_3[895:864]},
     {v0SelectBySew_3[863:832]},
     {v0SelectBySew_3[831:800]},
     {v0SelectBySew_3[799:768]},
     {v0SelectBySew_3[767:736]},
     {v0SelectBySew_3[735:704]},
     {v0SelectBySew_3[703:672]},
     {v0SelectBySew_3[671:640]},
     {v0SelectBySew_3[639:608]},
     {v0SelectBySew_3[607:576]},
     {v0SelectBySew_3[575:544]},
     {v0SelectBySew_3[543:512]},
     {v0SelectBySew_3[511:480]},
     {v0SelectBySew_3[479:448]},
     {v0SelectBySew_3[447:416]},
     {v0SelectBySew_3[415:384]},
     {v0SelectBySew_3[383:352]},
     {v0SelectBySew_3[351:320]},
     {v0SelectBySew_3[319:288]},
     {v0SelectBySew_3[287:256]},
     {v0SelectBySew_3[255:224]},
     {v0SelectBySew_3[223:192]},
     {v0SelectBySew_3[191:160]},
     {v0SelectBySew_3[159:128]},
     {v0SelectBySew_3[127:96]},
     {v0SelectBySew_3[95:64]},
     {v0SelectBySew_3[63:32]},
     {v0SelectBySew_3[31:0]}};
  wire [3:0]         intLMULInput = 4'h1 << instReq_bits_vlmul[1:0];
  wire [15:0]        _dataPosition_T_1 = {3'h0, instReq_bits_readFromScala[12:0]} << instReq_bits_sew;
  wire [12:0]        dataPosition = _dataPosition_T_1[12:0];
  wire [3:0]         _sewOHInput_T = 4'h1 << instReq_bits_sew;
  wire [2:0]         sewOHInput = _sewOHInput_T[2:0];
  wire [1:0]         dataOffset = {dataPosition[1] & (|(sewOHInput[1:0])), dataPosition[0] & sewOHInput[0]};
  wire [1:0]         accessLane = dataPosition[3:2];
  wire [8:0]         dataGroup = dataPosition[12:4];
  wire [5:0]         offset = dataGroup[5:0];
  wire [2:0]         accessRegGrowth = dataGroup[8:6];
  wire [2:0]         reallyGrowth = accessRegGrowth;
  wire [7:0]         decimalProportion = {offset, accessLane};
  wire [2:0]         decimal = decimalProportion[7:5];
  wire               notNeedRead = |{instReq_bits_vlmul[2] & decimal >= intLMULInput[3:1] | ~(instReq_bits_vlmul[2]) & {1'h0, accessRegGrowth} >= intLMULInput, instReq_bits_readFromScala[31:13]};
  reg  [1:0]         gatherReadState;
  wire               gatherSRead = gatherReadState == 2'h1;
  wire               gatherWaiteRead = gatherReadState == 2'h2;
  assign gatherResponse = &gatherReadState;
  wire               gatherData_valid_0 = gatherResponse;
  reg  [1:0]         gatherDatOffset;
  reg  [1:0]         gatherLane;
  reg  [5:0]         gatherOffset;
  reg  [2:0]         gatherGrowth;
  reg  [2:0]         instReg_instructionIndex;
  wire [2:0]         exeResp_0_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_1_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_2_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_3_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_0_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_1_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_2_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_3_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         writeRequest_0_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_1_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_2_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_3_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_0_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_1_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_2_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_3_enq_bits_index = instReg_instructionIndex;
  reg                instReg_decodeResult_specialSlot;
  reg  [4:0]         instReg_decodeResult_topUop;
  reg                instReg_decodeResult_popCount;
  reg                instReg_decodeResult_ffo;
  reg                instReg_decodeResult_average;
  reg                instReg_decodeResult_reverse;
  reg                instReg_decodeResult_dontNeedExecuteInLane;
  reg                instReg_decodeResult_scheduler;
  reg                instReg_decodeResult_sReadVD;
  reg                instReg_decodeResult_vtype;
  reg                instReg_decodeResult_sWrite;
  reg                instReg_decodeResult_crossRead;
  reg                instReg_decodeResult_crossWrite;
  reg                instReg_decodeResult_maskUnit;
  reg                instReg_decodeResult_special;
  reg                instReg_decodeResult_saturate;
  reg                instReg_decodeResult_vwmacc;
  reg                instReg_decodeResult_readOnly;
  reg                instReg_decodeResult_maskSource;
  reg                instReg_decodeResult_maskDestination;
  reg                instReg_decodeResult_maskLogic;
  reg  [3:0]         instReg_decodeResult_uop;
  reg                instReg_decodeResult_iota;
  reg                instReg_decodeResult_mv;
  reg                instReg_decodeResult_extend;
  reg                instReg_decodeResult_unOrderWrite;
  reg                instReg_decodeResult_compress;
  reg                instReg_decodeResult_gather16;
  reg                instReg_decodeResult_gather;
  reg                instReg_decodeResult_slid;
  reg                instReg_decodeResult_targetRd;
  reg                instReg_decodeResult_widenReduce;
  reg                instReg_decodeResult_red;
  reg                instReg_decodeResult_nr;
  reg                instReg_decodeResult_itype;
  reg                instReg_decodeResult_unsigned1;
  reg                instReg_decodeResult_unsigned0;
  reg                instReg_decodeResult_other;
  reg                instReg_decodeResult_multiCycle;
  reg                instReg_decodeResult_divider;
  reg                instReg_decodeResult_multiplier;
  reg                instReg_decodeResult_shift;
  reg                instReg_decodeResult_adder;
  reg                instReg_decodeResult_logic;
  reg  [31:0]        instReg_readFromScala;
  reg  [1:0]         instReg_sew;
  reg  [2:0]         instReg_vlmul;
  reg                instReg_maskType;
  reg  [2:0]         instReg_vxrm;
  reg  [4:0]         instReg_vs2;
  reg  [4:0]         instReg_vs1;
  reg  [4:0]         instReg_vd;
  wire [4:0]         writeRequest_0_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_1_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_2_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_3_writeData_vd = instReg_vd;
  reg  [13:0]        instReg_vl;
  wire [13:0]        reduceLastDataNeed_byteForVl = instReg_vl;
  wire               enqMvRD = instReq_bits_decodeResult_topUop == 5'hB;
  reg                instVlValid;
  wire               gatherRequestFire = gatherReadState == 2'h0 & gatherRead & ~instVlValid;
  wire               viotaReq = instReq_bits_decodeResult_topUop == 5'h8;
  reg                readVS1Reg_dataValid;
  reg                readVS1Reg_requestSend;
  reg                readVS1Reg_sendToExecution;
  reg  [31:0]        readVS1Reg_data;
  reg  [8:0]         readVS1Reg_readIndex;
  wire [3:0]         _sew1H_T = 4'h1 << instReg_sew;
  wire [2:0]         sew1H = _sew1H_T[2:0];
  wire [3:0]         unitType = 4'h1 << instReg_decodeResult_topUop[4:3];
  wire [3:0]         subType = 4'h1 << instReg_decodeResult_topUop[2:1];
  wire               readType = unitType[0];
  wire               gather16 = instReg_decodeResult_topUop == 5'h5;
  wire               maskDestinationType = instReg_decodeResult_topUop == 5'h18;
  wire               compress = instReg_decodeResult_topUop[4:1] == 4'h4;
  wire               viota = instReg_decodeResult_topUop == 5'h8;
  wire               mv = instReg_decodeResult_topUop[4:1] == 4'h5;
  wire               mvRd = instReg_decodeResult_topUop == 5'hB;
  wire               mvVd = instReg_decodeResult_topUop == 5'hA;
  wire               orderReduce = {instReg_decodeResult_topUop[4:2], instReg_decodeResult_topUop[0]} == 4'hB;
  wire               ffo = instReg_decodeResult_topUop[4:1] == 4'h7;
  wire               extendType = unitType[3] & (subType[2] | subType[1]);
  wire               readValid = readType & instVlValid;
  wire               noSource = mv | viota;
  wire               allGroupExecute = maskDestinationType | unitType[2] | compress | ffo;
  wire               useDefaultSew = readType & ~gather16;
  wire [1:0]         _dataSplitSew_T_11 = useDefaultSew ? instReg_sew : 2'h0;
  wire [1:0]         dataSplitSew = {_dataSplitSew_T_11[1], _dataSplitSew_T_11[0] | unitType[3] & subType[1] | gather16} | {allGroupExecute, 1'h0};
  wire               sourceDataUseDefaultSew = ~(unitType[3] | gather16);
  wire [1:0]         _sourceDataEEW_T_6 = (sourceDataUseDefaultSew ? instReg_sew : 2'h0) | (unitType[3] ? instReg_sew >> subType[2:1] : 2'h0);
  wire [1:0]         sourceDataEEW = {_sourceDataEEW_T_6[1], _sourceDataEEW_T_6[0] | gather16};
  wire [3:0]         executeIndexGrowth = 4'h1 << dataSplitSew;
  wire [1:0]         lastExecuteIndex = {2{executeIndexGrowth[0]}} | {executeIndexGrowth[1], 1'h0};
  wire [3:0]         _sourceDataEEW1H_T = 4'h1 << sourceDataEEW;
  wire [2:0]         sourceDataEEW1H = _sourceDataEEW1H_T[2:0];
  wire [12:0]        lastElementIndex = instReg_vl[12:0] - {12'h0, |instReg_vl};
  wire [12:0]        processingVl_lastByteIndex = lastElementIndex;
  wire               maskFormatSource = ffo | maskDestinationType;
  wire [3:0]         processingVl_lastGroupRemaining = processingVl_lastByteIndex[3:0];
  wire [8:0]         processingVl_0_1 = processingVl_lastByteIndex[12:4];
  wire [1:0]         processingVl_lastLaneIndex = processingVl_lastGroupRemaining[3:2];
  wire [3:0]         _processingVl_lastGroupDataNeed_T = 4'h1 << processingVl_lastLaneIndex;
  wire [2:0]         _GEN_131 = _processingVl_lastGroupDataNeed_T[2:0] | _processingVl_lastGroupDataNeed_T[3:1];
  wire [3:0]         processingVl_0_2 = {_processingVl_lastGroupDataNeed_T[3], _GEN_131[2], _GEN_131[1:0] | {_processingVl_lastGroupDataNeed_T[3], _GEN_131[2]}};
  wire [13:0]        processingVl_lastByteIndex_1 = {lastElementIndex, 1'h0};
  wire [3:0]         processingVl_lastGroupRemaining_1 = processingVl_lastByteIndex_1[3:0];
  wire [9:0]         processingVl_1_1 = processingVl_lastByteIndex_1[13:4];
  wire [1:0]         processingVl_lastLaneIndex_1 = processingVl_lastGroupRemaining_1[3:2];
  wire [3:0]         _processingVl_lastGroupDataNeed_T_5 = 4'h1 << processingVl_lastLaneIndex_1;
  wire [2:0]         _GEN_132 = _processingVl_lastGroupDataNeed_T_5[2:0] | _processingVl_lastGroupDataNeed_T_5[3:1];
  wire [3:0]         processingVl_1_2 = {_processingVl_lastGroupDataNeed_T_5[3], _GEN_132[2], _GEN_132[1:0] | {_processingVl_lastGroupDataNeed_T_5[3], _GEN_132[2]}};
  wire [14:0]        processingVl_lastByteIndex_2 = {lastElementIndex, 2'h0};
  wire [3:0]         processingVl_lastGroupRemaining_2 = processingVl_lastByteIndex_2[3:0];
  wire [10:0]        processingVl_2_1 = processingVl_lastByteIndex_2[14:4];
  wire [1:0]         processingVl_lastLaneIndex_2 = processingVl_lastGroupRemaining_2[3:2];
  wire [3:0]         _processingVl_lastGroupDataNeed_T_10 = 4'h1 << processingVl_lastLaneIndex_2;
  wire [2:0]         _GEN_133 = _processingVl_lastGroupDataNeed_T_10[2:0] | _processingVl_lastGroupDataNeed_T_10[3:1];
  wire [3:0]         processingVl_2_2 = {_processingVl_lastGroupDataNeed_T_10[3], _GEN_133[2], _GEN_133[1:0] | {_processingVl_lastGroupDataNeed_T_10[3], _GEN_133[2]}};
  wire [6:0]         processingMaskVl_lastGroupRemaining = lastElementIndex[6:0];
  wire [6:0]         elementTailForMaskDestination = lastElementIndex[6:0];
  wire               processingMaskVl_lastGroupMisAlign = |processingMaskVl_lastGroupRemaining;
  wire [5:0]         processingMaskVl_0_1 = lastElementIndex[12:7];
  wire [1:0]         processingMaskVl_lastLaneIndex = processingMaskVl_lastGroupRemaining[6:5] - {1'h0, processingMaskVl_lastGroupRemaining[4:0] == 5'h0};
  wire [3:0]         _processingMaskVl_dataNeedForPL_T = 4'h1 << processingMaskVl_lastLaneIndex;
  wire [2:0]         _GEN_134 = _processingMaskVl_dataNeedForPL_T[2:0] | _processingMaskVl_dataNeedForPL_T[3:1];
  wire [3:0]         processingMaskVl_dataNeedForPL = {_processingMaskVl_dataNeedForPL_T[3], _GEN_134[2], _GEN_134[1:0] | {_processingMaskVl_dataNeedForPL_T[3], _GEN_134[2]}};
  wire               processingMaskVl_dataNeedForNPL_misAlign = |(processingMaskVl_lastGroupRemaining[1:0]);
  wire [5:0]         processingMaskVl_dataNeedForNPL_datapathSize = {1'h0, processingMaskVl_lastGroupRemaining[6:2]} + {5'h0, processingMaskVl_dataNeedForNPL_misAlign};
  wire               processingMaskVl_dataNeedForNPL_allNeed = |(processingMaskVl_dataNeedForNPL_datapathSize[5:2]);
  wire [1:0]         processingMaskVl_dataNeedForNPL_lastLaneIndex = processingMaskVl_dataNeedForNPL_datapathSize[1:0];
  wire [3:0]         _processingMaskVl_dataNeedForNPL_dataNeed_T = 4'h1 << processingMaskVl_dataNeedForNPL_lastLaneIndex;
  wire [3:0]         _processingMaskVl_dataNeedForNPL_dataNeed_T_3 = _processingMaskVl_dataNeedForNPL_dataNeed_T | {_processingMaskVl_dataNeedForNPL_dataNeed_T[2:0], 1'h0};
  wire [3:0]         processingMaskVl_dataNeedForNPL_dataNeed = ~(_processingMaskVl_dataNeedForNPL_dataNeed_T_3 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_3[1:0], 2'h0}) | {4{processingMaskVl_dataNeedForNPL_allNeed}};
  wire               processingMaskVl_dataNeedForNPL_misAlign_1 = processingMaskVl_lastGroupRemaining[0];
  wire [6:0]         processingMaskVl_dataNeedForNPL_datapathSize_1 = {1'h0, processingMaskVl_lastGroupRemaining[6:1]} + {6'h0, processingMaskVl_dataNeedForNPL_misAlign_1};
  wire               processingMaskVl_dataNeedForNPL_allNeed_1 = |(processingMaskVl_dataNeedForNPL_datapathSize_1[6:2]);
  wire [1:0]         processingMaskVl_dataNeedForNPL_lastLaneIndex_1 = processingMaskVl_dataNeedForNPL_datapathSize_1[1:0];
  wire [3:0]         _processingMaskVl_dataNeedForNPL_dataNeed_T_10 = 4'h1 << processingMaskVl_dataNeedForNPL_lastLaneIndex_1;
  wire [3:0]         _processingMaskVl_dataNeedForNPL_dataNeed_T_13 = _processingMaskVl_dataNeedForNPL_dataNeed_T_10 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_10[2:0], 1'h0};
  wire [3:0]         processingMaskVl_dataNeedForNPL_dataNeed_1 = ~(_processingMaskVl_dataNeedForNPL_dataNeed_T_13 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_13[1:0], 2'h0}) | {4{processingMaskVl_dataNeedForNPL_allNeed_1}};
  wire [7:0]         processingMaskVl_dataNeedForNPL_datapathSize_2 = {1'h0, processingMaskVl_lastGroupRemaining};
  wire               processingMaskVl_dataNeedForNPL_allNeed_2 = |(processingMaskVl_dataNeedForNPL_datapathSize_2[7:2]);
  wire [1:0]         processingMaskVl_dataNeedForNPL_lastLaneIndex_2 = processingMaskVl_dataNeedForNPL_datapathSize_2[1:0];
  wire [3:0]         _processingMaskVl_dataNeedForNPL_dataNeed_T_20 = 4'h1 << processingMaskVl_dataNeedForNPL_lastLaneIndex_2;
  wire [3:0]         _processingMaskVl_dataNeedForNPL_dataNeed_T_23 = _processingMaskVl_dataNeedForNPL_dataNeed_T_20 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_20[2:0], 1'h0};
  wire [3:0]         processingMaskVl_dataNeedForNPL_dataNeed_2 = ~(_processingMaskVl_dataNeedForNPL_dataNeed_T_23 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_23[1:0], 2'h0}) | {4{processingMaskVl_dataNeedForNPL_allNeed_2}};
  wire [3:0]         processingMaskVl_dataNeedForNPL =
    (sew1H[0] ? processingMaskVl_dataNeedForNPL_dataNeed : 4'h0) | (sew1H[1] ? processingMaskVl_dataNeedForNPL_dataNeed_1 : 4'h0) | (sew1H[2] ? processingMaskVl_dataNeedForNPL_dataNeed_2 : 4'h0);
  wire [3:0]         processingMaskVl_0_2 = ffo ? processingMaskVl_dataNeedForPL : processingMaskVl_dataNeedForNPL;
  wire               reduceLastDataNeed_vlMSB = |(reduceLastDataNeed_byteForVl[13:4]);
  wire [3:0]         reduceLastDataNeed_vlLSB = instReg_vl[3:0];
  wire [3:0]         reduceLastDataNeed_vlLSB_1 = instReg_vl[3:0];
  wire [3:0]         reduceLastDataNeed_vlLSB_2 = instReg_vl[3:0];
  wire [1:0]         reduceLastDataNeed_lsbDSize = reduceLastDataNeed_vlLSB[3:2] - {1'h0, reduceLastDataNeed_vlLSB[1:0] == 2'h0};
  wire [3:0]         _reduceLastDataNeed_T = 4'h1 << reduceLastDataNeed_lsbDSize;
  wire [2:0]         _GEN_135 = _reduceLastDataNeed_T[2:0] | _reduceLastDataNeed_T[3:1];
  wire [14:0]        reduceLastDataNeed_byteForVl_1 = {instReg_vl, 1'h0};
  wire               reduceLastDataNeed_vlMSB_1 = |(reduceLastDataNeed_byteForVl_1[14:4]);
  wire [1:0]         reduceLastDataNeed_lsbDSize_1 = reduceLastDataNeed_vlLSB_1[3:2] - {1'h0, reduceLastDataNeed_vlLSB_1[1:0] == 2'h0};
  wire [3:0]         _reduceLastDataNeed_T_8 = 4'h1 << reduceLastDataNeed_lsbDSize_1;
  wire [2:0]         _GEN_136 = _reduceLastDataNeed_T_8[2:0] | _reduceLastDataNeed_T_8[3:1];
  wire [15:0]        reduceLastDataNeed_byteForVl_2 = {instReg_vl, 2'h0};
  wire               reduceLastDataNeed_vlMSB_2 = |(reduceLastDataNeed_byteForVl_2[15:4]);
  wire [1:0]         reduceLastDataNeed_lsbDSize_2 = reduceLastDataNeed_vlLSB_2[3:2] - {1'h0, reduceLastDataNeed_vlLSB_2[1:0] == 2'h0};
  wire [3:0]         _reduceLastDataNeed_T_16 = 4'h1 << reduceLastDataNeed_lsbDSize_2;
  wire [2:0]         _GEN_137 = _reduceLastDataNeed_T_16[2:0] | _reduceLastDataNeed_T_16[3:1];
  wire [3:0]         reduceLastDataNeed =
    (sew1H[0] ? {_reduceLastDataNeed_T[3], _GEN_135[2], _GEN_135[1:0] | {_reduceLastDataNeed_T[3], _GEN_135[2]}} | {4{reduceLastDataNeed_vlMSB}} : 4'h0)
    | (sew1H[1] ? {_reduceLastDataNeed_T_8[3], _GEN_136[2], _GEN_136[1:0] | {_reduceLastDataNeed_T_8[3], _GEN_136[2]}} | {4{reduceLastDataNeed_vlMSB_1}} : 4'h0)
    | (sew1H[2] ? {_reduceLastDataNeed_T_16[3], _GEN_137[2], _GEN_137[1:0] | {_reduceLastDataNeed_T_16[3], _GEN_137[2]}} | {4{reduceLastDataNeed_vlMSB_2}} : 4'h0);
  wire [1:0]         dataSourceSew = unitType[3] ? instReg_sew - instReg_decodeResult_topUop[2:1] : gather16 ? 2'h1 : instReg_sew;
  wire [3:0]         _dataSourceSew1H_T = 4'h1 << dataSourceSew;
  wire [2:0]         dataSourceSew1H = _dataSourceSew1H_T[2:0];
  wire               unorderReduce = ~orderReduce & unitType[2];
  wire               normalFormat = ~maskFormatSource & ~unorderReduce & ~mv;
  wire [10:0]        lastGroupForInstruction =
    {1'h0, {1'h0, {3'h0, maskFormatSource ? processingMaskVl_0_1 : 6'h0} | (normalFormat & dataSourceSew1H[0] ? processingVl_0_1 : 9'h0)} | (normalFormat & dataSourceSew1H[1] ? processingVl_1_1 : 10'h0)}
    | (normalFormat & dataSourceSew1H[2] ? processingVl_2_1 : 11'h0);
  wire [7:0]         popDataNeed_dataPathGroups = lastElementIndex[12:5];
  wire [1:0]         popDataNeed_lastLaneIndex = popDataNeed_dataPathGroups[1:0];
  wire               popDataNeed_lagerThanDLen = |(popDataNeed_dataPathGroups[7:2]);
  wire [3:0]         _popDataNeed_T = 4'h1 << popDataNeed_lastLaneIndex;
  wire [2:0]         _GEN_138 = _popDataNeed_T[2:0] | _popDataNeed_T[3:1];
  wire [3:0]         popDataNeed = {_popDataNeed_T[3], _GEN_138[2], _GEN_138[1:0] | {_popDataNeed_T[3], _GEN_138[2]}} | {4{popDataNeed_lagerThanDLen}};
  wire [3:0]         lastGroupDataNeed =
    (unorderReduce & instReg_decodeResult_popCount ? popDataNeed : 4'h0) | (unorderReduce & ~instReg_decodeResult_popCount ? reduceLastDataNeed : 4'h0) | (maskFormatSource ? processingMaskVl_0_2 : 4'h0)
    | (normalFormat & dataSourceSew1H[0] ? processingVl_0_2 : 4'h0) | (normalFormat & dataSourceSew1H[1] ? processingVl_1_2 : 4'h0) | (normalFormat & dataSourceSew1H[2] ? processingVl_2_2 : 4'h0);
  wire [3:0]         exeRequestQueue_queue_dataIn_lo = {exeRequestQueue_0_enq_bits_index, exeRequestQueue_0_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi = {exeRequestQueue_0_enq_bits_source1, exeRequestQueue_0_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn = {exeRequestQueue_queue_dataIn_hi, exeRequestQueue_queue_dataIn_lo};
  wire               exeRequestQueue_queue_dataOut_ffo = _exeRequestQueue_queue_fifo_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_index = _exeRequestQueue_queue_fifo_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_source2 = _exeRequestQueue_queue_fifo_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_source1 = _exeRequestQueue_queue_fifo_data_out[67:36];
  wire               exeRequestQueue_0_enq_ready = ~_exeRequestQueue_queue_fifo_full;
  wire               exeRequestQueue_0_deq_ready;
  wire               exeRequestQueue_0_deq_valid = ~_exeRequestQueue_queue_fifo_empty | exeRequestQueue_0_enq_valid;
  wire [31:0]        exeRequestQueue_0_deq_bits_source1 = _exeRequestQueue_queue_fifo_empty ? exeRequestQueue_0_enq_bits_source1 : exeRequestQueue_queue_dataOut_source1;
  wire [31:0]        exeRequestQueue_0_deq_bits_source2 = _exeRequestQueue_queue_fifo_empty ? exeRequestQueue_0_enq_bits_source2 : exeRequestQueue_queue_dataOut_source2;
  wire [2:0]         exeRequestQueue_0_deq_bits_index = _exeRequestQueue_queue_fifo_empty ? exeRequestQueue_0_enq_bits_index : exeRequestQueue_queue_dataOut_index;
  wire               exeRequestQueue_0_deq_bits_ffo = _exeRequestQueue_queue_fifo_empty ? exeRequestQueue_0_enq_bits_ffo : exeRequestQueue_queue_dataOut_ffo;
  wire               tokenIO_0_maskRequestRelease_0 = exeRequestQueue_0_deq_ready & exeRequestQueue_0_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_1 = {exeRequestQueue_1_enq_bits_index, exeRequestQueue_1_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_1 = {exeRequestQueue_1_enq_bits_source1, exeRequestQueue_1_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_1 = {exeRequestQueue_queue_dataIn_hi_1, exeRequestQueue_queue_dataIn_lo_1};
  wire               exeRequestQueue_queue_dataOut_1_ffo = _exeRequestQueue_queue_fifo_1_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_1_index = _exeRequestQueue_queue_fifo_1_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_1_source2 = _exeRequestQueue_queue_fifo_1_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_1_source1 = _exeRequestQueue_queue_fifo_1_data_out[67:36];
  wire               exeRequestQueue_1_enq_ready = ~_exeRequestQueue_queue_fifo_1_full;
  wire               exeRequestQueue_1_deq_ready;
  wire               exeRequestQueue_1_deq_valid = ~_exeRequestQueue_queue_fifo_1_empty | exeRequestQueue_1_enq_valid;
  wire [31:0]        exeRequestQueue_1_deq_bits_source1 = _exeRequestQueue_queue_fifo_1_empty ? exeRequestQueue_1_enq_bits_source1 : exeRequestQueue_queue_dataOut_1_source1;
  wire [31:0]        exeRequestQueue_1_deq_bits_source2 = _exeRequestQueue_queue_fifo_1_empty ? exeRequestQueue_1_enq_bits_source2 : exeRequestQueue_queue_dataOut_1_source2;
  wire [2:0]         exeRequestQueue_1_deq_bits_index = _exeRequestQueue_queue_fifo_1_empty ? exeRequestQueue_1_enq_bits_index : exeRequestQueue_queue_dataOut_1_index;
  wire               exeRequestQueue_1_deq_bits_ffo = _exeRequestQueue_queue_fifo_1_empty ? exeRequestQueue_1_enq_bits_ffo : exeRequestQueue_queue_dataOut_1_ffo;
  wire               tokenIO_1_maskRequestRelease_0 = exeRequestQueue_1_deq_ready & exeRequestQueue_1_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_2 = {exeRequestQueue_2_enq_bits_index, exeRequestQueue_2_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_2 = {exeRequestQueue_2_enq_bits_source1, exeRequestQueue_2_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_2 = {exeRequestQueue_queue_dataIn_hi_2, exeRequestQueue_queue_dataIn_lo_2};
  wire               exeRequestQueue_queue_dataOut_2_ffo = _exeRequestQueue_queue_fifo_2_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_2_index = _exeRequestQueue_queue_fifo_2_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_2_source2 = _exeRequestQueue_queue_fifo_2_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_2_source1 = _exeRequestQueue_queue_fifo_2_data_out[67:36];
  wire               exeRequestQueue_2_enq_ready = ~_exeRequestQueue_queue_fifo_2_full;
  wire               exeRequestQueue_2_deq_ready;
  wire               exeRequestQueue_2_deq_valid = ~_exeRequestQueue_queue_fifo_2_empty | exeRequestQueue_2_enq_valid;
  wire [31:0]        exeRequestQueue_2_deq_bits_source1 = _exeRequestQueue_queue_fifo_2_empty ? exeRequestQueue_2_enq_bits_source1 : exeRequestQueue_queue_dataOut_2_source1;
  wire [31:0]        exeRequestQueue_2_deq_bits_source2 = _exeRequestQueue_queue_fifo_2_empty ? exeRequestQueue_2_enq_bits_source2 : exeRequestQueue_queue_dataOut_2_source2;
  wire [2:0]         exeRequestQueue_2_deq_bits_index = _exeRequestQueue_queue_fifo_2_empty ? exeRequestQueue_2_enq_bits_index : exeRequestQueue_queue_dataOut_2_index;
  wire               exeRequestQueue_2_deq_bits_ffo = _exeRequestQueue_queue_fifo_2_empty ? exeRequestQueue_2_enq_bits_ffo : exeRequestQueue_queue_dataOut_2_ffo;
  wire               tokenIO_2_maskRequestRelease_0 = exeRequestQueue_2_deq_ready & exeRequestQueue_2_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_3 = {exeRequestQueue_3_enq_bits_index, exeRequestQueue_3_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_3 = {exeRequestQueue_3_enq_bits_source1, exeRequestQueue_3_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_3 = {exeRequestQueue_queue_dataIn_hi_3, exeRequestQueue_queue_dataIn_lo_3};
  wire               exeRequestQueue_queue_dataOut_3_ffo = _exeRequestQueue_queue_fifo_3_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_3_index = _exeRequestQueue_queue_fifo_3_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_3_source2 = _exeRequestQueue_queue_fifo_3_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_3_source1 = _exeRequestQueue_queue_fifo_3_data_out[67:36];
  wire               exeRequestQueue_3_enq_ready = ~_exeRequestQueue_queue_fifo_3_full;
  wire               exeRequestQueue_3_deq_ready;
  wire               exeRequestQueue_3_deq_valid = ~_exeRequestQueue_queue_fifo_3_empty | exeRequestQueue_3_enq_valid;
  wire [31:0]        exeRequestQueue_3_deq_bits_source1 = _exeRequestQueue_queue_fifo_3_empty ? exeRequestQueue_3_enq_bits_source1 : exeRequestQueue_queue_dataOut_3_source1;
  wire [31:0]        exeRequestQueue_3_deq_bits_source2 = _exeRequestQueue_queue_fifo_3_empty ? exeRequestQueue_3_enq_bits_source2 : exeRequestQueue_queue_dataOut_3_source2;
  wire [2:0]         exeRequestQueue_3_deq_bits_index = _exeRequestQueue_queue_fifo_3_empty ? exeRequestQueue_3_enq_bits_index : exeRequestQueue_queue_dataOut_3_index;
  wire               exeRequestQueue_3_deq_bits_ffo = _exeRequestQueue_queue_fifo_3_empty ? exeRequestQueue_3_enq_bits_ffo : exeRequestQueue_queue_dataOut_3_ffo;
  wire               tokenIO_3_maskRequestRelease_0 = exeRequestQueue_3_deq_ready & exeRequestQueue_3_deq_valid;
  reg                exeReqReg_0_valid;
  reg  [31:0]        exeReqReg_0_bits_source1;
  reg  [31:0]        exeReqReg_0_bits_source2;
  reg  [2:0]         exeReqReg_0_bits_index;
  reg                exeReqReg_0_bits_ffo;
  reg                exeReqReg_1_valid;
  reg  [31:0]        exeReqReg_1_bits_source1;
  reg  [31:0]        exeReqReg_1_bits_source2;
  reg  [2:0]         exeReqReg_1_bits_index;
  reg                exeReqReg_1_bits_ffo;
  reg                exeReqReg_2_valid;
  reg  [31:0]        exeReqReg_2_bits_source1;
  reg  [31:0]        exeReqReg_2_bits_source2;
  reg  [2:0]         exeReqReg_2_bits_index;
  reg                exeReqReg_2_bits_ffo;
  reg                exeReqReg_3_valid;
  reg  [31:0]        exeReqReg_3_bits_source1;
  reg  [31:0]        exeReqReg_3_bits_source2;
  reg  [2:0]         exeReqReg_3_bits_index;
  reg                exeReqReg_3_bits_ffo;
  reg  [9:0]         requestCounter;
  wire [10:0]        _GEN_139 = {1'h0, requestCounter};
  wire               counterValid = _GEN_139 <= lastGroupForInstruction;
  wire               lastGroup = _GEN_139 == lastGroupForInstruction | ~orderReduce & unitType[2] | mv;
  wire [127:0]       slideAddressGen_slideMaskInput_lo_lo_lo_lo_lo_lo = {slideAddressGen_slideMaskInput_lo_lo_lo_lo_lo_lo_hi, slideAddressGen_slideMaskInput_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_lo_lo_lo_lo_hi = {slideAddressGen_slideMaskInput_lo_lo_lo_lo_lo_hi_hi, slideAddressGen_slideMaskInput_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_lo_lo_lo_lo_lo = {slideAddressGen_slideMaskInput_lo_lo_lo_lo_lo_hi, slideAddressGen_slideMaskInput_lo_lo_lo_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_lo_lo_lo_hi_lo = {slideAddressGen_slideMaskInput_lo_lo_lo_lo_hi_lo_hi, slideAddressGen_slideMaskInput_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_lo_lo_lo_hi_hi = {slideAddressGen_slideMaskInput_lo_lo_lo_lo_hi_hi_hi, slideAddressGen_slideMaskInput_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_lo_lo_lo_lo_hi = {slideAddressGen_slideMaskInput_lo_lo_lo_lo_hi_hi, slideAddressGen_slideMaskInput_lo_lo_lo_lo_hi_lo};
  wire [511:0]       slideAddressGen_slideMaskInput_lo_lo_lo_lo = {slideAddressGen_slideMaskInput_lo_lo_lo_lo_hi, slideAddressGen_slideMaskInput_lo_lo_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_lo_lo_hi_lo_lo = {slideAddressGen_slideMaskInput_lo_lo_lo_hi_lo_lo_hi, slideAddressGen_slideMaskInput_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_lo_lo_hi_lo_hi = {slideAddressGen_slideMaskInput_lo_lo_lo_hi_lo_hi_hi, slideAddressGen_slideMaskInput_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_lo_lo_lo_hi_lo = {slideAddressGen_slideMaskInput_lo_lo_lo_hi_lo_hi, slideAddressGen_slideMaskInput_lo_lo_lo_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_lo_lo_hi_hi_lo = {slideAddressGen_slideMaskInput_lo_lo_lo_hi_hi_lo_hi, slideAddressGen_slideMaskInput_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_lo_lo_hi_hi_hi = {slideAddressGen_slideMaskInput_lo_lo_lo_hi_hi_hi_hi, slideAddressGen_slideMaskInput_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_lo_lo_lo_hi_hi = {slideAddressGen_slideMaskInput_lo_lo_lo_hi_hi_hi, slideAddressGen_slideMaskInput_lo_lo_lo_hi_hi_lo};
  wire [511:0]       slideAddressGen_slideMaskInput_lo_lo_lo_hi = {slideAddressGen_slideMaskInput_lo_lo_lo_hi_hi, slideAddressGen_slideMaskInput_lo_lo_lo_hi_lo};
  wire [1023:0]      slideAddressGen_slideMaskInput_lo_lo_lo = {slideAddressGen_slideMaskInput_lo_lo_lo_hi, slideAddressGen_slideMaskInput_lo_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_lo_hi_lo_lo_lo = {slideAddressGen_slideMaskInput_lo_lo_hi_lo_lo_lo_hi, slideAddressGen_slideMaskInput_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_lo_hi_lo_lo_hi = {slideAddressGen_slideMaskInput_lo_lo_hi_lo_lo_hi_hi, slideAddressGen_slideMaskInput_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_lo_lo_hi_lo_lo = {slideAddressGen_slideMaskInput_lo_lo_hi_lo_lo_hi, slideAddressGen_slideMaskInput_lo_lo_hi_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_lo_hi_lo_hi_lo = {slideAddressGen_slideMaskInput_lo_lo_hi_lo_hi_lo_hi, slideAddressGen_slideMaskInput_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_lo_hi_lo_hi_hi = {slideAddressGen_slideMaskInput_lo_lo_hi_lo_hi_hi_hi, slideAddressGen_slideMaskInput_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_lo_lo_hi_lo_hi = {slideAddressGen_slideMaskInput_lo_lo_hi_lo_hi_hi, slideAddressGen_slideMaskInput_lo_lo_hi_lo_hi_lo};
  wire [511:0]       slideAddressGen_slideMaskInput_lo_lo_hi_lo = {slideAddressGen_slideMaskInput_lo_lo_hi_lo_hi, slideAddressGen_slideMaskInput_lo_lo_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_lo_hi_hi_lo_lo = {slideAddressGen_slideMaskInput_lo_lo_hi_hi_lo_lo_hi, slideAddressGen_slideMaskInput_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_lo_hi_hi_lo_hi = {slideAddressGen_slideMaskInput_lo_lo_hi_hi_lo_hi_hi, slideAddressGen_slideMaskInput_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_lo_lo_hi_hi_lo = {slideAddressGen_slideMaskInput_lo_lo_hi_hi_lo_hi, slideAddressGen_slideMaskInput_lo_lo_hi_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_lo_hi_hi_hi_lo = {slideAddressGen_slideMaskInput_lo_lo_hi_hi_hi_lo_hi, slideAddressGen_slideMaskInput_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_lo_hi_hi_hi_hi = {slideAddressGen_slideMaskInput_lo_lo_hi_hi_hi_hi_hi, slideAddressGen_slideMaskInput_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_lo_lo_hi_hi_hi = {slideAddressGen_slideMaskInput_lo_lo_hi_hi_hi_hi, slideAddressGen_slideMaskInput_lo_lo_hi_hi_hi_lo};
  wire [511:0]       slideAddressGen_slideMaskInput_lo_lo_hi_hi = {slideAddressGen_slideMaskInput_lo_lo_hi_hi_hi, slideAddressGen_slideMaskInput_lo_lo_hi_hi_lo};
  wire [1023:0]      slideAddressGen_slideMaskInput_lo_lo_hi = {slideAddressGen_slideMaskInput_lo_lo_hi_hi, slideAddressGen_slideMaskInput_lo_lo_hi_lo};
  wire [2047:0]      slideAddressGen_slideMaskInput_lo_lo = {slideAddressGen_slideMaskInput_lo_lo_hi, slideAddressGen_slideMaskInput_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_hi_lo_lo_lo_lo = {slideAddressGen_slideMaskInput_lo_hi_lo_lo_lo_lo_hi, slideAddressGen_slideMaskInput_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_hi_lo_lo_lo_hi = {slideAddressGen_slideMaskInput_lo_hi_lo_lo_lo_hi_hi, slideAddressGen_slideMaskInput_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_lo_hi_lo_lo_lo = {slideAddressGen_slideMaskInput_lo_hi_lo_lo_lo_hi, slideAddressGen_slideMaskInput_lo_hi_lo_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_hi_lo_lo_hi_lo = {slideAddressGen_slideMaskInput_lo_hi_lo_lo_hi_lo_hi, slideAddressGen_slideMaskInput_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_hi_lo_lo_hi_hi = {slideAddressGen_slideMaskInput_lo_hi_lo_lo_hi_hi_hi, slideAddressGen_slideMaskInput_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_lo_hi_lo_lo_hi = {slideAddressGen_slideMaskInput_lo_hi_lo_lo_hi_hi, slideAddressGen_slideMaskInput_lo_hi_lo_lo_hi_lo};
  wire [511:0]       slideAddressGen_slideMaskInput_lo_hi_lo_lo = {slideAddressGen_slideMaskInput_lo_hi_lo_lo_hi, slideAddressGen_slideMaskInput_lo_hi_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_hi_lo_hi_lo_lo = {slideAddressGen_slideMaskInput_lo_hi_lo_hi_lo_lo_hi, slideAddressGen_slideMaskInput_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_hi_lo_hi_lo_hi = {slideAddressGen_slideMaskInput_lo_hi_lo_hi_lo_hi_hi, slideAddressGen_slideMaskInput_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_lo_hi_lo_hi_lo = {slideAddressGen_slideMaskInput_lo_hi_lo_hi_lo_hi, slideAddressGen_slideMaskInput_lo_hi_lo_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_hi_lo_hi_hi_lo = {slideAddressGen_slideMaskInput_lo_hi_lo_hi_hi_lo_hi, slideAddressGen_slideMaskInput_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_hi_lo_hi_hi_hi = {slideAddressGen_slideMaskInput_lo_hi_lo_hi_hi_hi_hi, slideAddressGen_slideMaskInput_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_lo_hi_lo_hi_hi = {slideAddressGen_slideMaskInput_lo_hi_lo_hi_hi_hi, slideAddressGen_slideMaskInput_lo_hi_lo_hi_hi_lo};
  wire [511:0]       slideAddressGen_slideMaskInput_lo_hi_lo_hi = {slideAddressGen_slideMaskInput_lo_hi_lo_hi_hi, slideAddressGen_slideMaskInput_lo_hi_lo_hi_lo};
  wire [1023:0]      slideAddressGen_slideMaskInput_lo_hi_lo = {slideAddressGen_slideMaskInput_lo_hi_lo_hi, slideAddressGen_slideMaskInput_lo_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_hi_hi_lo_lo_lo = {slideAddressGen_slideMaskInput_lo_hi_hi_lo_lo_lo_hi, slideAddressGen_slideMaskInput_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_hi_hi_lo_lo_hi = {slideAddressGen_slideMaskInput_lo_hi_hi_lo_lo_hi_hi, slideAddressGen_slideMaskInput_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_lo_hi_hi_lo_lo = {slideAddressGen_slideMaskInput_lo_hi_hi_lo_lo_hi, slideAddressGen_slideMaskInput_lo_hi_hi_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_hi_hi_lo_hi_lo = {slideAddressGen_slideMaskInput_lo_hi_hi_lo_hi_lo_hi, slideAddressGen_slideMaskInput_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_hi_hi_lo_hi_hi = {slideAddressGen_slideMaskInput_lo_hi_hi_lo_hi_hi_hi, slideAddressGen_slideMaskInput_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_lo_hi_hi_lo_hi = {slideAddressGen_slideMaskInput_lo_hi_hi_lo_hi_hi, slideAddressGen_slideMaskInput_lo_hi_hi_lo_hi_lo};
  wire [511:0]       slideAddressGen_slideMaskInput_lo_hi_hi_lo = {slideAddressGen_slideMaskInput_lo_hi_hi_lo_hi, slideAddressGen_slideMaskInput_lo_hi_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_hi_hi_hi_lo_lo = {slideAddressGen_slideMaskInput_lo_hi_hi_hi_lo_lo_hi, slideAddressGen_slideMaskInput_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_hi_hi_hi_lo_hi = {slideAddressGen_slideMaskInput_lo_hi_hi_hi_lo_hi_hi, slideAddressGen_slideMaskInput_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_lo_hi_hi_hi_lo = {slideAddressGen_slideMaskInput_lo_hi_hi_hi_lo_hi, slideAddressGen_slideMaskInput_lo_hi_hi_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_hi_hi_hi_hi_lo = {slideAddressGen_slideMaskInput_lo_hi_hi_hi_hi_lo_hi, slideAddressGen_slideMaskInput_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_hi_hi_hi_hi_hi = {slideAddressGen_slideMaskInput_lo_hi_hi_hi_hi_hi_hi, slideAddressGen_slideMaskInput_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_lo_hi_hi_hi_hi = {slideAddressGen_slideMaskInput_lo_hi_hi_hi_hi_hi, slideAddressGen_slideMaskInput_lo_hi_hi_hi_hi_lo};
  wire [511:0]       slideAddressGen_slideMaskInput_lo_hi_hi_hi = {slideAddressGen_slideMaskInput_lo_hi_hi_hi_hi, slideAddressGen_slideMaskInput_lo_hi_hi_hi_lo};
  wire [1023:0]      slideAddressGen_slideMaskInput_lo_hi_hi = {slideAddressGen_slideMaskInput_lo_hi_hi_hi, slideAddressGen_slideMaskInput_lo_hi_hi_lo};
  wire [2047:0]      slideAddressGen_slideMaskInput_lo_hi = {slideAddressGen_slideMaskInput_lo_hi_hi, slideAddressGen_slideMaskInput_lo_hi_lo};
  wire [4095:0]      slideAddressGen_slideMaskInput_lo = {slideAddressGen_slideMaskInput_lo_hi, slideAddressGen_slideMaskInput_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_lo_lo_lo_lo_lo = {slideAddressGen_slideMaskInput_hi_lo_lo_lo_lo_lo_hi, slideAddressGen_slideMaskInput_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_lo_lo_lo_lo_hi = {slideAddressGen_slideMaskInput_hi_lo_lo_lo_lo_hi_hi, slideAddressGen_slideMaskInput_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_hi_lo_lo_lo_lo = {slideAddressGen_slideMaskInput_hi_lo_lo_lo_lo_hi, slideAddressGen_slideMaskInput_hi_lo_lo_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_lo_lo_lo_hi_lo = {slideAddressGen_slideMaskInput_hi_lo_lo_lo_hi_lo_hi, slideAddressGen_slideMaskInput_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_lo_lo_lo_hi_hi = {slideAddressGen_slideMaskInput_hi_lo_lo_lo_hi_hi_hi, slideAddressGen_slideMaskInput_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_hi_lo_lo_lo_hi = {slideAddressGen_slideMaskInput_hi_lo_lo_lo_hi_hi, slideAddressGen_slideMaskInput_hi_lo_lo_lo_hi_lo};
  wire [511:0]       slideAddressGen_slideMaskInput_hi_lo_lo_lo = {slideAddressGen_slideMaskInput_hi_lo_lo_lo_hi, slideAddressGen_slideMaskInput_hi_lo_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_lo_lo_hi_lo_lo = {slideAddressGen_slideMaskInput_hi_lo_lo_hi_lo_lo_hi, slideAddressGen_slideMaskInput_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_lo_lo_hi_lo_hi = {slideAddressGen_slideMaskInput_hi_lo_lo_hi_lo_hi_hi, slideAddressGen_slideMaskInput_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_hi_lo_lo_hi_lo = {slideAddressGen_slideMaskInput_hi_lo_lo_hi_lo_hi, slideAddressGen_slideMaskInput_hi_lo_lo_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_lo_lo_hi_hi_lo = {slideAddressGen_slideMaskInput_hi_lo_lo_hi_hi_lo_hi, slideAddressGen_slideMaskInput_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_lo_lo_hi_hi_hi = {slideAddressGen_slideMaskInput_hi_lo_lo_hi_hi_hi_hi, slideAddressGen_slideMaskInput_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_hi_lo_lo_hi_hi = {slideAddressGen_slideMaskInput_hi_lo_lo_hi_hi_hi, slideAddressGen_slideMaskInput_hi_lo_lo_hi_hi_lo};
  wire [511:0]       slideAddressGen_slideMaskInput_hi_lo_lo_hi = {slideAddressGen_slideMaskInput_hi_lo_lo_hi_hi, slideAddressGen_slideMaskInput_hi_lo_lo_hi_lo};
  wire [1023:0]      slideAddressGen_slideMaskInput_hi_lo_lo = {slideAddressGen_slideMaskInput_hi_lo_lo_hi, slideAddressGen_slideMaskInput_hi_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_lo_hi_lo_lo_lo = {slideAddressGen_slideMaskInput_hi_lo_hi_lo_lo_lo_hi, slideAddressGen_slideMaskInput_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_lo_hi_lo_lo_hi = {slideAddressGen_slideMaskInput_hi_lo_hi_lo_lo_hi_hi, slideAddressGen_slideMaskInput_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_hi_lo_hi_lo_lo = {slideAddressGen_slideMaskInput_hi_lo_hi_lo_lo_hi, slideAddressGen_slideMaskInput_hi_lo_hi_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_lo_hi_lo_hi_lo = {slideAddressGen_slideMaskInput_hi_lo_hi_lo_hi_lo_hi, slideAddressGen_slideMaskInput_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_lo_hi_lo_hi_hi = {slideAddressGen_slideMaskInput_hi_lo_hi_lo_hi_hi_hi, slideAddressGen_slideMaskInput_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_hi_lo_hi_lo_hi = {slideAddressGen_slideMaskInput_hi_lo_hi_lo_hi_hi, slideAddressGen_slideMaskInput_hi_lo_hi_lo_hi_lo};
  wire [511:0]       slideAddressGen_slideMaskInput_hi_lo_hi_lo = {slideAddressGen_slideMaskInput_hi_lo_hi_lo_hi, slideAddressGen_slideMaskInput_hi_lo_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_lo_hi_hi_lo_lo = {slideAddressGen_slideMaskInput_hi_lo_hi_hi_lo_lo_hi, slideAddressGen_slideMaskInput_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_lo_hi_hi_lo_hi = {slideAddressGen_slideMaskInput_hi_lo_hi_hi_lo_hi_hi, slideAddressGen_slideMaskInput_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_hi_lo_hi_hi_lo = {slideAddressGen_slideMaskInput_hi_lo_hi_hi_lo_hi, slideAddressGen_slideMaskInput_hi_lo_hi_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_lo_hi_hi_hi_lo = {slideAddressGen_slideMaskInput_hi_lo_hi_hi_hi_lo_hi, slideAddressGen_slideMaskInput_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_lo_hi_hi_hi_hi = {slideAddressGen_slideMaskInput_hi_lo_hi_hi_hi_hi_hi, slideAddressGen_slideMaskInput_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_hi_lo_hi_hi_hi = {slideAddressGen_slideMaskInput_hi_lo_hi_hi_hi_hi, slideAddressGen_slideMaskInput_hi_lo_hi_hi_hi_lo};
  wire [511:0]       slideAddressGen_slideMaskInput_hi_lo_hi_hi = {slideAddressGen_slideMaskInput_hi_lo_hi_hi_hi, slideAddressGen_slideMaskInput_hi_lo_hi_hi_lo};
  wire [1023:0]      slideAddressGen_slideMaskInput_hi_lo_hi = {slideAddressGen_slideMaskInput_hi_lo_hi_hi, slideAddressGen_slideMaskInput_hi_lo_hi_lo};
  wire [2047:0]      slideAddressGen_slideMaskInput_hi_lo = {slideAddressGen_slideMaskInput_hi_lo_hi, slideAddressGen_slideMaskInput_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_hi_lo_lo_lo_lo = {slideAddressGen_slideMaskInput_hi_hi_lo_lo_lo_lo_hi, slideAddressGen_slideMaskInput_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_hi_lo_lo_lo_hi = {slideAddressGen_slideMaskInput_hi_hi_lo_lo_lo_hi_hi, slideAddressGen_slideMaskInput_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_hi_hi_lo_lo_lo = {slideAddressGen_slideMaskInput_hi_hi_lo_lo_lo_hi, slideAddressGen_slideMaskInput_hi_hi_lo_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_hi_lo_lo_hi_lo = {slideAddressGen_slideMaskInput_hi_hi_lo_lo_hi_lo_hi, slideAddressGen_slideMaskInput_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_hi_lo_lo_hi_hi = {slideAddressGen_slideMaskInput_hi_hi_lo_lo_hi_hi_hi, slideAddressGen_slideMaskInput_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_hi_hi_lo_lo_hi = {slideAddressGen_slideMaskInput_hi_hi_lo_lo_hi_hi, slideAddressGen_slideMaskInput_hi_hi_lo_lo_hi_lo};
  wire [511:0]       slideAddressGen_slideMaskInput_hi_hi_lo_lo = {slideAddressGen_slideMaskInput_hi_hi_lo_lo_hi, slideAddressGen_slideMaskInput_hi_hi_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_hi_lo_hi_lo_lo = {slideAddressGen_slideMaskInput_hi_hi_lo_hi_lo_lo_hi, slideAddressGen_slideMaskInput_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_hi_lo_hi_lo_hi = {slideAddressGen_slideMaskInput_hi_hi_lo_hi_lo_hi_hi, slideAddressGen_slideMaskInput_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_hi_hi_lo_hi_lo = {slideAddressGen_slideMaskInput_hi_hi_lo_hi_lo_hi, slideAddressGen_slideMaskInput_hi_hi_lo_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_hi_lo_hi_hi_lo = {slideAddressGen_slideMaskInput_hi_hi_lo_hi_hi_lo_hi, slideAddressGen_slideMaskInput_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_hi_lo_hi_hi_hi = {slideAddressGen_slideMaskInput_hi_hi_lo_hi_hi_hi_hi, slideAddressGen_slideMaskInput_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_hi_hi_lo_hi_hi = {slideAddressGen_slideMaskInput_hi_hi_lo_hi_hi_hi, slideAddressGen_slideMaskInput_hi_hi_lo_hi_hi_lo};
  wire [511:0]       slideAddressGen_slideMaskInput_hi_hi_lo_hi = {slideAddressGen_slideMaskInput_hi_hi_lo_hi_hi, slideAddressGen_slideMaskInput_hi_hi_lo_hi_lo};
  wire [1023:0]      slideAddressGen_slideMaskInput_hi_hi_lo = {slideAddressGen_slideMaskInput_hi_hi_lo_hi, slideAddressGen_slideMaskInput_hi_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_hi_hi_lo_lo_lo = {slideAddressGen_slideMaskInput_hi_hi_hi_lo_lo_lo_hi, slideAddressGen_slideMaskInput_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_hi_hi_lo_lo_hi = {slideAddressGen_slideMaskInput_hi_hi_hi_lo_lo_hi_hi, slideAddressGen_slideMaskInput_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_hi_hi_hi_lo_lo = {slideAddressGen_slideMaskInput_hi_hi_hi_lo_lo_hi, slideAddressGen_slideMaskInput_hi_hi_hi_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_hi_hi_lo_hi_lo = {slideAddressGen_slideMaskInput_hi_hi_hi_lo_hi_lo_hi, slideAddressGen_slideMaskInput_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_hi_hi_lo_hi_hi = {slideAddressGen_slideMaskInput_hi_hi_hi_lo_hi_hi_hi, slideAddressGen_slideMaskInput_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_hi_hi_hi_lo_hi = {slideAddressGen_slideMaskInput_hi_hi_hi_lo_hi_hi, slideAddressGen_slideMaskInput_hi_hi_hi_lo_hi_lo};
  wire [511:0]       slideAddressGen_slideMaskInput_hi_hi_hi_lo = {slideAddressGen_slideMaskInput_hi_hi_hi_lo_hi, slideAddressGen_slideMaskInput_hi_hi_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_hi_hi_hi_lo_lo = {slideAddressGen_slideMaskInput_hi_hi_hi_hi_lo_lo_hi, slideAddressGen_slideMaskInput_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_hi_hi_hi_lo_hi = {slideAddressGen_slideMaskInput_hi_hi_hi_hi_lo_hi_hi, slideAddressGen_slideMaskInput_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_hi_hi_hi_hi_lo = {slideAddressGen_slideMaskInput_hi_hi_hi_hi_lo_hi, slideAddressGen_slideMaskInput_hi_hi_hi_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_hi_hi_hi_hi_lo = {slideAddressGen_slideMaskInput_hi_hi_hi_hi_hi_lo_hi, slideAddressGen_slideMaskInput_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_hi_hi_hi_hi_hi = {slideAddressGen_slideMaskInput_hi_hi_hi_hi_hi_hi_hi, slideAddressGen_slideMaskInput_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_hi_hi_hi_hi_hi = {slideAddressGen_slideMaskInput_hi_hi_hi_hi_hi_hi, slideAddressGen_slideMaskInput_hi_hi_hi_hi_hi_lo};
  wire [511:0]       slideAddressGen_slideMaskInput_hi_hi_hi_hi = {slideAddressGen_slideMaskInput_hi_hi_hi_hi_hi, slideAddressGen_slideMaskInput_hi_hi_hi_hi_lo};
  wire [1023:0]      slideAddressGen_slideMaskInput_hi_hi_hi = {slideAddressGen_slideMaskInput_hi_hi_hi_hi, slideAddressGen_slideMaskInput_hi_hi_hi_lo};
  wire [2047:0]      slideAddressGen_slideMaskInput_hi_hi = {slideAddressGen_slideMaskInput_hi_hi_hi, slideAddressGen_slideMaskInput_hi_hi_lo};
  wire [4095:0]      slideAddressGen_slideMaskInput_hi = {slideAddressGen_slideMaskInput_hi_hi, slideAddressGen_slideMaskInput_hi_lo};
  wire [2047:0][3:0] _GEN_140 =
    {{slideAddressGen_slideMaskInput_hi[4095:4092]},
     {slideAddressGen_slideMaskInput_hi[4091:4088]},
     {slideAddressGen_slideMaskInput_hi[4087:4084]},
     {slideAddressGen_slideMaskInput_hi[4083:4080]},
     {slideAddressGen_slideMaskInput_hi[4079:4076]},
     {slideAddressGen_slideMaskInput_hi[4075:4072]},
     {slideAddressGen_slideMaskInput_hi[4071:4068]},
     {slideAddressGen_slideMaskInput_hi[4067:4064]},
     {slideAddressGen_slideMaskInput_hi[4063:4060]},
     {slideAddressGen_slideMaskInput_hi[4059:4056]},
     {slideAddressGen_slideMaskInput_hi[4055:4052]},
     {slideAddressGen_slideMaskInput_hi[4051:4048]},
     {slideAddressGen_slideMaskInput_hi[4047:4044]},
     {slideAddressGen_slideMaskInput_hi[4043:4040]},
     {slideAddressGen_slideMaskInput_hi[4039:4036]},
     {slideAddressGen_slideMaskInput_hi[4035:4032]},
     {slideAddressGen_slideMaskInput_hi[4031:4028]},
     {slideAddressGen_slideMaskInput_hi[4027:4024]},
     {slideAddressGen_slideMaskInput_hi[4023:4020]},
     {slideAddressGen_slideMaskInput_hi[4019:4016]},
     {slideAddressGen_slideMaskInput_hi[4015:4012]},
     {slideAddressGen_slideMaskInput_hi[4011:4008]},
     {slideAddressGen_slideMaskInput_hi[4007:4004]},
     {slideAddressGen_slideMaskInput_hi[4003:4000]},
     {slideAddressGen_slideMaskInput_hi[3999:3996]},
     {slideAddressGen_slideMaskInput_hi[3995:3992]},
     {slideAddressGen_slideMaskInput_hi[3991:3988]},
     {slideAddressGen_slideMaskInput_hi[3987:3984]},
     {slideAddressGen_slideMaskInput_hi[3983:3980]},
     {slideAddressGen_slideMaskInput_hi[3979:3976]},
     {slideAddressGen_slideMaskInput_hi[3975:3972]},
     {slideAddressGen_slideMaskInput_hi[3971:3968]},
     {slideAddressGen_slideMaskInput_hi[3967:3964]},
     {slideAddressGen_slideMaskInput_hi[3963:3960]},
     {slideAddressGen_slideMaskInput_hi[3959:3956]},
     {slideAddressGen_slideMaskInput_hi[3955:3952]},
     {slideAddressGen_slideMaskInput_hi[3951:3948]},
     {slideAddressGen_slideMaskInput_hi[3947:3944]},
     {slideAddressGen_slideMaskInput_hi[3943:3940]},
     {slideAddressGen_slideMaskInput_hi[3939:3936]},
     {slideAddressGen_slideMaskInput_hi[3935:3932]},
     {slideAddressGen_slideMaskInput_hi[3931:3928]},
     {slideAddressGen_slideMaskInput_hi[3927:3924]},
     {slideAddressGen_slideMaskInput_hi[3923:3920]},
     {slideAddressGen_slideMaskInput_hi[3919:3916]},
     {slideAddressGen_slideMaskInput_hi[3915:3912]},
     {slideAddressGen_slideMaskInput_hi[3911:3908]},
     {slideAddressGen_slideMaskInput_hi[3907:3904]},
     {slideAddressGen_slideMaskInput_hi[3903:3900]},
     {slideAddressGen_slideMaskInput_hi[3899:3896]},
     {slideAddressGen_slideMaskInput_hi[3895:3892]},
     {slideAddressGen_slideMaskInput_hi[3891:3888]},
     {slideAddressGen_slideMaskInput_hi[3887:3884]},
     {slideAddressGen_slideMaskInput_hi[3883:3880]},
     {slideAddressGen_slideMaskInput_hi[3879:3876]},
     {slideAddressGen_slideMaskInput_hi[3875:3872]},
     {slideAddressGen_slideMaskInput_hi[3871:3868]},
     {slideAddressGen_slideMaskInput_hi[3867:3864]},
     {slideAddressGen_slideMaskInput_hi[3863:3860]},
     {slideAddressGen_slideMaskInput_hi[3859:3856]},
     {slideAddressGen_slideMaskInput_hi[3855:3852]},
     {slideAddressGen_slideMaskInput_hi[3851:3848]},
     {slideAddressGen_slideMaskInput_hi[3847:3844]},
     {slideAddressGen_slideMaskInput_hi[3843:3840]},
     {slideAddressGen_slideMaskInput_hi[3839:3836]},
     {slideAddressGen_slideMaskInput_hi[3835:3832]},
     {slideAddressGen_slideMaskInput_hi[3831:3828]},
     {slideAddressGen_slideMaskInput_hi[3827:3824]},
     {slideAddressGen_slideMaskInput_hi[3823:3820]},
     {slideAddressGen_slideMaskInput_hi[3819:3816]},
     {slideAddressGen_slideMaskInput_hi[3815:3812]},
     {slideAddressGen_slideMaskInput_hi[3811:3808]},
     {slideAddressGen_slideMaskInput_hi[3807:3804]},
     {slideAddressGen_slideMaskInput_hi[3803:3800]},
     {slideAddressGen_slideMaskInput_hi[3799:3796]},
     {slideAddressGen_slideMaskInput_hi[3795:3792]},
     {slideAddressGen_slideMaskInput_hi[3791:3788]},
     {slideAddressGen_slideMaskInput_hi[3787:3784]},
     {slideAddressGen_slideMaskInput_hi[3783:3780]},
     {slideAddressGen_slideMaskInput_hi[3779:3776]},
     {slideAddressGen_slideMaskInput_hi[3775:3772]},
     {slideAddressGen_slideMaskInput_hi[3771:3768]},
     {slideAddressGen_slideMaskInput_hi[3767:3764]},
     {slideAddressGen_slideMaskInput_hi[3763:3760]},
     {slideAddressGen_slideMaskInput_hi[3759:3756]},
     {slideAddressGen_slideMaskInput_hi[3755:3752]},
     {slideAddressGen_slideMaskInput_hi[3751:3748]},
     {slideAddressGen_slideMaskInput_hi[3747:3744]},
     {slideAddressGen_slideMaskInput_hi[3743:3740]},
     {slideAddressGen_slideMaskInput_hi[3739:3736]},
     {slideAddressGen_slideMaskInput_hi[3735:3732]},
     {slideAddressGen_slideMaskInput_hi[3731:3728]},
     {slideAddressGen_slideMaskInput_hi[3727:3724]},
     {slideAddressGen_slideMaskInput_hi[3723:3720]},
     {slideAddressGen_slideMaskInput_hi[3719:3716]},
     {slideAddressGen_slideMaskInput_hi[3715:3712]},
     {slideAddressGen_slideMaskInput_hi[3711:3708]},
     {slideAddressGen_slideMaskInput_hi[3707:3704]},
     {slideAddressGen_slideMaskInput_hi[3703:3700]},
     {slideAddressGen_slideMaskInput_hi[3699:3696]},
     {slideAddressGen_slideMaskInput_hi[3695:3692]},
     {slideAddressGen_slideMaskInput_hi[3691:3688]},
     {slideAddressGen_slideMaskInput_hi[3687:3684]},
     {slideAddressGen_slideMaskInput_hi[3683:3680]},
     {slideAddressGen_slideMaskInput_hi[3679:3676]},
     {slideAddressGen_slideMaskInput_hi[3675:3672]},
     {slideAddressGen_slideMaskInput_hi[3671:3668]},
     {slideAddressGen_slideMaskInput_hi[3667:3664]},
     {slideAddressGen_slideMaskInput_hi[3663:3660]},
     {slideAddressGen_slideMaskInput_hi[3659:3656]},
     {slideAddressGen_slideMaskInput_hi[3655:3652]},
     {slideAddressGen_slideMaskInput_hi[3651:3648]},
     {slideAddressGen_slideMaskInput_hi[3647:3644]},
     {slideAddressGen_slideMaskInput_hi[3643:3640]},
     {slideAddressGen_slideMaskInput_hi[3639:3636]},
     {slideAddressGen_slideMaskInput_hi[3635:3632]},
     {slideAddressGen_slideMaskInput_hi[3631:3628]},
     {slideAddressGen_slideMaskInput_hi[3627:3624]},
     {slideAddressGen_slideMaskInput_hi[3623:3620]},
     {slideAddressGen_slideMaskInput_hi[3619:3616]},
     {slideAddressGen_slideMaskInput_hi[3615:3612]},
     {slideAddressGen_slideMaskInput_hi[3611:3608]},
     {slideAddressGen_slideMaskInput_hi[3607:3604]},
     {slideAddressGen_slideMaskInput_hi[3603:3600]},
     {slideAddressGen_slideMaskInput_hi[3599:3596]},
     {slideAddressGen_slideMaskInput_hi[3595:3592]},
     {slideAddressGen_slideMaskInput_hi[3591:3588]},
     {slideAddressGen_slideMaskInput_hi[3587:3584]},
     {slideAddressGen_slideMaskInput_hi[3583:3580]},
     {slideAddressGen_slideMaskInput_hi[3579:3576]},
     {slideAddressGen_slideMaskInput_hi[3575:3572]},
     {slideAddressGen_slideMaskInput_hi[3571:3568]},
     {slideAddressGen_slideMaskInput_hi[3567:3564]},
     {slideAddressGen_slideMaskInput_hi[3563:3560]},
     {slideAddressGen_slideMaskInput_hi[3559:3556]},
     {slideAddressGen_slideMaskInput_hi[3555:3552]},
     {slideAddressGen_slideMaskInput_hi[3551:3548]},
     {slideAddressGen_slideMaskInput_hi[3547:3544]},
     {slideAddressGen_slideMaskInput_hi[3543:3540]},
     {slideAddressGen_slideMaskInput_hi[3539:3536]},
     {slideAddressGen_slideMaskInput_hi[3535:3532]},
     {slideAddressGen_slideMaskInput_hi[3531:3528]},
     {slideAddressGen_slideMaskInput_hi[3527:3524]},
     {slideAddressGen_slideMaskInput_hi[3523:3520]},
     {slideAddressGen_slideMaskInput_hi[3519:3516]},
     {slideAddressGen_slideMaskInput_hi[3515:3512]},
     {slideAddressGen_slideMaskInput_hi[3511:3508]},
     {slideAddressGen_slideMaskInput_hi[3507:3504]},
     {slideAddressGen_slideMaskInput_hi[3503:3500]},
     {slideAddressGen_slideMaskInput_hi[3499:3496]},
     {slideAddressGen_slideMaskInput_hi[3495:3492]},
     {slideAddressGen_slideMaskInput_hi[3491:3488]},
     {slideAddressGen_slideMaskInput_hi[3487:3484]},
     {slideAddressGen_slideMaskInput_hi[3483:3480]},
     {slideAddressGen_slideMaskInput_hi[3479:3476]},
     {slideAddressGen_slideMaskInput_hi[3475:3472]},
     {slideAddressGen_slideMaskInput_hi[3471:3468]},
     {slideAddressGen_slideMaskInput_hi[3467:3464]},
     {slideAddressGen_slideMaskInput_hi[3463:3460]},
     {slideAddressGen_slideMaskInput_hi[3459:3456]},
     {slideAddressGen_slideMaskInput_hi[3455:3452]},
     {slideAddressGen_slideMaskInput_hi[3451:3448]},
     {slideAddressGen_slideMaskInput_hi[3447:3444]},
     {slideAddressGen_slideMaskInput_hi[3443:3440]},
     {slideAddressGen_slideMaskInput_hi[3439:3436]},
     {slideAddressGen_slideMaskInput_hi[3435:3432]},
     {slideAddressGen_slideMaskInput_hi[3431:3428]},
     {slideAddressGen_slideMaskInput_hi[3427:3424]},
     {slideAddressGen_slideMaskInput_hi[3423:3420]},
     {slideAddressGen_slideMaskInput_hi[3419:3416]},
     {slideAddressGen_slideMaskInput_hi[3415:3412]},
     {slideAddressGen_slideMaskInput_hi[3411:3408]},
     {slideAddressGen_slideMaskInput_hi[3407:3404]},
     {slideAddressGen_slideMaskInput_hi[3403:3400]},
     {slideAddressGen_slideMaskInput_hi[3399:3396]},
     {slideAddressGen_slideMaskInput_hi[3395:3392]},
     {slideAddressGen_slideMaskInput_hi[3391:3388]},
     {slideAddressGen_slideMaskInput_hi[3387:3384]},
     {slideAddressGen_slideMaskInput_hi[3383:3380]},
     {slideAddressGen_slideMaskInput_hi[3379:3376]},
     {slideAddressGen_slideMaskInput_hi[3375:3372]},
     {slideAddressGen_slideMaskInput_hi[3371:3368]},
     {slideAddressGen_slideMaskInput_hi[3367:3364]},
     {slideAddressGen_slideMaskInput_hi[3363:3360]},
     {slideAddressGen_slideMaskInput_hi[3359:3356]},
     {slideAddressGen_slideMaskInput_hi[3355:3352]},
     {slideAddressGen_slideMaskInput_hi[3351:3348]},
     {slideAddressGen_slideMaskInput_hi[3347:3344]},
     {slideAddressGen_slideMaskInput_hi[3343:3340]},
     {slideAddressGen_slideMaskInput_hi[3339:3336]},
     {slideAddressGen_slideMaskInput_hi[3335:3332]},
     {slideAddressGen_slideMaskInput_hi[3331:3328]},
     {slideAddressGen_slideMaskInput_hi[3327:3324]},
     {slideAddressGen_slideMaskInput_hi[3323:3320]},
     {slideAddressGen_slideMaskInput_hi[3319:3316]},
     {slideAddressGen_slideMaskInput_hi[3315:3312]},
     {slideAddressGen_slideMaskInput_hi[3311:3308]},
     {slideAddressGen_slideMaskInput_hi[3307:3304]},
     {slideAddressGen_slideMaskInput_hi[3303:3300]},
     {slideAddressGen_slideMaskInput_hi[3299:3296]},
     {slideAddressGen_slideMaskInput_hi[3295:3292]},
     {slideAddressGen_slideMaskInput_hi[3291:3288]},
     {slideAddressGen_slideMaskInput_hi[3287:3284]},
     {slideAddressGen_slideMaskInput_hi[3283:3280]},
     {slideAddressGen_slideMaskInput_hi[3279:3276]},
     {slideAddressGen_slideMaskInput_hi[3275:3272]},
     {slideAddressGen_slideMaskInput_hi[3271:3268]},
     {slideAddressGen_slideMaskInput_hi[3267:3264]},
     {slideAddressGen_slideMaskInput_hi[3263:3260]},
     {slideAddressGen_slideMaskInput_hi[3259:3256]},
     {slideAddressGen_slideMaskInput_hi[3255:3252]},
     {slideAddressGen_slideMaskInput_hi[3251:3248]},
     {slideAddressGen_slideMaskInput_hi[3247:3244]},
     {slideAddressGen_slideMaskInput_hi[3243:3240]},
     {slideAddressGen_slideMaskInput_hi[3239:3236]},
     {slideAddressGen_slideMaskInput_hi[3235:3232]},
     {slideAddressGen_slideMaskInput_hi[3231:3228]},
     {slideAddressGen_slideMaskInput_hi[3227:3224]},
     {slideAddressGen_slideMaskInput_hi[3223:3220]},
     {slideAddressGen_slideMaskInput_hi[3219:3216]},
     {slideAddressGen_slideMaskInput_hi[3215:3212]},
     {slideAddressGen_slideMaskInput_hi[3211:3208]},
     {slideAddressGen_slideMaskInput_hi[3207:3204]},
     {slideAddressGen_slideMaskInput_hi[3203:3200]},
     {slideAddressGen_slideMaskInput_hi[3199:3196]},
     {slideAddressGen_slideMaskInput_hi[3195:3192]},
     {slideAddressGen_slideMaskInput_hi[3191:3188]},
     {slideAddressGen_slideMaskInput_hi[3187:3184]},
     {slideAddressGen_slideMaskInput_hi[3183:3180]},
     {slideAddressGen_slideMaskInput_hi[3179:3176]},
     {slideAddressGen_slideMaskInput_hi[3175:3172]},
     {slideAddressGen_slideMaskInput_hi[3171:3168]},
     {slideAddressGen_slideMaskInput_hi[3167:3164]},
     {slideAddressGen_slideMaskInput_hi[3163:3160]},
     {slideAddressGen_slideMaskInput_hi[3159:3156]},
     {slideAddressGen_slideMaskInput_hi[3155:3152]},
     {slideAddressGen_slideMaskInput_hi[3151:3148]},
     {slideAddressGen_slideMaskInput_hi[3147:3144]},
     {slideAddressGen_slideMaskInput_hi[3143:3140]},
     {slideAddressGen_slideMaskInput_hi[3139:3136]},
     {slideAddressGen_slideMaskInput_hi[3135:3132]},
     {slideAddressGen_slideMaskInput_hi[3131:3128]},
     {slideAddressGen_slideMaskInput_hi[3127:3124]},
     {slideAddressGen_slideMaskInput_hi[3123:3120]},
     {slideAddressGen_slideMaskInput_hi[3119:3116]},
     {slideAddressGen_slideMaskInput_hi[3115:3112]},
     {slideAddressGen_slideMaskInput_hi[3111:3108]},
     {slideAddressGen_slideMaskInput_hi[3107:3104]},
     {slideAddressGen_slideMaskInput_hi[3103:3100]},
     {slideAddressGen_slideMaskInput_hi[3099:3096]},
     {slideAddressGen_slideMaskInput_hi[3095:3092]},
     {slideAddressGen_slideMaskInput_hi[3091:3088]},
     {slideAddressGen_slideMaskInput_hi[3087:3084]},
     {slideAddressGen_slideMaskInput_hi[3083:3080]},
     {slideAddressGen_slideMaskInput_hi[3079:3076]},
     {slideAddressGen_slideMaskInput_hi[3075:3072]},
     {slideAddressGen_slideMaskInput_hi[3071:3068]},
     {slideAddressGen_slideMaskInput_hi[3067:3064]},
     {slideAddressGen_slideMaskInput_hi[3063:3060]},
     {slideAddressGen_slideMaskInput_hi[3059:3056]},
     {slideAddressGen_slideMaskInput_hi[3055:3052]},
     {slideAddressGen_slideMaskInput_hi[3051:3048]},
     {slideAddressGen_slideMaskInput_hi[3047:3044]},
     {slideAddressGen_slideMaskInput_hi[3043:3040]},
     {slideAddressGen_slideMaskInput_hi[3039:3036]},
     {slideAddressGen_slideMaskInput_hi[3035:3032]},
     {slideAddressGen_slideMaskInput_hi[3031:3028]},
     {slideAddressGen_slideMaskInput_hi[3027:3024]},
     {slideAddressGen_slideMaskInput_hi[3023:3020]},
     {slideAddressGen_slideMaskInput_hi[3019:3016]},
     {slideAddressGen_slideMaskInput_hi[3015:3012]},
     {slideAddressGen_slideMaskInput_hi[3011:3008]},
     {slideAddressGen_slideMaskInput_hi[3007:3004]},
     {slideAddressGen_slideMaskInput_hi[3003:3000]},
     {slideAddressGen_slideMaskInput_hi[2999:2996]},
     {slideAddressGen_slideMaskInput_hi[2995:2992]},
     {slideAddressGen_slideMaskInput_hi[2991:2988]},
     {slideAddressGen_slideMaskInput_hi[2987:2984]},
     {slideAddressGen_slideMaskInput_hi[2983:2980]},
     {slideAddressGen_slideMaskInput_hi[2979:2976]},
     {slideAddressGen_slideMaskInput_hi[2975:2972]},
     {slideAddressGen_slideMaskInput_hi[2971:2968]},
     {slideAddressGen_slideMaskInput_hi[2967:2964]},
     {slideAddressGen_slideMaskInput_hi[2963:2960]},
     {slideAddressGen_slideMaskInput_hi[2959:2956]},
     {slideAddressGen_slideMaskInput_hi[2955:2952]},
     {slideAddressGen_slideMaskInput_hi[2951:2948]},
     {slideAddressGen_slideMaskInput_hi[2947:2944]},
     {slideAddressGen_slideMaskInput_hi[2943:2940]},
     {slideAddressGen_slideMaskInput_hi[2939:2936]},
     {slideAddressGen_slideMaskInput_hi[2935:2932]},
     {slideAddressGen_slideMaskInput_hi[2931:2928]},
     {slideAddressGen_slideMaskInput_hi[2927:2924]},
     {slideAddressGen_slideMaskInput_hi[2923:2920]},
     {slideAddressGen_slideMaskInput_hi[2919:2916]},
     {slideAddressGen_slideMaskInput_hi[2915:2912]},
     {slideAddressGen_slideMaskInput_hi[2911:2908]},
     {slideAddressGen_slideMaskInput_hi[2907:2904]},
     {slideAddressGen_slideMaskInput_hi[2903:2900]},
     {slideAddressGen_slideMaskInput_hi[2899:2896]},
     {slideAddressGen_slideMaskInput_hi[2895:2892]},
     {slideAddressGen_slideMaskInput_hi[2891:2888]},
     {slideAddressGen_slideMaskInput_hi[2887:2884]},
     {slideAddressGen_slideMaskInput_hi[2883:2880]},
     {slideAddressGen_slideMaskInput_hi[2879:2876]},
     {slideAddressGen_slideMaskInput_hi[2875:2872]},
     {slideAddressGen_slideMaskInput_hi[2871:2868]},
     {slideAddressGen_slideMaskInput_hi[2867:2864]},
     {slideAddressGen_slideMaskInput_hi[2863:2860]},
     {slideAddressGen_slideMaskInput_hi[2859:2856]},
     {slideAddressGen_slideMaskInput_hi[2855:2852]},
     {slideAddressGen_slideMaskInput_hi[2851:2848]},
     {slideAddressGen_slideMaskInput_hi[2847:2844]},
     {slideAddressGen_slideMaskInput_hi[2843:2840]},
     {slideAddressGen_slideMaskInput_hi[2839:2836]},
     {slideAddressGen_slideMaskInput_hi[2835:2832]},
     {slideAddressGen_slideMaskInput_hi[2831:2828]},
     {slideAddressGen_slideMaskInput_hi[2827:2824]},
     {slideAddressGen_slideMaskInput_hi[2823:2820]},
     {slideAddressGen_slideMaskInput_hi[2819:2816]},
     {slideAddressGen_slideMaskInput_hi[2815:2812]},
     {slideAddressGen_slideMaskInput_hi[2811:2808]},
     {slideAddressGen_slideMaskInput_hi[2807:2804]},
     {slideAddressGen_slideMaskInput_hi[2803:2800]},
     {slideAddressGen_slideMaskInput_hi[2799:2796]},
     {slideAddressGen_slideMaskInput_hi[2795:2792]},
     {slideAddressGen_slideMaskInput_hi[2791:2788]},
     {slideAddressGen_slideMaskInput_hi[2787:2784]},
     {slideAddressGen_slideMaskInput_hi[2783:2780]},
     {slideAddressGen_slideMaskInput_hi[2779:2776]},
     {slideAddressGen_slideMaskInput_hi[2775:2772]},
     {slideAddressGen_slideMaskInput_hi[2771:2768]},
     {slideAddressGen_slideMaskInput_hi[2767:2764]},
     {slideAddressGen_slideMaskInput_hi[2763:2760]},
     {slideAddressGen_slideMaskInput_hi[2759:2756]},
     {slideAddressGen_slideMaskInput_hi[2755:2752]},
     {slideAddressGen_slideMaskInput_hi[2751:2748]},
     {slideAddressGen_slideMaskInput_hi[2747:2744]},
     {slideAddressGen_slideMaskInput_hi[2743:2740]},
     {slideAddressGen_slideMaskInput_hi[2739:2736]},
     {slideAddressGen_slideMaskInput_hi[2735:2732]},
     {slideAddressGen_slideMaskInput_hi[2731:2728]},
     {slideAddressGen_slideMaskInput_hi[2727:2724]},
     {slideAddressGen_slideMaskInput_hi[2723:2720]},
     {slideAddressGen_slideMaskInput_hi[2719:2716]},
     {slideAddressGen_slideMaskInput_hi[2715:2712]},
     {slideAddressGen_slideMaskInput_hi[2711:2708]},
     {slideAddressGen_slideMaskInput_hi[2707:2704]},
     {slideAddressGen_slideMaskInput_hi[2703:2700]},
     {slideAddressGen_slideMaskInput_hi[2699:2696]},
     {slideAddressGen_slideMaskInput_hi[2695:2692]},
     {slideAddressGen_slideMaskInput_hi[2691:2688]},
     {slideAddressGen_slideMaskInput_hi[2687:2684]},
     {slideAddressGen_slideMaskInput_hi[2683:2680]},
     {slideAddressGen_slideMaskInput_hi[2679:2676]},
     {slideAddressGen_slideMaskInput_hi[2675:2672]},
     {slideAddressGen_slideMaskInput_hi[2671:2668]},
     {slideAddressGen_slideMaskInput_hi[2667:2664]},
     {slideAddressGen_slideMaskInput_hi[2663:2660]},
     {slideAddressGen_slideMaskInput_hi[2659:2656]},
     {slideAddressGen_slideMaskInput_hi[2655:2652]},
     {slideAddressGen_slideMaskInput_hi[2651:2648]},
     {slideAddressGen_slideMaskInput_hi[2647:2644]},
     {slideAddressGen_slideMaskInput_hi[2643:2640]},
     {slideAddressGen_slideMaskInput_hi[2639:2636]},
     {slideAddressGen_slideMaskInput_hi[2635:2632]},
     {slideAddressGen_slideMaskInput_hi[2631:2628]},
     {slideAddressGen_slideMaskInput_hi[2627:2624]},
     {slideAddressGen_slideMaskInput_hi[2623:2620]},
     {slideAddressGen_slideMaskInput_hi[2619:2616]},
     {slideAddressGen_slideMaskInput_hi[2615:2612]},
     {slideAddressGen_slideMaskInput_hi[2611:2608]},
     {slideAddressGen_slideMaskInput_hi[2607:2604]},
     {slideAddressGen_slideMaskInput_hi[2603:2600]},
     {slideAddressGen_slideMaskInput_hi[2599:2596]},
     {slideAddressGen_slideMaskInput_hi[2595:2592]},
     {slideAddressGen_slideMaskInput_hi[2591:2588]},
     {slideAddressGen_slideMaskInput_hi[2587:2584]},
     {slideAddressGen_slideMaskInput_hi[2583:2580]},
     {slideAddressGen_slideMaskInput_hi[2579:2576]},
     {slideAddressGen_slideMaskInput_hi[2575:2572]},
     {slideAddressGen_slideMaskInput_hi[2571:2568]},
     {slideAddressGen_slideMaskInput_hi[2567:2564]},
     {slideAddressGen_slideMaskInput_hi[2563:2560]},
     {slideAddressGen_slideMaskInput_hi[2559:2556]},
     {slideAddressGen_slideMaskInput_hi[2555:2552]},
     {slideAddressGen_slideMaskInput_hi[2551:2548]},
     {slideAddressGen_slideMaskInput_hi[2547:2544]},
     {slideAddressGen_slideMaskInput_hi[2543:2540]},
     {slideAddressGen_slideMaskInput_hi[2539:2536]},
     {slideAddressGen_slideMaskInput_hi[2535:2532]},
     {slideAddressGen_slideMaskInput_hi[2531:2528]},
     {slideAddressGen_slideMaskInput_hi[2527:2524]},
     {slideAddressGen_slideMaskInput_hi[2523:2520]},
     {slideAddressGen_slideMaskInput_hi[2519:2516]},
     {slideAddressGen_slideMaskInput_hi[2515:2512]},
     {slideAddressGen_slideMaskInput_hi[2511:2508]},
     {slideAddressGen_slideMaskInput_hi[2507:2504]},
     {slideAddressGen_slideMaskInput_hi[2503:2500]},
     {slideAddressGen_slideMaskInput_hi[2499:2496]},
     {slideAddressGen_slideMaskInput_hi[2495:2492]},
     {slideAddressGen_slideMaskInput_hi[2491:2488]},
     {slideAddressGen_slideMaskInput_hi[2487:2484]},
     {slideAddressGen_slideMaskInput_hi[2483:2480]},
     {slideAddressGen_slideMaskInput_hi[2479:2476]},
     {slideAddressGen_slideMaskInput_hi[2475:2472]},
     {slideAddressGen_slideMaskInput_hi[2471:2468]},
     {slideAddressGen_slideMaskInput_hi[2467:2464]},
     {slideAddressGen_slideMaskInput_hi[2463:2460]},
     {slideAddressGen_slideMaskInput_hi[2459:2456]},
     {slideAddressGen_slideMaskInput_hi[2455:2452]},
     {slideAddressGen_slideMaskInput_hi[2451:2448]},
     {slideAddressGen_slideMaskInput_hi[2447:2444]},
     {slideAddressGen_slideMaskInput_hi[2443:2440]},
     {slideAddressGen_slideMaskInput_hi[2439:2436]},
     {slideAddressGen_slideMaskInput_hi[2435:2432]},
     {slideAddressGen_slideMaskInput_hi[2431:2428]},
     {slideAddressGen_slideMaskInput_hi[2427:2424]},
     {slideAddressGen_slideMaskInput_hi[2423:2420]},
     {slideAddressGen_slideMaskInput_hi[2419:2416]},
     {slideAddressGen_slideMaskInput_hi[2415:2412]},
     {slideAddressGen_slideMaskInput_hi[2411:2408]},
     {slideAddressGen_slideMaskInput_hi[2407:2404]},
     {slideAddressGen_slideMaskInput_hi[2403:2400]},
     {slideAddressGen_slideMaskInput_hi[2399:2396]},
     {slideAddressGen_slideMaskInput_hi[2395:2392]},
     {slideAddressGen_slideMaskInput_hi[2391:2388]},
     {slideAddressGen_slideMaskInput_hi[2387:2384]},
     {slideAddressGen_slideMaskInput_hi[2383:2380]},
     {slideAddressGen_slideMaskInput_hi[2379:2376]},
     {slideAddressGen_slideMaskInput_hi[2375:2372]},
     {slideAddressGen_slideMaskInput_hi[2371:2368]},
     {slideAddressGen_slideMaskInput_hi[2367:2364]},
     {slideAddressGen_slideMaskInput_hi[2363:2360]},
     {slideAddressGen_slideMaskInput_hi[2359:2356]},
     {slideAddressGen_slideMaskInput_hi[2355:2352]},
     {slideAddressGen_slideMaskInput_hi[2351:2348]},
     {slideAddressGen_slideMaskInput_hi[2347:2344]},
     {slideAddressGen_slideMaskInput_hi[2343:2340]},
     {slideAddressGen_slideMaskInput_hi[2339:2336]},
     {slideAddressGen_slideMaskInput_hi[2335:2332]},
     {slideAddressGen_slideMaskInput_hi[2331:2328]},
     {slideAddressGen_slideMaskInput_hi[2327:2324]},
     {slideAddressGen_slideMaskInput_hi[2323:2320]},
     {slideAddressGen_slideMaskInput_hi[2319:2316]},
     {slideAddressGen_slideMaskInput_hi[2315:2312]},
     {slideAddressGen_slideMaskInput_hi[2311:2308]},
     {slideAddressGen_slideMaskInput_hi[2307:2304]},
     {slideAddressGen_slideMaskInput_hi[2303:2300]},
     {slideAddressGen_slideMaskInput_hi[2299:2296]},
     {slideAddressGen_slideMaskInput_hi[2295:2292]},
     {slideAddressGen_slideMaskInput_hi[2291:2288]},
     {slideAddressGen_slideMaskInput_hi[2287:2284]},
     {slideAddressGen_slideMaskInput_hi[2283:2280]},
     {slideAddressGen_slideMaskInput_hi[2279:2276]},
     {slideAddressGen_slideMaskInput_hi[2275:2272]},
     {slideAddressGen_slideMaskInput_hi[2271:2268]},
     {slideAddressGen_slideMaskInput_hi[2267:2264]},
     {slideAddressGen_slideMaskInput_hi[2263:2260]},
     {slideAddressGen_slideMaskInput_hi[2259:2256]},
     {slideAddressGen_slideMaskInput_hi[2255:2252]},
     {slideAddressGen_slideMaskInput_hi[2251:2248]},
     {slideAddressGen_slideMaskInput_hi[2247:2244]},
     {slideAddressGen_slideMaskInput_hi[2243:2240]},
     {slideAddressGen_slideMaskInput_hi[2239:2236]},
     {slideAddressGen_slideMaskInput_hi[2235:2232]},
     {slideAddressGen_slideMaskInput_hi[2231:2228]},
     {slideAddressGen_slideMaskInput_hi[2227:2224]},
     {slideAddressGen_slideMaskInput_hi[2223:2220]},
     {slideAddressGen_slideMaskInput_hi[2219:2216]},
     {slideAddressGen_slideMaskInput_hi[2215:2212]},
     {slideAddressGen_slideMaskInput_hi[2211:2208]},
     {slideAddressGen_slideMaskInput_hi[2207:2204]},
     {slideAddressGen_slideMaskInput_hi[2203:2200]},
     {slideAddressGen_slideMaskInput_hi[2199:2196]},
     {slideAddressGen_slideMaskInput_hi[2195:2192]},
     {slideAddressGen_slideMaskInput_hi[2191:2188]},
     {slideAddressGen_slideMaskInput_hi[2187:2184]},
     {slideAddressGen_slideMaskInput_hi[2183:2180]},
     {slideAddressGen_slideMaskInput_hi[2179:2176]},
     {slideAddressGen_slideMaskInput_hi[2175:2172]},
     {slideAddressGen_slideMaskInput_hi[2171:2168]},
     {slideAddressGen_slideMaskInput_hi[2167:2164]},
     {slideAddressGen_slideMaskInput_hi[2163:2160]},
     {slideAddressGen_slideMaskInput_hi[2159:2156]},
     {slideAddressGen_slideMaskInput_hi[2155:2152]},
     {slideAddressGen_slideMaskInput_hi[2151:2148]},
     {slideAddressGen_slideMaskInput_hi[2147:2144]},
     {slideAddressGen_slideMaskInput_hi[2143:2140]},
     {slideAddressGen_slideMaskInput_hi[2139:2136]},
     {slideAddressGen_slideMaskInput_hi[2135:2132]},
     {slideAddressGen_slideMaskInput_hi[2131:2128]},
     {slideAddressGen_slideMaskInput_hi[2127:2124]},
     {slideAddressGen_slideMaskInput_hi[2123:2120]},
     {slideAddressGen_slideMaskInput_hi[2119:2116]},
     {slideAddressGen_slideMaskInput_hi[2115:2112]},
     {slideAddressGen_slideMaskInput_hi[2111:2108]},
     {slideAddressGen_slideMaskInput_hi[2107:2104]},
     {slideAddressGen_slideMaskInput_hi[2103:2100]},
     {slideAddressGen_slideMaskInput_hi[2099:2096]},
     {slideAddressGen_slideMaskInput_hi[2095:2092]},
     {slideAddressGen_slideMaskInput_hi[2091:2088]},
     {slideAddressGen_slideMaskInput_hi[2087:2084]},
     {slideAddressGen_slideMaskInput_hi[2083:2080]},
     {slideAddressGen_slideMaskInput_hi[2079:2076]},
     {slideAddressGen_slideMaskInput_hi[2075:2072]},
     {slideAddressGen_slideMaskInput_hi[2071:2068]},
     {slideAddressGen_slideMaskInput_hi[2067:2064]},
     {slideAddressGen_slideMaskInput_hi[2063:2060]},
     {slideAddressGen_slideMaskInput_hi[2059:2056]},
     {slideAddressGen_slideMaskInput_hi[2055:2052]},
     {slideAddressGen_slideMaskInput_hi[2051:2048]},
     {slideAddressGen_slideMaskInput_hi[2047:2044]},
     {slideAddressGen_slideMaskInput_hi[2043:2040]},
     {slideAddressGen_slideMaskInput_hi[2039:2036]},
     {slideAddressGen_slideMaskInput_hi[2035:2032]},
     {slideAddressGen_slideMaskInput_hi[2031:2028]},
     {slideAddressGen_slideMaskInput_hi[2027:2024]},
     {slideAddressGen_slideMaskInput_hi[2023:2020]},
     {slideAddressGen_slideMaskInput_hi[2019:2016]},
     {slideAddressGen_slideMaskInput_hi[2015:2012]},
     {slideAddressGen_slideMaskInput_hi[2011:2008]},
     {slideAddressGen_slideMaskInput_hi[2007:2004]},
     {slideAddressGen_slideMaskInput_hi[2003:2000]},
     {slideAddressGen_slideMaskInput_hi[1999:1996]},
     {slideAddressGen_slideMaskInput_hi[1995:1992]},
     {slideAddressGen_slideMaskInput_hi[1991:1988]},
     {slideAddressGen_slideMaskInput_hi[1987:1984]},
     {slideAddressGen_slideMaskInput_hi[1983:1980]},
     {slideAddressGen_slideMaskInput_hi[1979:1976]},
     {slideAddressGen_slideMaskInput_hi[1975:1972]},
     {slideAddressGen_slideMaskInput_hi[1971:1968]},
     {slideAddressGen_slideMaskInput_hi[1967:1964]},
     {slideAddressGen_slideMaskInput_hi[1963:1960]},
     {slideAddressGen_slideMaskInput_hi[1959:1956]},
     {slideAddressGen_slideMaskInput_hi[1955:1952]},
     {slideAddressGen_slideMaskInput_hi[1951:1948]},
     {slideAddressGen_slideMaskInput_hi[1947:1944]},
     {slideAddressGen_slideMaskInput_hi[1943:1940]},
     {slideAddressGen_slideMaskInput_hi[1939:1936]},
     {slideAddressGen_slideMaskInput_hi[1935:1932]},
     {slideAddressGen_slideMaskInput_hi[1931:1928]},
     {slideAddressGen_slideMaskInput_hi[1927:1924]},
     {slideAddressGen_slideMaskInput_hi[1923:1920]},
     {slideAddressGen_slideMaskInput_hi[1919:1916]},
     {slideAddressGen_slideMaskInput_hi[1915:1912]},
     {slideAddressGen_slideMaskInput_hi[1911:1908]},
     {slideAddressGen_slideMaskInput_hi[1907:1904]},
     {slideAddressGen_slideMaskInput_hi[1903:1900]},
     {slideAddressGen_slideMaskInput_hi[1899:1896]},
     {slideAddressGen_slideMaskInput_hi[1895:1892]},
     {slideAddressGen_slideMaskInput_hi[1891:1888]},
     {slideAddressGen_slideMaskInput_hi[1887:1884]},
     {slideAddressGen_slideMaskInput_hi[1883:1880]},
     {slideAddressGen_slideMaskInput_hi[1879:1876]},
     {slideAddressGen_slideMaskInput_hi[1875:1872]},
     {slideAddressGen_slideMaskInput_hi[1871:1868]},
     {slideAddressGen_slideMaskInput_hi[1867:1864]},
     {slideAddressGen_slideMaskInput_hi[1863:1860]},
     {slideAddressGen_slideMaskInput_hi[1859:1856]},
     {slideAddressGen_slideMaskInput_hi[1855:1852]},
     {slideAddressGen_slideMaskInput_hi[1851:1848]},
     {slideAddressGen_slideMaskInput_hi[1847:1844]},
     {slideAddressGen_slideMaskInput_hi[1843:1840]},
     {slideAddressGen_slideMaskInput_hi[1839:1836]},
     {slideAddressGen_slideMaskInput_hi[1835:1832]},
     {slideAddressGen_slideMaskInput_hi[1831:1828]},
     {slideAddressGen_slideMaskInput_hi[1827:1824]},
     {slideAddressGen_slideMaskInput_hi[1823:1820]},
     {slideAddressGen_slideMaskInput_hi[1819:1816]},
     {slideAddressGen_slideMaskInput_hi[1815:1812]},
     {slideAddressGen_slideMaskInput_hi[1811:1808]},
     {slideAddressGen_slideMaskInput_hi[1807:1804]},
     {slideAddressGen_slideMaskInput_hi[1803:1800]},
     {slideAddressGen_slideMaskInput_hi[1799:1796]},
     {slideAddressGen_slideMaskInput_hi[1795:1792]},
     {slideAddressGen_slideMaskInput_hi[1791:1788]},
     {slideAddressGen_slideMaskInput_hi[1787:1784]},
     {slideAddressGen_slideMaskInput_hi[1783:1780]},
     {slideAddressGen_slideMaskInput_hi[1779:1776]},
     {slideAddressGen_slideMaskInput_hi[1775:1772]},
     {slideAddressGen_slideMaskInput_hi[1771:1768]},
     {slideAddressGen_slideMaskInput_hi[1767:1764]},
     {slideAddressGen_slideMaskInput_hi[1763:1760]},
     {slideAddressGen_slideMaskInput_hi[1759:1756]},
     {slideAddressGen_slideMaskInput_hi[1755:1752]},
     {slideAddressGen_slideMaskInput_hi[1751:1748]},
     {slideAddressGen_slideMaskInput_hi[1747:1744]},
     {slideAddressGen_slideMaskInput_hi[1743:1740]},
     {slideAddressGen_slideMaskInput_hi[1739:1736]},
     {slideAddressGen_slideMaskInput_hi[1735:1732]},
     {slideAddressGen_slideMaskInput_hi[1731:1728]},
     {slideAddressGen_slideMaskInput_hi[1727:1724]},
     {slideAddressGen_slideMaskInput_hi[1723:1720]},
     {slideAddressGen_slideMaskInput_hi[1719:1716]},
     {slideAddressGen_slideMaskInput_hi[1715:1712]},
     {slideAddressGen_slideMaskInput_hi[1711:1708]},
     {slideAddressGen_slideMaskInput_hi[1707:1704]},
     {slideAddressGen_slideMaskInput_hi[1703:1700]},
     {slideAddressGen_slideMaskInput_hi[1699:1696]},
     {slideAddressGen_slideMaskInput_hi[1695:1692]},
     {slideAddressGen_slideMaskInput_hi[1691:1688]},
     {slideAddressGen_slideMaskInput_hi[1687:1684]},
     {slideAddressGen_slideMaskInput_hi[1683:1680]},
     {slideAddressGen_slideMaskInput_hi[1679:1676]},
     {slideAddressGen_slideMaskInput_hi[1675:1672]},
     {slideAddressGen_slideMaskInput_hi[1671:1668]},
     {slideAddressGen_slideMaskInput_hi[1667:1664]},
     {slideAddressGen_slideMaskInput_hi[1663:1660]},
     {slideAddressGen_slideMaskInput_hi[1659:1656]},
     {slideAddressGen_slideMaskInput_hi[1655:1652]},
     {slideAddressGen_slideMaskInput_hi[1651:1648]},
     {slideAddressGen_slideMaskInput_hi[1647:1644]},
     {slideAddressGen_slideMaskInput_hi[1643:1640]},
     {slideAddressGen_slideMaskInput_hi[1639:1636]},
     {slideAddressGen_slideMaskInput_hi[1635:1632]},
     {slideAddressGen_slideMaskInput_hi[1631:1628]},
     {slideAddressGen_slideMaskInput_hi[1627:1624]},
     {slideAddressGen_slideMaskInput_hi[1623:1620]},
     {slideAddressGen_slideMaskInput_hi[1619:1616]},
     {slideAddressGen_slideMaskInput_hi[1615:1612]},
     {slideAddressGen_slideMaskInput_hi[1611:1608]},
     {slideAddressGen_slideMaskInput_hi[1607:1604]},
     {slideAddressGen_slideMaskInput_hi[1603:1600]},
     {slideAddressGen_slideMaskInput_hi[1599:1596]},
     {slideAddressGen_slideMaskInput_hi[1595:1592]},
     {slideAddressGen_slideMaskInput_hi[1591:1588]},
     {slideAddressGen_slideMaskInput_hi[1587:1584]},
     {slideAddressGen_slideMaskInput_hi[1583:1580]},
     {slideAddressGen_slideMaskInput_hi[1579:1576]},
     {slideAddressGen_slideMaskInput_hi[1575:1572]},
     {slideAddressGen_slideMaskInput_hi[1571:1568]},
     {slideAddressGen_slideMaskInput_hi[1567:1564]},
     {slideAddressGen_slideMaskInput_hi[1563:1560]},
     {slideAddressGen_slideMaskInput_hi[1559:1556]},
     {slideAddressGen_slideMaskInput_hi[1555:1552]},
     {slideAddressGen_slideMaskInput_hi[1551:1548]},
     {slideAddressGen_slideMaskInput_hi[1547:1544]},
     {slideAddressGen_slideMaskInput_hi[1543:1540]},
     {slideAddressGen_slideMaskInput_hi[1539:1536]},
     {slideAddressGen_slideMaskInput_hi[1535:1532]},
     {slideAddressGen_slideMaskInput_hi[1531:1528]},
     {slideAddressGen_slideMaskInput_hi[1527:1524]},
     {slideAddressGen_slideMaskInput_hi[1523:1520]},
     {slideAddressGen_slideMaskInput_hi[1519:1516]},
     {slideAddressGen_slideMaskInput_hi[1515:1512]},
     {slideAddressGen_slideMaskInput_hi[1511:1508]},
     {slideAddressGen_slideMaskInput_hi[1507:1504]},
     {slideAddressGen_slideMaskInput_hi[1503:1500]},
     {slideAddressGen_slideMaskInput_hi[1499:1496]},
     {slideAddressGen_slideMaskInput_hi[1495:1492]},
     {slideAddressGen_slideMaskInput_hi[1491:1488]},
     {slideAddressGen_slideMaskInput_hi[1487:1484]},
     {slideAddressGen_slideMaskInput_hi[1483:1480]},
     {slideAddressGen_slideMaskInput_hi[1479:1476]},
     {slideAddressGen_slideMaskInput_hi[1475:1472]},
     {slideAddressGen_slideMaskInput_hi[1471:1468]},
     {slideAddressGen_slideMaskInput_hi[1467:1464]},
     {slideAddressGen_slideMaskInput_hi[1463:1460]},
     {slideAddressGen_slideMaskInput_hi[1459:1456]},
     {slideAddressGen_slideMaskInput_hi[1455:1452]},
     {slideAddressGen_slideMaskInput_hi[1451:1448]},
     {slideAddressGen_slideMaskInput_hi[1447:1444]},
     {slideAddressGen_slideMaskInput_hi[1443:1440]},
     {slideAddressGen_slideMaskInput_hi[1439:1436]},
     {slideAddressGen_slideMaskInput_hi[1435:1432]},
     {slideAddressGen_slideMaskInput_hi[1431:1428]},
     {slideAddressGen_slideMaskInput_hi[1427:1424]},
     {slideAddressGen_slideMaskInput_hi[1423:1420]},
     {slideAddressGen_slideMaskInput_hi[1419:1416]},
     {slideAddressGen_slideMaskInput_hi[1415:1412]},
     {slideAddressGen_slideMaskInput_hi[1411:1408]},
     {slideAddressGen_slideMaskInput_hi[1407:1404]},
     {slideAddressGen_slideMaskInput_hi[1403:1400]},
     {slideAddressGen_slideMaskInput_hi[1399:1396]},
     {slideAddressGen_slideMaskInput_hi[1395:1392]},
     {slideAddressGen_slideMaskInput_hi[1391:1388]},
     {slideAddressGen_slideMaskInput_hi[1387:1384]},
     {slideAddressGen_slideMaskInput_hi[1383:1380]},
     {slideAddressGen_slideMaskInput_hi[1379:1376]},
     {slideAddressGen_slideMaskInput_hi[1375:1372]},
     {slideAddressGen_slideMaskInput_hi[1371:1368]},
     {slideAddressGen_slideMaskInput_hi[1367:1364]},
     {slideAddressGen_slideMaskInput_hi[1363:1360]},
     {slideAddressGen_slideMaskInput_hi[1359:1356]},
     {slideAddressGen_slideMaskInput_hi[1355:1352]},
     {slideAddressGen_slideMaskInput_hi[1351:1348]},
     {slideAddressGen_slideMaskInput_hi[1347:1344]},
     {slideAddressGen_slideMaskInput_hi[1343:1340]},
     {slideAddressGen_slideMaskInput_hi[1339:1336]},
     {slideAddressGen_slideMaskInput_hi[1335:1332]},
     {slideAddressGen_slideMaskInput_hi[1331:1328]},
     {slideAddressGen_slideMaskInput_hi[1327:1324]},
     {slideAddressGen_slideMaskInput_hi[1323:1320]},
     {slideAddressGen_slideMaskInput_hi[1319:1316]},
     {slideAddressGen_slideMaskInput_hi[1315:1312]},
     {slideAddressGen_slideMaskInput_hi[1311:1308]},
     {slideAddressGen_slideMaskInput_hi[1307:1304]},
     {slideAddressGen_slideMaskInput_hi[1303:1300]},
     {slideAddressGen_slideMaskInput_hi[1299:1296]},
     {slideAddressGen_slideMaskInput_hi[1295:1292]},
     {slideAddressGen_slideMaskInput_hi[1291:1288]},
     {slideAddressGen_slideMaskInput_hi[1287:1284]},
     {slideAddressGen_slideMaskInput_hi[1283:1280]},
     {slideAddressGen_slideMaskInput_hi[1279:1276]},
     {slideAddressGen_slideMaskInput_hi[1275:1272]},
     {slideAddressGen_slideMaskInput_hi[1271:1268]},
     {slideAddressGen_slideMaskInput_hi[1267:1264]},
     {slideAddressGen_slideMaskInput_hi[1263:1260]},
     {slideAddressGen_slideMaskInput_hi[1259:1256]},
     {slideAddressGen_slideMaskInput_hi[1255:1252]},
     {slideAddressGen_slideMaskInput_hi[1251:1248]},
     {slideAddressGen_slideMaskInput_hi[1247:1244]},
     {slideAddressGen_slideMaskInput_hi[1243:1240]},
     {slideAddressGen_slideMaskInput_hi[1239:1236]},
     {slideAddressGen_slideMaskInput_hi[1235:1232]},
     {slideAddressGen_slideMaskInput_hi[1231:1228]},
     {slideAddressGen_slideMaskInput_hi[1227:1224]},
     {slideAddressGen_slideMaskInput_hi[1223:1220]},
     {slideAddressGen_slideMaskInput_hi[1219:1216]},
     {slideAddressGen_slideMaskInput_hi[1215:1212]},
     {slideAddressGen_slideMaskInput_hi[1211:1208]},
     {slideAddressGen_slideMaskInput_hi[1207:1204]},
     {slideAddressGen_slideMaskInput_hi[1203:1200]},
     {slideAddressGen_slideMaskInput_hi[1199:1196]},
     {slideAddressGen_slideMaskInput_hi[1195:1192]},
     {slideAddressGen_slideMaskInput_hi[1191:1188]},
     {slideAddressGen_slideMaskInput_hi[1187:1184]},
     {slideAddressGen_slideMaskInput_hi[1183:1180]},
     {slideAddressGen_slideMaskInput_hi[1179:1176]},
     {slideAddressGen_slideMaskInput_hi[1175:1172]},
     {slideAddressGen_slideMaskInput_hi[1171:1168]},
     {slideAddressGen_slideMaskInput_hi[1167:1164]},
     {slideAddressGen_slideMaskInput_hi[1163:1160]},
     {slideAddressGen_slideMaskInput_hi[1159:1156]},
     {slideAddressGen_slideMaskInput_hi[1155:1152]},
     {slideAddressGen_slideMaskInput_hi[1151:1148]},
     {slideAddressGen_slideMaskInput_hi[1147:1144]},
     {slideAddressGen_slideMaskInput_hi[1143:1140]},
     {slideAddressGen_slideMaskInput_hi[1139:1136]},
     {slideAddressGen_slideMaskInput_hi[1135:1132]},
     {slideAddressGen_slideMaskInput_hi[1131:1128]},
     {slideAddressGen_slideMaskInput_hi[1127:1124]},
     {slideAddressGen_slideMaskInput_hi[1123:1120]},
     {slideAddressGen_slideMaskInput_hi[1119:1116]},
     {slideAddressGen_slideMaskInput_hi[1115:1112]},
     {slideAddressGen_slideMaskInput_hi[1111:1108]},
     {slideAddressGen_slideMaskInput_hi[1107:1104]},
     {slideAddressGen_slideMaskInput_hi[1103:1100]},
     {slideAddressGen_slideMaskInput_hi[1099:1096]},
     {slideAddressGen_slideMaskInput_hi[1095:1092]},
     {slideAddressGen_slideMaskInput_hi[1091:1088]},
     {slideAddressGen_slideMaskInput_hi[1087:1084]},
     {slideAddressGen_slideMaskInput_hi[1083:1080]},
     {slideAddressGen_slideMaskInput_hi[1079:1076]},
     {slideAddressGen_slideMaskInput_hi[1075:1072]},
     {slideAddressGen_slideMaskInput_hi[1071:1068]},
     {slideAddressGen_slideMaskInput_hi[1067:1064]},
     {slideAddressGen_slideMaskInput_hi[1063:1060]},
     {slideAddressGen_slideMaskInput_hi[1059:1056]},
     {slideAddressGen_slideMaskInput_hi[1055:1052]},
     {slideAddressGen_slideMaskInput_hi[1051:1048]},
     {slideAddressGen_slideMaskInput_hi[1047:1044]},
     {slideAddressGen_slideMaskInput_hi[1043:1040]},
     {slideAddressGen_slideMaskInput_hi[1039:1036]},
     {slideAddressGen_slideMaskInput_hi[1035:1032]},
     {slideAddressGen_slideMaskInput_hi[1031:1028]},
     {slideAddressGen_slideMaskInput_hi[1027:1024]},
     {slideAddressGen_slideMaskInput_hi[1023:1020]},
     {slideAddressGen_slideMaskInput_hi[1019:1016]},
     {slideAddressGen_slideMaskInput_hi[1015:1012]},
     {slideAddressGen_slideMaskInput_hi[1011:1008]},
     {slideAddressGen_slideMaskInput_hi[1007:1004]},
     {slideAddressGen_slideMaskInput_hi[1003:1000]},
     {slideAddressGen_slideMaskInput_hi[999:996]},
     {slideAddressGen_slideMaskInput_hi[995:992]},
     {slideAddressGen_slideMaskInput_hi[991:988]},
     {slideAddressGen_slideMaskInput_hi[987:984]},
     {slideAddressGen_slideMaskInput_hi[983:980]},
     {slideAddressGen_slideMaskInput_hi[979:976]},
     {slideAddressGen_slideMaskInput_hi[975:972]},
     {slideAddressGen_slideMaskInput_hi[971:968]},
     {slideAddressGen_slideMaskInput_hi[967:964]},
     {slideAddressGen_slideMaskInput_hi[963:960]},
     {slideAddressGen_slideMaskInput_hi[959:956]},
     {slideAddressGen_slideMaskInput_hi[955:952]},
     {slideAddressGen_slideMaskInput_hi[951:948]},
     {slideAddressGen_slideMaskInput_hi[947:944]},
     {slideAddressGen_slideMaskInput_hi[943:940]},
     {slideAddressGen_slideMaskInput_hi[939:936]},
     {slideAddressGen_slideMaskInput_hi[935:932]},
     {slideAddressGen_slideMaskInput_hi[931:928]},
     {slideAddressGen_slideMaskInput_hi[927:924]},
     {slideAddressGen_slideMaskInput_hi[923:920]},
     {slideAddressGen_slideMaskInput_hi[919:916]},
     {slideAddressGen_slideMaskInput_hi[915:912]},
     {slideAddressGen_slideMaskInput_hi[911:908]},
     {slideAddressGen_slideMaskInput_hi[907:904]},
     {slideAddressGen_slideMaskInput_hi[903:900]},
     {slideAddressGen_slideMaskInput_hi[899:896]},
     {slideAddressGen_slideMaskInput_hi[895:892]},
     {slideAddressGen_slideMaskInput_hi[891:888]},
     {slideAddressGen_slideMaskInput_hi[887:884]},
     {slideAddressGen_slideMaskInput_hi[883:880]},
     {slideAddressGen_slideMaskInput_hi[879:876]},
     {slideAddressGen_slideMaskInput_hi[875:872]},
     {slideAddressGen_slideMaskInput_hi[871:868]},
     {slideAddressGen_slideMaskInput_hi[867:864]},
     {slideAddressGen_slideMaskInput_hi[863:860]},
     {slideAddressGen_slideMaskInput_hi[859:856]},
     {slideAddressGen_slideMaskInput_hi[855:852]},
     {slideAddressGen_slideMaskInput_hi[851:848]},
     {slideAddressGen_slideMaskInput_hi[847:844]},
     {slideAddressGen_slideMaskInput_hi[843:840]},
     {slideAddressGen_slideMaskInput_hi[839:836]},
     {slideAddressGen_slideMaskInput_hi[835:832]},
     {slideAddressGen_slideMaskInput_hi[831:828]},
     {slideAddressGen_slideMaskInput_hi[827:824]},
     {slideAddressGen_slideMaskInput_hi[823:820]},
     {slideAddressGen_slideMaskInput_hi[819:816]},
     {slideAddressGen_slideMaskInput_hi[815:812]},
     {slideAddressGen_slideMaskInput_hi[811:808]},
     {slideAddressGen_slideMaskInput_hi[807:804]},
     {slideAddressGen_slideMaskInput_hi[803:800]},
     {slideAddressGen_slideMaskInput_hi[799:796]},
     {slideAddressGen_slideMaskInput_hi[795:792]},
     {slideAddressGen_slideMaskInput_hi[791:788]},
     {slideAddressGen_slideMaskInput_hi[787:784]},
     {slideAddressGen_slideMaskInput_hi[783:780]},
     {slideAddressGen_slideMaskInput_hi[779:776]},
     {slideAddressGen_slideMaskInput_hi[775:772]},
     {slideAddressGen_slideMaskInput_hi[771:768]},
     {slideAddressGen_slideMaskInput_hi[767:764]},
     {slideAddressGen_slideMaskInput_hi[763:760]},
     {slideAddressGen_slideMaskInput_hi[759:756]},
     {slideAddressGen_slideMaskInput_hi[755:752]},
     {slideAddressGen_slideMaskInput_hi[751:748]},
     {slideAddressGen_slideMaskInput_hi[747:744]},
     {slideAddressGen_slideMaskInput_hi[743:740]},
     {slideAddressGen_slideMaskInput_hi[739:736]},
     {slideAddressGen_slideMaskInput_hi[735:732]},
     {slideAddressGen_slideMaskInput_hi[731:728]},
     {slideAddressGen_slideMaskInput_hi[727:724]},
     {slideAddressGen_slideMaskInput_hi[723:720]},
     {slideAddressGen_slideMaskInput_hi[719:716]},
     {slideAddressGen_slideMaskInput_hi[715:712]},
     {slideAddressGen_slideMaskInput_hi[711:708]},
     {slideAddressGen_slideMaskInput_hi[707:704]},
     {slideAddressGen_slideMaskInput_hi[703:700]},
     {slideAddressGen_slideMaskInput_hi[699:696]},
     {slideAddressGen_slideMaskInput_hi[695:692]},
     {slideAddressGen_slideMaskInput_hi[691:688]},
     {slideAddressGen_slideMaskInput_hi[687:684]},
     {slideAddressGen_slideMaskInput_hi[683:680]},
     {slideAddressGen_slideMaskInput_hi[679:676]},
     {slideAddressGen_slideMaskInput_hi[675:672]},
     {slideAddressGen_slideMaskInput_hi[671:668]},
     {slideAddressGen_slideMaskInput_hi[667:664]},
     {slideAddressGen_slideMaskInput_hi[663:660]},
     {slideAddressGen_slideMaskInput_hi[659:656]},
     {slideAddressGen_slideMaskInput_hi[655:652]},
     {slideAddressGen_slideMaskInput_hi[651:648]},
     {slideAddressGen_slideMaskInput_hi[647:644]},
     {slideAddressGen_slideMaskInput_hi[643:640]},
     {slideAddressGen_slideMaskInput_hi[639:636]},
     {slideAddressGen_slideMaskInput_hi[635:632]},
     {slideAddressGen_slideMaskInput_hi[631:628]},
     {slideAddressGen_slideMaskInput_hi[627:624]},
     {slideAddressGen_slideMaskInput_hi[623:620]},
     {slideAddressGen_slideMaskInput_hi[619:616]},
     {slideAddressGen_slideMaskInput_hi[615:612]},
     {slideAddressGen_slideMaskInput_hi[611:608]},
     {slideAddressGen_slideMaskInput_hi[607:604]},
     {slideAddressGen_slideMaskInput_hi[603:600]},
     {slideAddressGen_slideMaskInput_hi[599:596]},
     {slideAddressGen_slideMaskInput_hi[595:592]},
     {slideAddressGen_slideMaskInput_hi[591:588]},
     {slideAddressGen_slideMaskInput_hi[587:584]},
     {slideAddressGen_slideMaskInput_hi[583:580]},
     {slideAddressGen_slideMaskInput_hi[579:576]},
     {slideAddressGen_slideMaskInput_hi[575:572]},
     {slideAddressGen_slideMaskInput_hi[571:568]},
     {slideAddressGen_slideMaskInput_hi[567:564]},
     {slideAddressGen_slideMaskInput_hi[563:560]},
     {slideAddressGen_slideMaskInput_hi[559:556]},
     {slideAddressGen_slideMaskInput_hi[555:552]},
     {slideAddressGen_slideMaskInput_hi[551:548]},
     {slideAddressGen_slideMaskInput_hi[547:544]},
     {slideAddressGen_slideMaskInput_hi[543:540]},
     {slideAddressGen_slideMaskInput_hi[539:536]},
     {slideAddressGen_slideMaskInput_hi[535:532]},
     {slideAddressGen_slideMaskInput_hi[531:528]},
     {slideAddressGen_slideMaskInput_hi[527:524]},
     {slideAddressGen_slideMaskInput_hi[523:520]},
     {slideAddressGen_slideMaskInput_hi[519:516]},
     {slideAddressGen_slideMaskInput_hi[515:512]},
     {slideAddressGen_slideMaskInput_hi[511:508]},
     {slideAddressGen_slideMaskInput_hi[507:504]},
     {slideAddressGen_slideMaskInput_hi[503:500]},
     {slideAddressGen_slideMaskInput_hi[499:496]},
     {slideAddressGen_slideMaskInput_hi[495:492]},
     {slideAddressGen_slideMaskInput_hi[491:488]},
     {slideAddressGen_slideMaskInput_hi[487:484]},
     {slideAddressGen_slideMaskInput_hi[483:480]},
     {slideAddressGen_slideMaskInput_hi[479:476]},
     {slideAddressGen_slideMaskInput_hi[475:472]},
     {slideAddressGen_slideMaskInput_hi[471:468]},
     {slideAddressGen_slideMaskInput_hi[467:464]},
     {slideAddressGen_slideMaskInput_hi[463:460]},
     {slideAddressGen_slideMaskInput_hi[459:456]},
     {slideAddressGen_slideMaskInput_hi[455:452]},
     {slideAddressGen_slideMaskInput_hi[451:448]},
     {slideAddressGen_slideMaskInput_hi[447:444]},
     {slideAddressGen_slideMaskInput_hi[443:440]},
     {slideAddressGen_slideMaskInput_hi[439:436]},
     {slideAddressGen_slideMaskInput_hi[435:432]},
     {slideAddressGen_slideMaskInput_hi[431:428]},
     {slideAddressGen_slideMaskInput_hi[427:424]},
     {slideAddressGen_slideMaskInput_hi[423:420]},
     {slideAddressGen_slideMaskInput_hi[419:416]},
     {slideAddressGen_slideMaskInput_hi[415:412]},
     {slideAddressGen_slideMaskInput_hi[411:408]},
     {slideAddressGen_slideMaskInput_hi[407:404]},
     {slideAddressGen_slideMaskInput_hi[403:400]},
     {slideAddressGen_slideMaskInput_hi[399:396]},
     {slideAddressGen_slideMaskInput_hi[395:392]},
     {slideAddressGen_slideMaskInput_hi[391:388]},
     {slideAddressGen_slideMaskInput_hi[387:384]},
     {slideAddressGen_slideMaskInput_hi[383:380]},
     {slideAddressGen_slideMaskInput_hi[379:376]},
     {slideAddressGen_slideMaskInput_hi[375:372]},
     {slideAddressGen_slideMaskInput_hi[371:368]},
     {slideAddressGen_slideMaskInput_hi[367:364]},
     {slideAddressGen_slideMaskInput_hi[363:360]},
     {slideAddressGen_slideMaskInput_hi[359:356]},
     {slideAddressGen_slideMaskInput_hi[355:352]},
     {slideAddressGen_slideMaskInput_hi[351:348]},
     {slideAddressGen_slideMaskInput_hi[347:344]},
     {slideAddressGen_slideMaskInput_hi[343:340]},
     {slideAddressGen_slideMaskInput_hi[339:336]},
     {slideAddressGen_slideMaskInput_hi[335:332]},
     {slideAddressGen_slideMaskInput_hi[331:328]},
     {slideAddressGen_slideMaskInput_hi[327:324]},
     {slideAddressGen_slideMaskInput_hi[323:320]},
     {slideAddressGen_slideMaskInput_hi[319:316]},
     {slideAddressGen_slideMaskInput_hi[315:312]},
     {slideAddressGen_slideMaskInput_hi[311:308]},
     {slideAddressGen_slideMaskInput_hi[307:304]},
     {slideAddressGen_slideMaskInput_hi[303:300]},
     {slideAddressGen_slideMaskInput_hi[299:296]},
     {slideAddressGen_slideMaskInput_hi[295:292]},
     {slideAddressGen_slideMaskInput_hi[291:288]},
     {slideAddressGen_slideMaskInput_hi[287:284]},
     {slideAddressGen_slideMaskInput_hi[283:280]},
     {slideAddressGen_slideMaskInput_hi[279:276]},
     {slideAddressGen_slideMaskInput_hi[275:272]},
     {slideAddressGen_slideMaskInput_hi[271:268]},
     {slideAddressGen_slideMaskInput_hi[267:264]},
     {slideAddressGen_slideMaskInput_hi[263:260]},
     {slideAddressGen_slideMaskInput_hi[259:256]},
     {slideAddressGen_slideMaskInput_hi[255:252]},
     {slideAddressGen_slideMaskInput_hi[251:248]},
     {slideAddressGen_slideMaskInput_hi[247:244]},
     {slideAddressGen_slideMaskInput_hi[243:240]},
     {slideAddressGen_slideMaskInput_hi[239:236]},
     {slideAddressGen_slideMaskInput_hi[235:232]},
     {slideAddressGen_slideMaskInput_hi[231:228]},
     {slideAddressGen_slideMaskInput_hi[227:224]},
     {slideAddressGen_slideMaskInput_hi[223:220]},
     {slideAddressGen_slideMaskInput_hi[219:216]},
     {slideAddressGen_slideMaskInput_hi[215:212]},
     {slideAddressGen_slideMaskInput_hi[211:208]},
     {slideAddressGen_slideMaskInput_hi[207:204]},
     {slideAddressGen_slideMaskInput_hi[203:200]},
     {slideAddressGen_slideMaskInput_hi[199:196]},
     {slideAddressGen_slideMaskInput_hi[195:192]},
     {slideAddressGen_slideMaskInput_hi[191:188]},
     {slideAddressGen_slideMaskInput_hi[187:184]},
     {slideAddressGen_slideMaskInput_hi[183:180]},
     {slideAddressGen_slideMaskInput_hi[179:176]},
     {slideAddressGen_slideMaskInput_hi[175:172]},
     {slideAddressGen_slideMaskInput_hi[171:168]},
     {slideAddressGen_slideMaskInput_hi[167:164]},
     {slideAddressGen_slideMaskInput_hi[163:160]},
     {slideAddressGen_slideMaskInput_hi[159:156]},
     {slideAddressGen_slideMaskInput_hi[155:152]},
     {slideAddressGen_slideMaskInput_hi[151:148]},
     {slideAddressGen_slideMaskInput_hi[147:144]},
     {slideAddressGen_slideMaskInput_hi[143:140]},
     {slideAddressGen_slideMaskInput_hi[139:136]},
     {slideAddressGen_slideMaskInput_hi[135:132]},
     {slideAddressGen_slideMaskInput_hi[131:128]},
     {slideAddressGen_slideMaskInput_hi[127:124]},
     {slideAddressGen_slideMaskInput_hi[123:120]},
     {slideAddressGen_slideMaskInput_hi[119:116]},
     {slideAddressGen_slideMaskInput_hi[115:112]},
     {slideAddressGen_slideMaskInput_hi[111:108]},
     {slideAddressGen_slideMaskInput_hi[107:104]},
     {slideAddressGen_slideMaskInput_hi[103:100]},
     {slideAddressGen_slideMaskInput_hi[99:96]},
     {slideAddressGen_slideMaskInput_hi[95:92]},
     {slideAddressGen_slideMaskInput_hi[91:88]},
     {slideAddressGen_slideMaskInput_hi[87:84]},
     {slideAddressGen_slideMaskInput_hi[83:80]},
     {slideAddressGen_slideMaskInput_hi[79:76]},
     {slideAddressGen_slideMaskInput_hi[75:72]},
     {slideAddressGen_slideMaskInput_hi[71:68]},
     {slideAddressGen_slideMaskInput_hi[67:64]},
     {slideAddressGen_slideMaskInput_hi[63:60]},
     {slideAddressGen_slideMaskInput_hi[59:56]},
     {slideAddressGen_slideMaskInput_hi[55:52]},
     {slideAddressGen_slideMaskInput_hi[51:48]},
     {slideAddressGen_slideMaskInput_hi[47:44]},
     {slideAddressGen_slideMaskInput_hi[43:40]},
     {slideAddressGen_slideMaskInput_hi[39:36]},
     {slideAddressGen_slideMaskInput_hi[35:32]},
     {slideAddressGen_slideMaskInput_hi[31:28]},
     {slideAddressGen_slideMaskInput_hi[27:24]},
     {slideAddressGen_slideMaskInput_hi[23:20]},
     {slideAddressGen_slideMaskInput_hi[19:16]},
     {slideAddressGen_slideMaskInput_hi[15:12]},
     {slideAddressGen_slideMaskInput_hi[11:8]},
     {slideAddressGen_slideMaskInput_hi[7:4]},
     {slideAddressGen_slideMaskInput_hi[3:0]},
     {slideAddressGen_slideMaskInput_lo[4095:4092]},
     {slideAddressGen_slideMaskInput_lo[4091:4088]},
     {slideAddressGen_slideMaskInput_lo[4087:4084]},
     {slideAddressGen_slideMaskInput_lo[4083:4080]},
     {slideAddressGen_slideMaskInput_lo[4079:4076]},
     {slideAddressGen_slideMaskInput_lo[4075:4072]},
     {slideAddressGen_slideMaskInput_lo[4071:4068]},
     {slideAddressGen_slideMaskInput_lo[4067:4064]},
     {slideAddressGen_slideMaskInput_lo[4063:4060]},
     {slideAddressGen_slideMaskInput_lo[4059:4056]},
     {slideAddressGen_slideMaskInput_lo[4055:4052]},
     {slideAddressGen_slideMaskInput_lo[4051:4048]},
     {slideAddressGen_slideMaskInput_lo[4047:4044]},
     {slideAddressGen_slideMaskInput_lo[4043:4040]},
     {slideAddressGen_slideMaskInput_lo[4039:4036]},
     {slideAddressGen_slideMaskInput_lo[4035:4032]},
     {slideAddressGen_slideMaskInput_lo[4031:4028]},
     {slideAddressGen_slideMaskInput_lo[4027:4024]},
     {slideAddressGen_slideMaskInput_lo[4023:4020]},
     {slideAddressGen_slideMaskInput_lo[4019:4016]},
     {slideAddressGen_slideMaskInput_lo[4015:4012]},
     {slideAddressGen_slideMaskInput_lo[4011:4008]},
     {slideAddressGen_slideMaskInput_lo[4007:4004]},
     {slideAddressGen_slideMaskInput_lo[4003:4000]},
     {slideAddressGen_slideMaskInput_lo[3999:3996]},
     {slideAddressGen_slideMaskInput_lo[3995:3992]},
     {slideAddressGen_slideMaskInput_lo[3991:3988]},
     {slideAddressGen_slideMaskInput_lo[3987:3984]},
     {slideAddressGen_slideMaskInput_lo[3983:3980]},
     {slideAddressGen_slideMaskInput_lo[3979:3976]},
     {slideAddressGen_slideMaskInput_lo[3975:3972]},
     {slideAddressGen_slideMaskInput_lo[3971:3968]},
     {slideAddressGen_slideMaskInput_lo[3967:3964]},
     {slideAddressGen_slideMaskInput_lo[3963:3960]},
     {slideAddressGen_slideMaskInput_lo[3959:3956]},
     {slideAddressGen_slideMaskInput_lo[3955:3952]},
     {slideAddressGen_slideMaskInput_lo[3951:3948]},
     {slideAddressGen_slideMaskInput_lo[3947:3944]},
     {slideAddressGen_slideMaskInput_lo[3943:3940]},
     {slideAddressGen_slideMaskInput_lo[3939:3936]},
     {slideAddressGen_slideMaskInput_lo[3935:3932]},
     {slideAddressGen_slideMaskInput_lo[3931:3928]},
     {slideAddressGen_slideMaskInput_lo[3927:3924]},
     {slideAddressGen_slideMaskInput_lo[3923:3920]},
     {slideAddressGen_slideMaskInput_lo[3919:3916]},
     {slideAddressGen_slideMaskInput_lo[3915:3912]},
     {slideAddressGen_slideMaskInput_lo[3911:3908]},
     {slideAddressGen_slideMaskInput_lo[3907:3904]},
     {slideAddressGen_slideMaskInput_lo[3903:3900]},
     {slideAddressGen_slideMaskInput_lo[3899:3896]},
     {slideAddressGen_slideMaskInput_lo[3895:3892]},
     {slideAddressGen_slideMaskInput_lo[3891:3888]},
     {slideAddressGen_slideMaskInput_lo[3887:3884]},
     {slideAddressGen_slideMaskInput_lo[3883:3880]},
     {slideAddressGen_slideMaskInput_lo[3879:3876]},
     {slideAddressGen_slideMaskInput_lo[3875:3872]},
     {slideAddressGen_slideMaskInput_lo[3871:3868]},
     {slideAddressGen_slideMaskInput_lo[3867:3864]},
     {slideAddressGen_slideMaskInput_lo[3863:3860]},
     {slideAddressGen_slideMaskInput_lo[3859:3856]},
     {slideAddressGen_slideMaskInput_lo[3855:3852]},
     {slideAddressGen_slideMaskInput_lo[3851:3848]},
     {slideAddressGen_slideMaskInput_lo[3847:3844]},
     {slideAddressGen_slideMaskInput_lo[3843:3840]},
     {slideAddressGen_slideMaskInput_lo[3839:3836]},
     {slideAddressGen_slideMaskInput_lo[3835:3832]},
     {slideAddressGen_slideMaskInput_lo[3831:3828]},
     {slideAddressGen_slideMaskInput_lo[3827:3824]},
     {slideAddressGen_slideMaskInput_lo[3823:3820]},
     {slideAddressGen_slideMaskInput_lo[3819:3816]},
     {slideAddressGen_slideMaskInput_lo[3815:3812]},
     {slideAddressGen_slideMaskInput_lo[3811:3808]},
     {slideAddressGen_slideMaskInput_lo[3807:3804]},
     {slideAddressGen_slideMaskInput_lo[3803:3800]},
     {slideAddressGen_slideMaskInput_lo[3799:3796]},
     {slideAddressGen_slideMaskInput_lo[3795:3792]},
     {slideAddressGen_slideMaskInput_lo[3791:3788]},
     {slideAddressGen_slideMaskInput_lo[3787:3784]},
     {slideAddressGen_slideMaskInput_lo[3783:3780]},
     {slideAddressGen_slideMaskInput_lo[3779:3776]},
     {slideAddressGen_slideMaskInput_lo[3775:3772]},
     {slideAddressGen_slideMaskInput_lo[3771:3768]},
     {slideAddressGen_slideMaskInput_lo[3767:3764]},
     {slideAddressGen_slideMaskInput_lo[3763:3760]},
     {slideAddressGen_slideMaskInput_lo[3759:3756]},
     {slideAddressGen_slideMaskInput_lo[3755:3752]},
     {slideAddressGen_slideMaskInput_lo[3751:3748]},
     {slideAddressGen_slideMaskInput_lo[3747:3744]},
     {slideAddressGen_slideMaskInput_lo[3743:3740]},
     {slideAddressGen_slideMaskInput_lo[3739:3736]},
     {slideAddressGen_slideMaskInput_lo[3735:3732]},
     {slideAddressGen_slideMaskInput_lo[3731:3728]},
     {slideAddressGen_slideMaskInput_lo[3727:3724]},
     {slideAddressGen_slideMaskInput_lo[3723:3720]},
     {slideAddressGen_slideMaskInput_lo[3719:3716]},
     {slideAddressGen_slideMaskInput_lo[3715:3712]},
     {slideAddressGen_slideMaskInput_lo[3711:3708]},
     {slideAddressGen_slideMaskInput_lo[3707:3704]},
     {slideAddressGen_slideMaskInput_lo[3703:3700]},
     {slideAddressGen_slideMaskInput_lo[3699:3696]},
     {slideAddressGen_slideMaskInput_lo[3695:3692]},
     {slideAddressGen_slideMaskInput_lo[3691:3688]},
     {slideAddressGen_slideMaskInput_lo[3687:3684]},
     {slideAddressGen_slideMaskInput_lo[3683:3680]},
     {slideAddressGen_slideMaskInput_lo[3679:3676]},
     {slideAddressGen_slideMaskInput_lo[3675:3672]},
     {slideAddressGen_slideMaskInput_lo[3671:3668]},
     {slideAddressGen_slideMaskInput_lo[3667:3664]},
     {slideAddressGen_slideMaskInput_lo[3663:3660]},
     {slideAddressGen_slideMaskInput_lo[3659:3656]},
     {slideAddressGen_slideMaskInput_lo[3655:3652]},
     {slideAddressGen_slideMaskInput_lo[3651:3648]},
     {slideAddressGen_slideMaskInput_lo[3647:3644]},
     {slideAddressGen_slideMaskInput_lo[3643:3640]},
     {slideAddressGen_slideMaskInput_lo[3639:3636]},
     {slideAddressGen_slideMaskInput_lo[3635:3632]},
     {slideAddressGen_slideMaskInput_lo[3631:3628]},
     {slideAddressGen_slideMaskInput_lo[3627:3624]},
     {slideAddressGen_slideMaskInput_lo[3623:3620]},
     {slideAddressGen_slideMaskInput_lo[3619:3616]},
     {slideAddressGen_slideMaskInput_lo[3615:3612]},
     {slideAddressGen_slideMaskInput_lo[3611:3608]},
     {slideAddressGen_slideMaskInput_lo[3607:3604]},
     {slideAddressGen_slideMaskInput_lo[3603:3600]},
     {slideAddressGen_slideMaskInput_lo[3599:3596]},
     {slideAddressGen_slideMaskInput_lo[3595:3592]},
     {slideAddressGen_slideMaskInput_lo[3591:3588]},
     {slideAddressGen_slideMaskInput_lo[3587:3584]},
     {slideAddressGen_slideMaskInput_lo[3583:3580]},
     {slideAddressGen_slideMaskInput_lo[3579:3576]},
     {slideAddressGen_slideMaskInput_lo[3575:3572]},
     {slideAddressGen_slideMaskInput_lo[3571:3568]},
     {slideAddressGen_slideMaskInput_lo[3567:3564]},
     {slideAddressGen_slideMaskInput_lo[3563:3560]},
     {slideAddressGen_slideMaskInput_lo[3559:3556]},
     {slideAddressGen_slideMaskInput_lo[3555:3552]},
     {slideAddressGen_slideMaskInput_lo[3551:3548]},
     {slideAddressGen_slideMaskInput_lo[3547:3544]},
     {slideAddressGen_slideMaskInput_lo[3543:3540]},
     {slideAddressGen_slideMaskInput_lo[3539:3536]},
     {slideAddressGen_slideMaskInput_lo[3535:3532]},
     {slideAddressGen_slideMaskInput_lo[3531:3528]},
     {slideAddressGen_slideMaskInput_lo[3527:3524]},
     {slideAddressGen_slideMaskInput_lo[3523:3520]},
     {slideAddressGen_slideMaskInput_lo[3519:3516]},
     {slideAddressGen_slideMaskInput_lo[3515:3512]},
     {slideAddressGen_slideMaskInput_lo[3511:3508]},
     {slideAddressGen_slideMaskInput_lo[3507:3504]},
     {slideAddressGen_slideMaskInput_lo[3503:3500]},
     {slideAddressGen_slideMaskInput_lo[3499:3496]},
     {slideAddressGen_slideMaskInput_lo[3495:3492]},
     {slideAddressGen_slideMaskInput_lo[3491:3488]},
     {slideAddressGen_slideMaskInput_lo[3487:3484]},
     {slideAddressGen_slideMaskInput_lo[3483:3480]},
     {slideAddressGen_slideMaskInput_lo[3479:3476]},
     {slideAddressGen_slideMaskInput_lo[3475:3472]},
     {slideAddressGen_slideMaskInput_lo[3471:3468]},
     {slideAddressGen_slideMaskInput_lo[3467:3464]},
     {slideAddressGen_slideMaskInput_lo[3463:3460]},
     {slideAddressGen_slideMaskInput_lo[3459:3456]},
     {slideAddressGen_slideMaskInput_lo[3455:3452]},
     {slideAddressGen_slideMaskInput_lo[3451:3448]},
     {slideAddressGen_slideMaskInput_lo[3447:3444]},
     {slideAddressGen_slideMaskInput_lo[3443:3440]},
     {slideAddressGen_slideMaskInput_lo[3439:3436]},
     {slideAddressGen_slideMaskInput_lo[3435:3432]},
     {slideAddressGen_slideMaskInput_lo[3431:3428]},
     {slideAddressGen_slideMaskInput_lo[3427:3424]},
     {slideAddressGen_slideMaskInput_lo[3423:3420]},
     {slideAddressGen_slideMaskInput_lo[3419:3416]},
     {slideAddressGen_slideMaskInput_lo[3415:3412]},
     {slideAddressGen_slideMaskInput_lo[3411:3408]},
     {slideAddressGen_slideMaskInput_lo[3407:3404]},
     {slideAddressGen_slideMaskInput_lo[3403:3400]},
     {slideAddressGen_slideMaskInput_lo[3399:3396]},
     {slideAddressGen_slideMaskInput_lo[3395:3392]},
     {slideAddressGen_slideMaskInput_lo[3391:3388]},
     {slideAddressGen_slideMaskInput_lo[3387:3384]},
     {slideAddressGen_slideMaskInput_lo[3383:3380]},
     {slideAddressGen_slideMaskInput_lo[3379:3376]},
     {slideAddressGen_slideMaskInput_lo[3375:3372]},
     {slideAddressGen_slideMaskInput_lo[3371:3368]},
     {slideAddressGen_slideMaskInput_lo[3367:3364]},
     {slideAddressGen_slideMaskInput_lo[3363:3360]},
     {slideAddressGen_slideMaskInput_lo[3359:3356]},
     {slideAddressGen_slideMaskInput_lo[3355:3352]},
     {slideAddressGen_slideMaskInput_lo[3351:3348]},
     {slideAddressGen_slideMaskInput_lo[3347:3344]},
     {slideAddressGen_slideMaskInput_lo[3343:3340]},
     {slideAddressGen_slideMaskInput_lo[3339:3336]},
     {slideAddressGen_slideMaskInput_lo[3335:3332]},
     {slideAddressGen_slideMaskInput_lo[3331:3328]},
     {slideAddressGen_slideMaskInput_lo[3327:3324]},
     {slideAddressGen_slideMaskInput_lo[3323:3320]},
     {slideAddressGen_slideMaskInput_lo[3319:3316]},
     {slideAddressGen_slideMaskInput_lo[3315:3312]},
     {slideAddressGen_slideMaskInput_lo[3311:3308]},
     {slideAddressGen_slideMaskInput_lo[3307:3304]},
     {slideAddressGen_slideMaskInput_lo[3303:3300]},
     {slideAddressGen_slideMaskInput_lo[3299:3296]},
     {slideAddressGen_slideMaskInput_lo[3295:3292]},
     {slideAddressGen_slideMaskInput_lo[3291:3288]},
     {slideAddressGen_slideMaskInput_lo[3287:3284]},
     {slideAddressGen_slideMaskInput_lo[3283:3280]},
     {slideAddressGen_slideMaskInput_lo[3279:3276]},
     {slideAddressGen_slideMaskInput_lo[3275:3272]},
     {slideAddressGen_slideMaskInput_lo[3271:3268]},
     {slideAddressGen_slideMaskInput_lo[3267:3264]},
     {slideAddressGen_slideMaskInput_lo[3263:3260]},
     {slideAddressGen_slideMaskInput_lo[3259:3256]},
     {slideAddressGen_slideMaskInput_lo[3255:3252]},
     {slideAddressGen_slideMaskInput_lo[3251:3248]},
     {slideAddressGen_slideMaskInput_lo[3247:3244]},
     {slideAddressGen_slideMaskInput_lo[3243:3240]},
     {slideAddressGen_slideMaskInput_lo[3239:3236]},
     {slideAddressGen_slideMaskInput_lo[3235:3232]},
     {slideAddressGen_slideMaskInput_lo[3231:3228]},
     {slideAddressGen_slideMaskInput_lo[3227:3224]},
     {slideAddressGen_slideMaskInput_lo[3223:3220]},
     {slideAddressGen_slideMaskInput_lo[3219:3216]},
     {slideAddressGen_slideMaskInput_lo[3215:3212]},
     {slideAddressGen_slideMaskInput_lo[3211:3208]},
     {slideAddressGen_slideMaskInput_lo[3207:3204]},
     {slideAddressGen_slideMaskInput_lo[3203:3200]},
     {slideAddressGen_slideMaskInput_lo[3199:3196]},
     {slideAddressGen_slideMaskInput_lo[3195:3192]},
     {slideAddressGen_slideMaskInput_lo[3191:3188]},
     {slideAddressGen_slideMaskInput_lo[3187:3184]},
     {slideAddressGen_slideMaskInput_lo[3183:3180]},
     {slideAddressGen_slideMaskInput_lo[3179:3176]},
     {slideAddressGen_slideMaskInput_lo[3175:3172]},
     {slideAddressGen_slideMaskInput_lo[3171:3168]},
     {slideAddressGen_slideMaskInput_lo[3167:3164]},
     {slideAddressGen_slideMaskInput_lo[3163:3160]},
     {slideAddressGen_slideMaskInput_lo[3159:3156]},
     {slideAddressGen_slideMaskInput_lo[3155:3152]},
     {slideAddressGen_slideMaskInput_lo[3151:3148]},
     {slideAddressGen_slideMaskInput_lo[3147:3144]},
     {slideAddressGen_slideMaskInput_lo[3143:3140]},
     {slideAddressGen_slideMaskInput_lo[3139:3136]},
     {slideAddressGen_slideMaskInput_lo[3135:3132]},
     {slideAddressGen_slideMaskInput_lo[3131:3128]},
     {slideAddressGen_slideMaskInput_lo[3127:3124]},
     {slideAddressGen_slideMaskInput_lo[3123:3120]},
     {slideAddressGen_slideMaskInput_lo[3119:3116]},
     {slideAddressGen_slideMaskInput_lo[3115:3112]},
     {slideAddressGen_slideMaskInput_lo[3111:3108]},
     {slideAddressGen_slideMaskInput_lo[3107:3104]},
     {slideAddressGen_slideMaskInput_lo[3103:3100]},
     {slideAddressGen_slideMaskInput_lo[3099:3096]},
     {slideAddressGen_slideMaskInput_lo[3095:3092]},
     {slideAddressGen_slideMaskInput_lo[3091:3088]},
     {slideAddressGen_slideMaskInput_lo[3087:3084]},
     {slideAddressGen_slideMaskInput_lo[3083:3080]},
     {slideAddressGen_slideMaskInput_lo[3079:3076]},
     {slideAddressGen_slideMaskInput_lo[3075:3072]},
     {slideAddressGen_slideMaskInput_lo[3071:3068]},
     {slideAddressGen_slideMaskInput_lo[3067:3064]},
     {slideAddressGen_slideMaskInput_lo[3063:3060]},
     {slideAddressGen_slideMaskInput_lo[3059:3056]},
     {slideAddressGen_slideMaskInput_lo[3055:3052]},
     {slideAddressGen_slideMaskInput_lo[3051:3048]},
     {slideAddressGen_slideMaskInput_lo[3047:3044]},
     {slideAddressGen_slideMaskInput_lo[3043:3040]},
     {slideAddressGen_slideMaskInput_lo[3039:3036]},
     {slideAddressGen_slideMaskInput_lo[3035:3032]},
     {slideAddressGen_slideMaskInput_lo[3031:3028]},
     {slideAddressGen_slideMaskInput_lo[3027:3024]},
     {slideAddressGen_slideMaskInput_lo[3023:3020]},
     {slideAddressGen_slideMaskInput_lo[3019:3016]},
     {slideAddressGen_slideMaskInput_lo[3015:3012]},
     {slideAddressGen_slideMaskInput_lo[3011:3008]},
     {slideAddressGen_slideMaskInput_lo[3007:3004]},
     {slideAddressGen_slideMaskInput_lo[3003:3000]},
     {slideAddressGen_slideMaskInput_lo[2999:2996]},
     {slideAddressGen_slideMaskInput_lo[2995:2992]},
     {slideAddressGen_slideMaskInput_lo[2991:2988]},
     {slideAddressGen_slideMaskInput_lo[2987:2984]},
     {slideAddressGen_slideMaskInput_lo[2983:2980]},
     {slideAddressGen_slideMaskInput_lo[2979:2976]},
     {slideAddressGen_slideMaskInput_lo[2975:2972]},
     {slideAddressGen_slideMaskInput_lo[2971:2968]},
     {slideAddressGen_slideMaskInput_lo[2967:2964]},
     {slideAddressGen_slideMaskInput_lo[2963:2960]},
     {slideAddressGen_slideMaskInput_lo[2959:2956]},
     {slideAddressGen_slideMaskInput_lo[2955:2952]},
     {slideAddressGen_slideMaskInput_lo[2951:2948]},
     {slideAddressGen_slideMaskInput_lo[2947:2944]},
     {slideAddressGen_slideMaskInput_lo[2943:2940]},
     {slideAddressGen_slideMaskInput_lo[2939:2936]},
     {slideAddressGen_slideMaskInput_lo[2935:2932]},
     {slideAddressGen_slideMaskInput_lo[2931:2928]},
     {slideAddressGen_slideMaskInput_lo[2927:2924]},
     {slideAddressGen_slideMaskInput_lo[2923:2920]},
     {slideAddressGen_slideMaskInput_lo[2919:2916]},
     {slideAddressGen_slideMaskInput_lo[2915:2912]},
     {slideAddressGen_slideMaskInput_lo[2911:2908]},
     {slideAddressGen_slideMaskInput_lo[2907:2904]},
     {slideAddressGen_slideMaskInput_lo[2903:2900]},
     {slideAddressGen_slideMaskInput_lo[2899:2896]},
     {slideAddressGen_slideMaskInput_lo[2895:2892]},
     {slideAddressGen_slideMaskInput_lo[2891:2888]},
     {slideAddressGen_slideMaskInput_lo[2887:2884]},
     {slideAddressGen_slideMaskInput_lo[2883:2880]},
     {slideAddressGen_slideMaskInput_lo[2879:2876]},
     {slideAddressGen_slideMaskInput_lo[2875:2872]},
     {slideAddressGen_slideMaskInput_lo[2871:2868]},
     {slideAddressGen_slideMaskInput_lo[2867:2864]},
     {slideAddressGen_slideMaskInput_lo[2863:2860]},
     {slideAddressGen_slideMaskInput_lo[2859:2856]},
     {slideAddressGen_slideMaskInput_lo[2855:2852]},
     {slideAddressGen_slideMaskInput_lo[2851:2848]},
     {slideAddressGen_slideMaskInput_lo[2847:2844]},
     {slideAddressGen_slideMaskInput_lo[2843:2840]},
     {slideAddressGen_slideMaskInput_lo[2839:2836]},
     {slideAddressGen_slideMaskInput_lo[2835:2832]},
     {slideAddressGen_slideMaskInput_lo[2831:2828]},
     {slideAddressGen_slideMaskInput_lo[2827:2824]},
     {slideAddressGen_slideMaskInput_lo[2823:2820]},
     {slideAddressGen_slideMaskInput_lo[2819:2816]},
     {slideAddressGen_slideMaskInput_lo[2815:2812]},
     {slideAddressGen_slideMaskInput_lo[2811:2808]},
     {slideAddressGen_slideMaskInput_lo[2807:2804]},
     {slideAddressGen_slideMaskInput_lo[2803:2800]},
     {slideAddressGen_slideMaskInput_lo[2799:2796]},
     {slideAddressGen_slideMaskInput_lo[2795:2792]},
     {slideAddressGen_slideMaskInput_lo[2791:2788]},
     {slideAddressGen_slideMaskInput_lo[2787:2784]},
     {slideAddressGen_slideMaskInput_lo[2783:2780]},
     {slideAddressGen_slideMaskInput_lo[2779:2776]},
     {slideAddressGen_slideMaskInput_lo[2775:2772]},
     {slideAddressGen_slideMaskInput_lo[2771:2768]},
     {slideAddressGen_slideMaskInput_lo[2767:2764]},
     {slideAddressGen_slideMaskInput_lo[2763:2760]},
     {slideAddressGen_slideMaskInput_lo[2759:2756]},
     {slideAddressGen_slideMaskInput_lo[2755:2752]},
     {slideAddressGen_slideMaskInput_lo[2751:2748]},
     {slideAddressGen_slideMaskInput_lo[2747:2744]},
     {slideAddressGen_slideMaskInput_lo[2743:2740]},
     {slideAddressGen_slideMaskInput_lo[2739:2736]},
     {slideAddressGen_slideMaskInput_lo[2735:2732]},
     {slideAddressGen_slideMaskInput_lo[2731:2728]},
     {slideAddressGen_slideMaskInput_lo[2727:2724]},
     {slideAddressGen_slideMaskInput_lo[2723:2720]},
     {slideAddressGen_slideMaskInput_lo[2719:2716]},
     {slideAddressGen_slideMaskInput_lo[2715:2712]},
     {slideAddressGen_slideMaskInput_lo[2711:2708]},
     {slideAddressGen_slideMaskInput_lo[2707:2704]},
     {slideAddressGen_slideMaskInput_lo[2703:2700]},
     {slideAddressGen_slideMaskInput_lo[2699:2696]},
     {slideAddressGen_slideMaskInput_lo[2695:2692]},
     {slideAddressGen_slideMaskInput_lo[2691:2688]},
     {slideAddressGen_slideMaskInput_lo[2687:2684]},
     {slideAddressGen_slideMaskInput_lo[2683:2680]},
     {slideAddressGen_slideMaskInput_lo[2679:2676]},
     {slideAddressGen_slideMaskInput_lo[2675:2672]},
     {slideAddressGen_slideMaskInput_lo[2671:2668]},
     {slideAddressGen_slideMaskInput_lo[2667:2664]},
     {slideAddressGen_slideMaskInput_lo[2663:2660]},
     {slideAddressGen_slideMaskInput_lo[2659:2656]},
     {slideAddressGen_slideMaskInput_lo[2655:2652]},
     {slideAddressGen_slideMaskInput_lo[2651:2648]},
     {slideAddressGen_slideMaskInput_lo[2647:2644]},
     {slideAddressGen_slideMaskInput_lo[2643:2640]},
     {slideAddressGen_slideMaskInput_lo[2639:2636]},
     {slideAddressGen_slideMaskInput_lo[2635:2632]},
     {slideAddressGen_slideMaskInput_lo[2631:2628]},
     {slideAddressGen_slideMaskInput_lo[2627:2624]},
     {slideAddressGen_slideMaskInput_lo[2623:2620]},
     {slideAddressGen_slideMaskInput_lo[2619:2616]},
     {slideAddressGen_slideMaskInput_lo[2615:2612]},
     {slideAddressGen_slideMaskInput_lo[2611:2608]},
     {slideAddressGen_slideMaskInput_lo[2607:2604]},
     {slideAddressGen_slideMaskInput_lo[2603:2600]},
     {slideAddressGen_slideMaskInput_lo[2599:2596]},
     {slideAddressGen_slideMaskInput_lo[2595:2592]},
     {slideAddressGen_slideMaskInput_lo[2591:2588]},
     {slideAddressGen_slideMaskInput_lo[2587:2584]},
     {slideAddressGen_slideMaskInput_lo[2583:2580]},
     {slideAddressGen_slideMaskInput_lo[2579:2576]},
     {slideAddressGen_slideMaskInput_lo[2575:2572]},
     {slideAddressGen_slideMaskInput_lo[2571:2568]},
     {slideAddressGen_slideMaskInput_lo[2567:2564]},
     {slideAddressGen_slideMaskInput_lo[2563:2560]},
     {slideAddressGen_slideMaskInput_lo[2559:2556]},
     {slideAddressGen_slideMaskInput_lo[2555:2552]},
     {slideAddressGen_slideMaskInput_lo[2551:2548]},
     {slideAddressGen_slideMaskInput_lo[2547:2544]},
     {slideAddressGen_slideMaskInput_lo[2543:2540]},
     {slideAddressGen_slideMaskInput_lo[2539:2536]},
     {slideAddressGen_slideMaskInput_lo[2535:2532]},
     {slideAddressGen_slideMaskInput_lo[2531:2528]},
     {slideAddressGen_slideMaskInput_lo[2527:2524]},
     {slideAddressGen_slideMaskInput_lo[2523:2520]},
     {slideAddressGen_slideMaskInput_lo[2519:2516]},
     {slideAddressGen_slideMaskInput_lo[2515:2512]},
     {slideAddressGen_slideMaskInput_lo[2511:2508]},
     {slideAddressGen_slideMaskInput_lo[2507:2504]},
     {slideAddressGen_slideMaskInput_lo[2503:2500]},
     {slideAddressGen_slideMaskInput_lo[2499:2496]},
     {slideAddressGen_slideMaskInput_lo[2495:2492]},
     {slideAddressGen_slideMaskInput_lo[2491:2488]},
     {slideAddressGen_slideMaskInput_lo[2487:2484]},
     {slideAddressGen_slideMaskInput_lo[2483:2480]},
     {slideAddressGen_slideMaskInput_lo[2479:2476]},
     {slideAddressGen_slideMaskInput_lo[2475:2472]},
     {slideAddressGen_slideMaskInput_lo[2471:2468]},
     {slideAddressGen_slideMaskInput_lo[2467:2464]},
     {slideAddressGen_slideMaskInput_lo[2463:2460]},
     {slideAddressGen_slideMaskInput_lo[2459:2456]},
     {slideAddressGen_slideMaskInput_lo[2455:2452]},
     {slideAddressGen_slideMaskInput_lo[2451:2448]},
     {slideAddressGen_slideMaskInput_lo[2447:2444]},
     {slideAddressGen_slideMaskInput_lo[2443:2440]},
     {slideAddressGen_slideMaskInput_lo[2439:2436]},
     {slideAddressGen_slideMaskInput_lo[2435:2432]},
     {slideAddressGen_slideMaskInput_lo[2431:2428]},
     {slideAddressGen_slideMaskInput_lo[2427:2424]},
     {slideAddressGen_slideMaskInput_lo[2423:2420]},
     {slideAddressGen_slideMaskInput_lo[2419:2416]},
     {slideAddressGen_slideMaskInput_lo[2415:2412]},
     {slideAddressGen_slideMaskInput_lo[2411:2408]},
     {slideAddressGen_slideMaskInput_lo[2407:2404]},
     {slideAddressGen_slideMaskInput_lo[2403:2400]},
     {slideAddressGen_slideMaskInput_lo[2399:2396]},
     {slideAddressGen_slideMaskInput_lo[2395:2392]},
     {slideAddressGen_slideMaskInput_lo[2391:2388]},
     {slideAddressGen_slideMaskInput_lo[2387:2384]},
     {slideAddressGen_slideMaskInput_lo[2383:2380]},
     {slideAddressGen_slideMaskInput_lo[2379:2376]},
     {slideAddressGen_slideMaskInput_lo[2375:2372]},
     {slideAddressGen_slideMaskInput_lo[2371:2368]},
     {slideAddressGen_slideMaskInput_lo[2367:2364]},
     {slideAddressGen_slideMaskInput_lo[2363:2360]},
     {slideAddressGen_slideMaskInput_lo[2359:2356]},
     {slideAddressGen_slideMaskInput_lo[2355:2352]},
     {slideAddressGen_slideMaskInput_lo[2351:2348]},
     {slideAddressGen_slideMaskInput_lo[2347:2344]},
     {slideAddressGen_slideMaskInput_lo[2343:2340]},
     {slideAddressGen_slideMaskInput_lo[2339:2336]},
     {slideAddressGen_slideMaskInput_lo[2335:2332]},
     {slideAddressGen_slideMaskInput_lo[2331:2328]},
     {slideAddressGen_slideMaskInput_lo[2327:2324]},
     {slideAddressGen_slideMaskInput_lo[2323:2320]},
     {slideAddressGen_slideMaskInput_lo[2319:2316]},
     {slideAddressGen_slideMaskInput_lo[2315:2312]},
     {slideAddressGen_slideMaskInput_lo[2311:2308]},
     {slideAddressGen_slideMaskInput_lo[2307:2304]},
     {slideAddressGen_slideMaskInput_lo[2303:2300]},
     {slideAddressGen_slideMaskInput_lo[2299:2296]},
     {slideAddressGen_slideMaskInput_lo[2295:2292]},
     {slideAddressGen_slideMaskInput_lo[2291:2288]},
     {slideAddressGen_slideMaskInput_lo[2287:2284]},
     {slideAddressGen_slideMaskInput_lo[2283:2280]},
     {slideAddressGen_slideMaskInput_lo[2279:2276]},
     {slideAddressGen_slideMaskInput_lo[2275:2272]},
     {slideAddressGen_slideMaskInput_lo[2271:2268]},
     {slideAddressGen_slideMaskInput_lo[2267:2264]},
     {slideAddressGen_slideMaskInput_lo[2263:2260]},
     {slideAddressGen_slideMaskInput_lo[2259:2256]},
     {slideAddressGen_slideMaskInput_lo[2255:2252]},
     {slideAddressGen_slideMaskInput_lo[2251:2248]},
     {slideAddressGen_slideMaskInput_lo[2247:2244]},
     {slideAddressGen_slideMaskInput_lo[2243:2240]},
     {slideAddressGen_slideMaskInput_lo[2239:2236]},
     {slideAddressGen_slideMaskInput_lo[2235:2232]},
     {slideAddressGen_slideMaskInput_lo[2231:2228]},
     {slideAddressGen_slideMaskInput_lo[2227:2224]},
     {slideAddressGen_slideMaskInput_lo[2223:2220]},
     {slideAddressGen_slideMaskInput_lo[2219:2216]},
     {slideAddressGen_slideMaskInput_lo[2215:2212]},
     {slideAddressGen_slideMaskInput_lo[2211:2208]},
     {slideAddressGen_slideMaskInput_lo[2207:2204]},
     {slideAddressGen_slideMaskInput_lo[2203:2200]},
     {slideAddressGen_slideMaskInput_lo[2199:2196]},
     {slideAddressGen_slideMaskInput_lo[2195:2192]},
     {slideAddressGen_slideMaskInput_lo[2191:2188]},
     {slideAddressGen_slideMaskInput_lo[2187:2184]},
     {slideAddressGen_slideMaskInput_lo[2183:2180]},
     {slideAddressGen_slideMaskInput_lo[2179:2176]},
     {slideAddressGen_slideMaskInput_lo[2175:2172]},
     {slideAddressGen_slideMaskInput_lo[2171:2168]},
     {slideAddressGen_slideMaskInput_lo[2167:2164]},
     {slideAddressGen_slideMaskInput_lo[2163:2160]},
     {slideAddressGen_slideMaskInput_lo[2159:2156]},
     {slideAddressGen_slideMaskInput_lo[2155:2152]},
     {slideAddressGen_slideMaskInput_lo[2151:2148]},
     {slideAddressGen_slideMaskInput_lo[2147:2144]},
     {slideAddressGen_slideMaskInput_lo[2143:2140]},
     {slideAddressGen_slideMaskInput_lo[2139:2136]},
     {slideAddressGen_slideMaskInput_lo[2135:2132]},
     {slideAddressGen_slideMaskInput_lo[2131:2128]},
     {slideAddressGen_slideMaskInput_lo[2127:2124]},
     {slideAddressGen_slideMaskInput_lo[2123:2120]},
     {slideAddressGen_slideMaskInput_lo[2119:2116]},
     {slideAddressGen_slideMaskInput_lo[2115:2112]},
     {slideAddressGen_slideMaskInput_lo[2111:2108]},
     {slideAddressGen_slideMaskInput_lo[2107:2104]},
     {slideAddressGen_slideMaskInput_lo[2103:2100]},
     {slideAddressGen_slideMaskInput_lo[2099:2096]},
     {slideAddressGen_slideMaskInput_lo[2095:2092]},
     {slideAddressGen_slideMaskInput_lo[2091:2088]},
     {slideAddressGen_slideMaskInput_lo[2087:2084]},
     {slideAddressGen_slideMaskInput_lo[2083:2080]},
     {slideAddressGen_slideMaskInput_lo[2079:2076]},
     {slideAddressGen_slideMaskInput_lo[2075:2072]},
     {slideAddressGen_slideMaskInput_lo[2071:2068]},
     {slideAddressGen_slideMaskInput_lo[2067:2064]},
     {slideAddressGen_slideMaskInput_lo[2063:2060]},
     {slideAddressGen_slideMaskInput_lo[2059:2056]},
     {slideAddressGen_slideMaskInput_lo[2055:2052]},
     {slideAddressGen_slideMaskInput_lo[2051:2048]},
     {slideAddressGen_slideMaskInput_lo[2047:2044]},
     {slideAddressGen_slideMaskInput_lo[2043:2040]},
     {slideAddressGen_slideMaskInput_lo[2039:2036]},
     {slideAddressGen_slideMaskInput_lo[2035:2032]},
     {slideAddressGen_slideMaskInput_lo[2031:2028]},
     {slideAddressGen_slideMaskInput_lo[2027:2024]},
     {slideAddressGen_slideMaskInput_lo[2023:2020]},
     {slideAddressGen_slideMaskInput_lo[2019:2016]},
     {slideAddressGen_slideMaskInput_lo[2015:2012]},
     {slideAddressGen_slideMaskInput_lo[2011:2008]},
     {slideAddressGen_slideMaskInput_lo[2007:2004]},
     {slideAddressGen_slideMaskInput_lo[2003:2000]},
     {slideAddressGen_slideMaskInput_lo[1999:1996]},
     {slideAddressGen_slideMaskInput_lo[1995:1992]},
     {slideAddressGen_slideMaskInput_lo[1991:1988]},
     {slideAddressGen_slideMaskInput_lo[1987:1984]},
     {slideAddressGen_slideMaskInput_lo[1983:1980]},
     {slideAddressGen_slideMaskInput_lo[1979:1976]},
     {slideAddressGen_slideMaskInput_lo[1975:1972]},
     {slideAddressGen_slideMaskInput_lo[1971:1968]},
     {slideAddressGen_slideMaskInput_lo[1967:1964]},
     {slideAddressGen_slideMaskInput_lo[1963:1960]},
     {slideAddressGen_slideMaskInput_lo[1959:1956]},
     {slideAddressGen_slideMaskInput_lo[1955:1952]},
     {slideAddressGen_slideMaskInput_lo[1951:1948]},
     {slideAddressGen_slideMaskInput_lo[1947:1944]},
     {slideAddressGen_slideMaskInput_lo[1943:1940]},
     {slideAddressGen_slideMaskInput_lo[1939:1936]},
     {slideAddressGen_slideMaskInput_lo[1935:1932]},
     {slideAddressGen_slideMaskInput_lo[1931:1928]},
     {slideAddressGen_slideMaskInput_lo[1927:1924]},
     {slideAddressGen_slideMaskInput_lo[1923:1920]},
     {slideAddressGen_slideMaskInput_lo[1919:1916]},
     {slideAddressGen_slideMaskInput_lo[1915:1912]},
     {slideAddressGen_slideMaskInput_lo[1911:1908]},
     {slideAddressGen_slideMaskInput_lo[1907:1904]},
     {slideAddressGen_slideMaskInput_lo[1903:1900]},
     {slideAddressGen_slideMaskInput_lo[1899:1896]},
     {slideAddressGen_slideMaskInput_lo[1895:1892]},
     {slideAddressGen_slideMaskInput_lo[1891:1888]},
     {slideAddressGen_slideMaskInput_lo[1887:1884]},
     {slideAddressGen_slideMaskInput_lo[1883:1880]},
     {slideAddressGen_slideMaskInput_lo[1879:1876]},
     {slideAddressGen_slideMaskInput_lo[1875:1872]},
     {slideAddressGen_slideMaskInput_lo[1871:1868]},
     {slideAddressGen_slideMaskInput_lo[1867:1864]},
     {slideAddressGen_slideMaskInput_lo[1863:1860]},
     {slideAddressGen_slideMaskInput_lo[1859:1856]},
     {slideAddressGen_slideMaskInput_lo[1855:1852]},
     {slideAddressGen_slideMaskInput_lo[1851:1848]},
     {slideAddressGen_slideMaskInput_lo[1847:1844]},
     {slideAddressGen_slideMaskInput_lo[1843:1840]},
     {slideAddressGen_slideMaskInput_lo[1839:1836]},
     {slideAddressGen_slideMaskInput_lo[1835:1832]},
     {slideAddressGen_slideMaskInput_lo[1831:1828]},
     {slideAddressGen_slideMaskInput_lo[1827:1824]},
     {slideAddressGen_slideMaskInput_lo[1823:1820]},
     {slideAddressGen_slideMaskInput_lo[1819:1816]},
     {slideAddressGen_slideMaskInput_lo[1815:1812]},
     {slideAddressGen_slideMaskInput_lo[1811:1808]},
     {slideAddressGen_slideMaskInput_lo[1807:1804]},
     {slideAddressGen_slideMaskInput_lo[1803:1800]},
     {slideAddressGen_slideMaskInput_lo[1799:1796]},
     {slideAddressGen_slideMaskInput_lo[1795:1792]},
     {slideAddressGen_slideMaskInput_lo[1791:1788]},
     {slideAddressGen_slideMaskInput_lo[1787:1784]},
     {slideAddressGen_slideMaskInput_lo[1783:1780]},
     {slideAddressGen_slideMaskInput_lo[1779:1776]},
     {slideAddressGen_slideMaskInput_lo[1775:1772]},
     {slideAddressGen_slideMaskInput_lo[1771:1768]},
     {slideAddressGen_slideMaskInput_lo[1767:1764]},
     {slideAddressGen_slideMaskInput_lo[1763:1760]},
     {slideAddressGen_slideMaskInput_lo[1759:1756]},
     {slideAddressGen_slideMaskInput_lo[1755:1752]},
     {slideAddressGen_slideMaskInput_lo[1751:1748]},
     {slideAddressGen_slideMaskInput_lo[1747:1744]},
     {slideAddressGen_slideMaskInput_lo[1743:1740]},
     {slideAddressGen_slideMaskInput_lo[1739:1736]},
     {slideAddressGen_slideMaskInput_lo[1735:1732]},
     {slideAddressGen_slideMaskInput_lo[1731:1728]},
     {slideAddressGen_slideMaskInput_lo[1727:1724]},
     {slideAddressGen_slideMaskInput_lo[1723:1720]},
     {slideAddressGen_slideMaskInput_lo[1719:1716]},
     {slideAddressGen_slideMaskInput_lo[1715:1712]},
     {slideAddressGen_slideMaskInput_lo[1711:1708]},
     {slideAddressGen_slideMaskInput_lo[1707:1704]},
     {slideAddressGen_slideMaskInput_lo[1703:1700]},
     {slideAddressGen_slideMaskInput_lo[1699:1696]},
     {slideAddressGen_slideMaskInput_lo[1695:1692]},
     {slideAddressGen_slideMaskInput_lo[1691:1688]},
     {slideAddressGen_slideMaskInput_lo[1687:1684]},
     {slideAddressGen_slideMaskInput_lo[1683:1680]},
     {slideAddressGen_slideMaskInput_lo[1679:1676]},
     {slideAddressGen_slideMaskInput_lo[1675:1672]},
     {slideAddressGen_slideMaskInput_lo[1671:1668]},
     {slideAddressGen_slideMaskInput_lo[1667:1664]},
     {slideAddressGen_slideMaskInput_lo[1663:1660]},
     {slideAddressGen_slideMaskInput_lo[1659:1656]},
     {slideAddressGen_slideMaskInput_lo[1655:1652]},
     {slideAddressGen_slideMaskInput_lo[1651:1648]},
     {slideAddressGen_slideMaskInput_lo[1647:1644]},
     {slideAddressGen_slideMaskInput_lo[1643:1640]},
     {slideAddressGen_slideMaskInput_lo[1639:1636]},
     {slideAddressGen_slideMaskInput_lo[1635:1632]},
     {slideAddressGen_slideMaskInput_lo[1631:1628]},
     {slideAddressGen_slideMaskInput_lo[1627:1624]},
     {slideAddressGen_slideMaskInput_lo[1623:1620]},
     {slideAddressGen_slideMaskInput_lo[1619:1616]},
     {slideAddressGen_slideMaskInput_lo[1615:1612]},
     {slideAddressGen_slideMaskInput_lo[1611:1608]},
     {slideAddressGen_slideMaskInput_lo[1607:1604]},
     {slideAddressGen_slideMaskInput_lo[1603:1600]},
     {slideAddressGen_slideMaskInput_lo[1599:1596]},
     {slideAddressGen_slideMaskInput_lo[1595:1592]},
     {slideAddressGen_slideMaskInput_lo[1591:1588]},
     {slideAddressGen_slideMaskInput_lo[1587:1584]},
     {slideAddressGen_slideMaskInput_lo[1583:1580]},
     {slideAddressGen_slideMaskInput_lo[1579:1576]},
     {slideAddressGen_slideMaskInput_lo[1575:1572]},
     {slideAddressGen_slideMaskInput_lo[1571:1568]},
     {slideAddressGen_slideMaskInput_lo[1567:1564]},
     {slideAddressGen_slideMaskInput_lo[1563:1560]},
     {slideAddressGen_slideMaskInput_lo[1559:1556]},
     {slideAddressGen_slideMaskInput_lo[1555:1552]},
     {slideAddressGen_slideMaskInput_lo[1551:1548]},
     {slideAddressGen_slideMaskInput_lo[1547:1544]},
     {slideAddressGen_slideMaskInput_lo[1543:1540]},
     {slideAddressGen_slideMaskInput_lo[1539:1536]},
     {slideAddressGen_slideMaskInput_lo[1535:1532]},
     {slideAddressGen_slideMaskInput_lo[1531:1528]},
     {slideAddressGen_slideMaskInput_lo[1527:1524]},
     {slideAddressGen_slideMaskInput_lo[1523:1520]},
     {slideAddressGen_slideMaskInput_lo[1519:1516]},
     {slideAddressGen_slideMaskInput_lo[1515:1512]},
     {slideAddressGen_slideMaskInput_lo[1511:1508]},
     {slideAddressGen_slideMaskInput_lo[1507:1504]},
     {slideAddressGen_slideMaskInput_lo[1503:1500]},
     {slideAddressGen_slideMaskInput_lo[1499:1496]},
     {slideAddressGen_slideMaskInput_lo[1495:1492]},
     {slideAddressGen_slideMaskInput_lo[1491:1488]},
     {slideAddressGen_slideMaskInput_lo[1487:1484]},
     {slideAddressGen_slideMaskInput_lo[1483:1480]},
     {slideAddressGen_slideMaskInput_lo[1479:1476]},
     {slideAddressGen_slideMaskInput_lo[1475:1472]},
     {slideAddressGen_slideMaskInput_lo[1471:1468]},
     {slideAddressGen_slideMaskInput_lo[1467:1464]},
     {slideAddressGen_slideMaskInput_lo[1463:1460]},
     {slideAddressGen_slideMaskInput_lo[1459:1456]},
     {slideAddressGen_slideMaskInput_lo[1455:1452]},
     {slideAddressGen_slideMaskInput_lo[1451:1448]},
     {slideAddressGen_slideMaskInput_lo[1447:1444]},
     {slideAddressGen_slideMaskInput_lo[1443:1440]},
     {slideAddressGen_slideMaskInput_lo[1439:1436]},
     {slideAddressGen_slideMaskInput_lo[1435:1432]},
     {slideAddressGen_slideMaskInput_lo[1431:1428]},
     {slideAddressGen_slideMaskInput_lo[1427:1424]},
     {slideAddressGen_slideMaskInput_lo[1423:1420]},
     {slideAddressGen_slideMaskInput_lo[1419:1416]},
     {slideAddressGen_slideMaskInput_lo[1415:1412]},
     {slideAddressGen_slideMaskInput_lo[1411:1408]},
     {slideAddressGen_slideMaskInput_lo[1407:1404]},
     {slideAddressGen_slideMaskInput_lo[1403:1400]},
     {slideAddressGen_slideMaskInput_lo[1399:1396]},
     {slideAddressGen_slideMaskInput_lo[1395:1392]},
     {slideAddressGen_slideMaskInput_lo[1391:1388]},
     {slideAddressGen_slideMaskInput_lo[1387:1384]},
     {slideAddressGen_slideMaskInput_lo[1383:1380]},
     {slideAddressGen_slideMaskInput_lo[1379:1376]},
     {slideAddressGen_slideMaskInput_lo[1375:1372]},
     {slideAddressGen_slideMaskInput_lo[1371:1368]},
     {slideAddressGen_slideMaskInput_lo[1367:1364]},
     {slideAddressGen_slideMaskInput_lo[1363:1360]},
     {slideAddressGen_slideMaskInput_lo[1359:1356]},
     {slideAddressGen_slideMaskInput_lo[1355:1352]},
     {slideAddressGen_slideMaskInput_lo[1351:1348]},
     {slideAddressGen_slideMaskInput_lo[1347:1344]},
     {slideAddressGen_slideMaskInput_lo[1343:1340]},
     {slideAddressGen_slideMaskInput_lo[1339:1336]},
     {slideAddressGen_slideMaskInput_lo[1335:1332]},
     {slideAddressGen_slideMaskInput_lo[1331:1328]},
     {slideAddressGen_slideMaskInput_lo[1327:1324]},
     {slideAddressGen_slideMaskInput_lo[1323:1320]},
     {slideAddressGen_slideMaskInput_lo[1319:1316]},
     {slideAddressGen_slideMaskInput_lo[1315:1312]},
     {slideAddressGen_slideMaskInput_lo[1311:1308]},
     {slideAddressGen_slideMaskInput_lo[1307:1304]},
     {slideAddressGen_slideMaskInput_lo[1303:1300]},
     {slideAddressGen_slideMaskInput_lo[1299:1296]},
     {slideAddressGen_slideMaskInput_lo[1295:1292]},
     {slideAddressGen_slideMaskInput_lo[1291:1288]},
     {slideAddressGen_slideMaskInput_lo[1287:1284]},
     {slideAddressGen_slideMaskInput_lo[1283:1280]},
     {slideAddressGen_slideMaskInput_lo[1279:1276]},
     {slideAddressGen_slideMaskInput_lo[1275:1272]},
     {slideAddressGen_slideMaskInput_lo[1271:1268]},
     {slideAddressGen_slideMaskInput_lo[1267:1264]},
     {slideAddressGen_slideMaskInput_lo[1263:1260]},
     {slideAddressGen_slideMaskInput_lo[1259:1256]},
     {slideAddressGen_slideMaskInput_lo[1255:1252]},
     {slideAddressGen_slideMaskInput_lo[1251:1248]},
     {slideAddressGen_slideMaskInput_lo[1247:1244]},
     {slideAddressGen_slideMaskInput_lo[1243:1240]},
     {slideAddressGen_slideMaskInput_lo[1239:1236]},
     {slideAddressGen_slideMaskInput_lo[1235:1232]},
     {slideAddressGen_slideMaskInput_lo[1231:1228]},
     {slideAddressGen_slideMaskInput_lo[1227:1224]},
     {slideAddressGen_slideMaskInput_lo[1223:1220]},
     {slideAddressGen_slideMaskInput_lo[1219:1216]},
     {slideAddressGen_slideMaskInput_lo[1215:1212]},
     {slideAddressGen_slideMaskInput_lo[1211:1208]},
     {slideAddressGen_slideMaskInput_lo[1207:1204]},
     {slideAddressGen_slideMaskInput_lo[1203:1200]},
     {slideAddressGen_slideMaskInput_lo[1199:1196]},
     {slideAddressGen_slideMaskInput_lo[1195:1192]},
     {slideAddressGen_slideMaskInput_lo[1191:1188]},
     {slideAddressGen_slideMaskInput_lo[1187:1184]},
     {slideAddressGen_slideMaskInput_lo[1183:1180]},
     {slideAddressGen_slideMaskInput_lo[1179:1176]},
     {slideAddressGen_slideMaskInput_lo[1175:1172]},
     {slideAddressGen_slideMaskInput_lo[1171:1168]},
     {slideAddressGen_slideMaskInput_lo[1167:1164]},
     {slideAddressGen_slideMaskInput_lo[1163:1160]},
     {slideAddressGen_slideMaskInput_lo[1159:1156]},
     {slideAddressGen_slideMaskInput_lo[1155:1152]},
     {slideAddressGen_slideMaskInput_lo[1151:1148]},
     {slideAddressGen_slideMaskInput_lo[1147:1144]},
     {slideAddressGen_slideMaskInput_lo[1143:1140]},
     {slideAddressGen_slideMaskInput_lo[1139:1136]},
     {slideAddressGen_slideMaskInput_lo[1135:1132]},
     {slideAddressGen_slideMaskInput_lo[1131:1128]},
     {slideAddressGen_slideMaskInput_lo[1127:1124]},
     {slideAddressGen_slideMaskInput_lo[1123:1120]},
     {slideAddressGen_slideMaskInput_lo[1119:1116]},
     {slideAddressGen_slideMaskInput_lo[1115:1112]},
     {slideAddressGen_slideMaskInput_lo[1111:1108]},
     {slideAddressGen_slideMaskInput_lo[1107:1104]},
     {slideAddressGen_slideMaskInput_lo[1103:1100]},
     {slideAddressGen_slideMaskInput_lo[1099:1096]},
     {slideAddressGen_slideMaskInput_lo[1095:1092]},
     {slideAddressGen_slideMaskInput_lo[1091:1088]},
     {slideAddressGen_slideMaskInput_lo[1087:1084]},
     {slideAddressGen_slideMaskInput_lo[1083:1080]},
     {slideAddressGen_slideMaskInput_lo[1079:1076]},
     {slideAddressGen_slideMaskInput_lo[1075:1072]},
     {slideAddressGen_slideMaskInput_lo[1071:1068]},
     {slideAddressGen_slideMaskInput_lo[1067:1064]},
     {slideAddressGen_slideMaskInput_lo[1063:1060]},
     {slideAddressGen_slideMaskInput_lo[1059:1056]},
     {slideAddressGen_slideMaskInput_lo[1055:1052]},
     {slideAddressGen_slideMaskInput_lo[1051:1048]},
     {slideAddressGen_slideMaskInput_lo[1047:1044]},
     {slideAddressGen_slideMaskInput_lo[1043:1040]},
     {slideAddressGen_slideMaskInput_lo[1039:1036]},
     {slideAddressGen_slideMaskInput_lo[1035:1032]},
     {slideAddressGen_slideMaskInput_lo[1031:1028]},
     {slideAddressGen_slideMaskInput_lo[1027:1024]},
     {slideAddressGen_slideMaskInput_lo[1023:1020]},
     {slideAddressGen_slideMaskInput_lo[1019:1016]},
     {slideAddressGen_slideMaskInput_lo[1015:1012]},
     {slideAddressGen_slideMaskInput_lo[1011:1008]},
     {slideAddressGen_slideMaskInput_lo[1007:1004]},
     {slideAddressGen_slideMaskInput_lo[1003:1000]},
     {slideAddressGen_slideMaskInput_lo[999:996]},
     {slideAddressGen_slideMaskInput_lo[995:992]},
     {slideAddressGen_slideMaskInput_lo[991:988]},
     {slideAddressGen_slideMaskInput_lo[987:984]},
     {slideAddressGen_slideMaskInput_lo[983:980]},
     {slideAddressGen_slideMaskInput_lo[979:976]},
     {slideAddressGen_slideMaskInput_lo[975:972]},
     {slideAddressGen_slideMaskInput_lo[971:968]},
     {slideAddressGen_slideMaskInput_lo[967:964]},
     {slideAddressGen_slideMaskInput_lo[963:960]},
     {slideAddressGen_slideMaskInput_lo[959:956]},
     {slideAddressGen_slideMaskInput_lo[955:952]},
     {slideAddressGen_slideMaskInput_lo[951:948]},
     {slideAddressGen_slideMaskInput_lo[947:944]},
     {slideAddressGen_slideMaskInput_lo[943:940]},
     {slideAddressGen_slideMaskInput_lo[939:936]},
     {slideAddressGen_slideMaskInput_lo[935:932]},
     {slideAddressGen_slideMaskInput_lo[931:928]},
     {slideAddressGen_slideMaskInput_lo[927:924]},
     {slideAddressGen_slideMaskInput_lo[923:920]},
     {slideAddressGen_slideMaskInput_lo[919:916]},
     {slideAddressGen_slideMaskInput_lo[915:912]},
     {slideAddressGen_slideMaskInput_lo[911:908]},
     {slideAddressGen_slideMaskInput_lo[907:904]},
     {slideAddressGen_slideMaskInput_lo[903:900]},
     {slideAddressGen_slideMaskInput_lo[899:896]},
     {slideAddressGen_slideMaskInput_lo[895:892]},
     {slideAddressGen_slideMaskInput_lo[891:888]},
     {slideAddressGen_slideMaskInput_lo[887:884]},
     {slideAddressGen_slideMaskInput_lo[883:880]},
     {slideAddressGen_slideMaskInput_lo[879:876]},
     {slideAddressGen_slideMaskInput_lo[875:872]},
     {slideAddressGen_slideMaskInput_lo[871:868]},
     {slideAddressGen_slideMaskInput_lo[867:864]},
     {slideAddressGen_slideMaskInput_lo[863:860]},
     {slideAddressGen_slideMaskInput_lo[859:856]},
     {slideAddressGen_slideMaskInput_lo[855:852]},
     {slideAddressGen_slideMaskInput_lo[851:848]},
     {slideAddressGen_slideMaskInput_lo[847:844]},
     {slideAddressGen_slideMaskInput_lo[843:840]},
     {slideAddressGen_slideMaskInput_lo[839:836]},
     {slideAddressGen_slideMaskInput_lo[835:832]},
     {slideAddressGen_slideMaskInput_lo[831:828]},
     {slideAddressGen_slideMaskInput_lo[827:824]},
     {slideAddressGen_slideMaskInput_lo[823:820]},
     {slideAddressGen_slideMaskInput_lo[819:816]},
     {slideAddressGen_slideMaskInput_lo[815:812]},
     {slideAddressGen_slideMaskInput_lo[811:808]},
     {slideAddressGen_slideMaskInput_lo[807:804]},
     {slideAddressGen_slideMaskInput_lo[803:800]},
     {slideAddressGen_slideMaskInput_lo[799:796]},
     {slideAddressGen_slideMaskInput_lo[795:792]},
     {slideAddressGen_slideMaskInput_lo[791:788]},
     {slideAddressGen_slideMaskInput_lo[787:784]},
     {slideAddressGen_slideMaskInput_lo[783:780]},
     {slideAddressGen_slideMaskInput_lo[779:776]},
     {slideAddressGen_slideMaskInput_lo[775:772]},
     {slideAddressGen_slideMaskInput_lo[771:768]},
     {slideAddressGen_slideMaskInput_lo[767:764]},
     {slideAddressGen_slideMaskInput_lo[763:760]},
     {slideAddressGen_slideMaskInput_lo[759:756]},
     {slideAddressGen_slideMaskInput_lo[755:752]},
     {slideAddressGen_slideMaskInput_lo[751:748]},
     {slideAddressGen_slideMaskInput_lo[747:744]},
     {slideAddressGen_slideMaskInput_lo[743:740]},
     {slideAddressGen_slideMaskInput_lo[739:736]},
     {slideAddressGen_slideMaskInput_lo[735:732]},
     {slideAddressGen_slideMaskInput_lo[731:728]},
     {slideAddressGen_slideMaskInput_lo[727:724]},
     {slideAddressGen_slideMaskInput_lo[723:720]},
     {slideAddressGen_slideMaskInput_lo[719:716]},
     {slideAddressGen_slideMaskInput_lo[715:712]},
     {slideAddressGen_slideMaskInput_lo[711:708]},
     {slideAddressGen_slideMaskInput_lo[707:704]},
     {slideAddressGen_slideMaskInput_lo[703:700]},
     {slideAddressGen_slideMaskInput_lo[699:696]},
     {slideAddressGen_slideMaskInput_lo[695:692]},
     {slideAddressGen_slideMaskInput_lo[691:688]},
     {slideAddressGen_slideMaskInput_lo[687:684]},
     {slideAddressGen_slideMaskInput_lo[683:680]},
     {slideAddressGen_slideMaskInput_lo[679:676]},
     {slideAddressGen_slideMaskInput_lo[675:672]},
     {slideAddressGen_slideMaskInput_lo[671:668]},
     {slideAddressGen_slideMaskInput_lo[667:664]},
     {slideAddressGen_slideMaskInput_lo[663:660]},
     {slideAddressGen_slideMaskInput_lo[659:656]},
     {slideAddressGen_slideMaskInput_lo[655:652]},
     {slideAddressGen_slideMaskInput_lo[651:648]},
     {slideAddressGen_slideMaskInput_lo[647:644]},
     {slideAddressGen_slideMaskInput_lo[643:640]},
     {slideAddressGen_slideMaskInput_lo[639:636]},
     {slideAddressGen_slideMaskInput_lo[635:632]},
     {slideAddressGen_slideMaskInput_lo[631:628]},
     {slideAddressGen_slideMaskInput_lo[627:624]},
     {slideAddressGen_slideMaskInput_lo[623:620]},
     {slideAddressGen_slideMaskInput_lo[619:616]},
     {slideAddressGen_slideMaskInput_lo[615:612]},
     {slideAddressGen_slideMaskInput_lo[611:608]},
     {slideAddressGen_slideMaskInput_lo[607:604]},
     {slideAddressGen_slideMaskInput_lo[603:600]},
     {slideAddressGen_slideMaskInput_lo[599:596]},
     {slideAddressGen_slideMaskInput_lo[595:592]},
     {slideAddressGen_slideMaskInput_lo[591:588]},
     {slideAddressGen_slideMaskInput_lo[587:584]},
     {slideAddressGen_slideMaskInput_lo[583:580]},
     {slideAddressGen_slideMaskInput_lo[579:576]},
     {slideAddressGen_slideMaskInput_lo[575:572]},
     {slideAddressGen_slideMaskInput_lo[571:568]},
     {slideAddressGen_slideMaskInput_lo[567:564]},
     {slideAddressGen_slideMaskInput_lo[563:560]},
     {slideAddressGen_slideMaskInput_lo[559:556]},
     {slideAddressGen_slideMaskInput_lo[555:552]},
     {slideAddressGen_slideMaskInput_lo[551:548]},
     {slideAddressGen_slideMaskInput_lo[547:544]},
     {slideAddressGen_slideMaskInput_lo[543:540]},
     {slideAddressGen_slideMaskInput_lo[539:536]},
     {slideAddressGen_slideMaskInput_lo[535:532]},
     {slideAddressGen_slideMaskInput_lo[531:528]},
     {slideAddressGen_slideMaskInput_lo[527:524]},
     {slideAddressGen_slideMaskInput_lo[523:520]},
     {slideAddressGen_slideMaskInput_lo[519:516]},
     {slideAddressGen_slideMaskInput_lo[515:512]},
     {slideAddressGen_slideMaskInput_lo[511:508]},
     {slideAddressGen_slideMaskInput_lo[507:504]},
     {slideAddressGen_slideMaskInput_lo[503:500]},
     {slideAddressGen_slideMaskInput_lo[499:496]},
     {slideAddressGen_slideMaskInput_lo[495:492]},
     {slideAddressGen_slideMaskInput_lo[491:488]},
     {slideAddressGen_slideMaskInput_lo[487:484]},
     {slideAddressGen_slideMaskInput_lo[483:480]},
     {slideAddressGen_slideMaskInput_lo[479:476]},
     {slideAddressGen_slideMaskInput_lo[475:472]},
     {slideAddressGen_slideMaskInput_lo[471:468]},
     {slideAddressGen_slideMaskInput_lo[467:464]},
     {slideAddressGen_slideMaskInput_lo[463:460]},
     {slideAddressGen_slideMaskInput_lo[459:456]},
     {slideAddressGen_slideMaskInput_lo[455:452]},
     {slideAddressGen_slideMaskInput_lo[451:448]},
     {slideAddressGen_slideMaskInput_lo[447:444]},
     {slideAddressGen_slideMaskInput_lo[443:440]},
     {slideAddressGen_slideMaskInput_lo[439:436]},
     {slideAddressGen_slideMaskInput_lo[435:432]},
     {slideAddressGen_slideMaskInput_lo[431:428]},
     {slideAddressGen_slideMaskInput_lo[427:424]},
     {slideAddressGen_slideMaskInput_lo[423:420]},
     {slideAddressGen_slideMaskInput_lo[419:416]},
     {slideAddressGen_slideMaskInput_lo[415:412]},
     {slideAddressGen_slideMaskInput_lo[411:408]},
     {slideAddressGen_slideMaskInput_lo[407:404]},
     {slideAddressGen_slideMaskInput_lo[403:400]},
     {slideAddressGen_slideMaskInput_lo[399:396]},
     {slideAddressGen_slideMaskInput_lo[395:392]},
     {slideAddressGen_slideMaskInput_lo[391:388]},
     {slideAddressGen_slideMaskInput_lo[387:384]},
     {slideAddressGen_slideMaskInput_lo[383:380]},
     {slideAddressGen_slideMaskInput_lo[379:376]},
     {slideAddressGen_slideMaskInput_lo[375:372]},
     {slideAddressGen_slideMaskInput_lo[371:368]},
     {slideAddressGen_slideMaskInput_lo[367:364]},
     {slideAddressGen_slideMaskInput_lo[363:360]},
     {slideAddressGen_slideMaskInput_lo[359:356]},
     {slideAddressGen_slideMaskInput_lo[355:352]},
     {slideAddressGen_slideMaskInput_lo[351:348]},
     {slideAddressGen_slideMaskInput_lo[347:344]},
     {slideAddressGen_slideMaskInput_lo[343:340]},
     {slideAddressGen_slideMaskInput_lo[339:336]},
     {slideAddressGen_slideMaskInput_lo[335:332]},
     {slideAddressGen_slideMaskInput_lo[331:328]},
     {slideAddressGen_slideMaskInput_lo[327:324]},
     {slideAddressGen_slideMaskInput_lo[323:320]},
     {slideAddressGen_slideMaskInput_lo[319:316]},
     {slideAddressGen_slideMaskInput_lo[315:312]},
     {slideAddressGen_slideMaskInput_lo[311:308]},
     {slideAddressGen_slideMaskInput_lo[307:304]},
     {slideAddressGen_slideMaskInput_lo[303:300]},
     {slideAddressGen_slideMaskInput_lo[299:296]},
     {slideAddressGen_slideMaskInput_lo[295:292]},
     {slideAddressGen_slideMaskInput_lo[291:288]},
     {slideAddressGen_slideMaskInput_lo[287:284]},
     {slideAddressGen_slideMaskInput_lo[283:280]},
     {slideAddressGen_slideMaskInput_lo[279:276]},
     {slideAddressGen_slideMaskInput_lo[275:272]},
     {slideAddressGen_slideMaskInput_lo[271:268]},
     {slideAddressGen_slideMaskInput_lo[267:264]},
     {slideAddressGen_slideMaskInput_lo[263:260]},
     {slideAddressGen_slideMaskInput_lo[259:256]},
     {slideAddressGen_slideMaskInput_lo[255:252]},
     {slideAddressGen_slideMaskInput_lo[251:248]},
     {slideAddressGen_slideMaskInput_lo[247:244]},
     {slideAddressGen_slideMaskInput_lo[243:240]},
     {slideAddressGen_slideMaskInput_lo[239:236]},
     {slideAddressGen_slideMaskInput_lo[235:232]},
     {slideAddressGen_slideMaskInput_lo[231:228]},
     {slideAddressGen_slideMaskInput_lo[227:224]},
     {slideAddressGen_slideMaskInput_lo[223:220]},
     {slideAddressGen_slideMaskInput_lo[219:216]},
     {slideAddressGen_slideMaskInput_lo[215:212]},
     {slideAddressGen_slideMaskInput_lo[211:208]},
     {slideAddressGen_slideMaskInput_lo[207:204]},
     {slideAddressGen_slideMaskInput_lo[203:200]},
     {slideAddressGen_slideMaskInput_lo[199:196]},
     {slideAddressGen_slideMaskInput_lo[195:192]},
     {slideAddressGen_slideMaskInput_lo[191:188]},
     {slideAddressGen_slideMaskInput_lo[187:184]},
     {slideAddressGen_slideMaskInput_lo[183:180]},
     {slideAddressGen_slideMaskInput_lo[179:176]},
     {slideAddressGen_slideMaskInput_lo[175:172]},
     {slideAddressGen_slideMaskInput_lo[171:168]},
     {slideAddressGen_slideMaskInput_lo[167:164]},
     {slideAddressGen_slideMaskInput_lo[163:160]},
     {slideAddressGen_slideMaskInput_lo[159:156]},
     {slideAddressGen_slideMaskInput_lo[155:152]},
     {slideAddressGen_slideMaskInput_lo[151:148]},
     {slideAddressGen_slideMaskInput_lo[147:144]},
     {slideAddressGen_slideMaskInput_lo[143:140]},
     {slideAddressGen_slideMaskInput_lo[139:136]},
     {slideAddressGen_slideMaskInput_lo[135:132]},
     {slideAddressGen_slideMaskInput_lo[131:128]},
     {slideAddressGen_slideMaskInput_lo[127:124]},
     {slideAddressGen_slideMaskInput_lo[123:120]},
     {slideAddressGen_slideMaskInput_lo[119:116]},
     {slideAddressGen_slideMaskInput_lo[115:112]},
     {slideAddressGen_slideMaskInput_lo[111:108]},
     {slideAddressGen_slideMaskInput_lo[107:104]},
     {slideAddressGen_slideMaskInput_lo[103:100]},
     {slideAddressGen_slideMaskInput_lo[99:96]},
     {slideAddressGen_slideMaskInput_lo[95:92]},
     {slideAddressGen_slideMaskInput_lo[91:88]},
     {slideAddressGen_slideMaskInput_lo[87:84]},
     {slideAddressGen_slideMaskInput_lo[83:80]},
     {slideAddressGen_slideMaskInput_lo[79:76]},
     {slideAddressGen_slideMaskInput_lo[75:72]},
     {slideAddressGen_slideMaskInput_lo[71:68]},
     {slideAddressGen_slideMaskInput_lo[67:64]},
     {slideAddressGen_slideMaskInput_lo[63:60]},
     {slideAddressGen_slideMaskInput_lo[59:56]},
     {slideAddressGen_slideMaskInput_lo[55:52]},
     {slideAddressGen_slideMaskInput_lo[51:48]},
     {slideAddressGen_slideMaskInput_lo[47:44]},
     {slideAddressGen_slideMaskInput_lo[43:40]},
     {slideAddressGen_slideMaskInput_lo[39:36]},
     {slideAddressGen_slideMaskInput_lo[35:32]},
     {slideAddressGen_slideMaskInput_lo[31:28]},
     {slideAddressGen_slideMaskInput_lo[27:24]},
     {slideAddressGen_slideMaskInput_lo[23:20]},
     {slideAddressGen_slideMaskInput_lo[19:16]},
     {slideAddressGen_slideMaskInput_lo[15:12]},
     {slideAddressGen_slideMaskInput_lo[11:8]},
     {slideAddressGen_slideMaskInput_lo[7:4]},
     {slideAddressGen_slideMaskInput_lo[3:0]}};
  wire               lastExecuteGroupDeq;
  wire               viotaCounterAdd;
  wire               groupCounterAdd = noSource ? viotaCounterAdd : lastExecuteGroupDeq;
  wire [3:0]         groupDataNeed = lastGroup ? lastGroupDataNeed : 4'hF;
  reg  [1:0]         executeIndex;
  reg  [3:0]         readIssueStageState_groupReadState;
  reg  [3:0]         readIssueStageState_needRead;
  wire [3:0]         readWaitQueue_enq_bits_needRead = readIssueStageState_needRead;
  reg  [3:0]         readIssueStageState_elementValid;
  wire [3:0]         readWaitQueue_enq_bits_sourceValid = readIssueStageState_elementValid;
  reg  [3:0]         readIssueStageState_replaceVs1;
  wire [3:0]         readWaitQueue_enq_bits_replaceVs1 = readIssueStageState_replaceVs1;
  reg  [23:0]        readIssueStageState_readOffset;
  reg  [1:0]         readIssueStageState_accessLane_0;
  reg  [1:0]         readIssueStageState_accessLane_1;
  wire [1:0]         selectExecuteReq_1_bits_readLane = readIssueStageState_accessLane_1;
  reg  [1:0]         readIssueStageState_accessLane_2;
  wire [1:0]         selectExecuteReq_2_bits_readLane = readIssueStageState_accessLane_2;
  reg  [1:0]         readIssueStageState_accessLane_3;
  wire [1:0]         selectExecuteReq_3_bits_readLane = readIssueStageState_accessLane_3;
  reg  [2:0]         readIssueStageState_vsGrowth_0;
  reg  [2:0]         readIssueStageState_vsGrowth_1;
  reg  [2:0]         readIssueStageState_vsGrowth_2;
  reg  [2:0]         readIssueStageState_vsGrowth_3;
  reg  [11:0]        readIssueStageState_executeGroup;
  wire [11:0]        readWaitQueue_enq_bits_executeGroup = readIssueStageState_executeGroup;
  reg  [7:0]         readIssueStageState_readDataOffset;
  reg                readIssueStageState_last;
  wire               readWaitQueue_enq_bits_last = readIssueStageState_last;
  reg                readIssueStageValid;
  wire [2:0]         accessCountQueue_enq_bits_0 = accessCountEnq_0;
  wire [2:0]         accessCountQueue_enq_bits_1 = accessCountEnq_1;
  wire [2:0]         accessCountQueue_enq_bits_2 = accessCountEnq_2;
  wire [2:0]         accessCountQueue_enq_bits_3 = accessCountEnq_3;
  wire               readIssueStageEnq;
  wire               accessCountQueue_deq_valid;
  assign accessCountQueue_deq_valid = ~_accessCountQueue_fifo_empty;
  wire [2:0]         accessCountQueue_dataOut_0;
  wire [2:0]         accessCountQueue_dataOut_1;
  wire [2:0]         accessCountQueue_dataOut_2;
  wire [2:0]         accessCountQueue_dataOut_3;
  wire [5:0]         accessCountQueue_dataIn_lo = {accessCountQueue_enq_bits_1, accessCountQueue_enq_bits_0};
  wire [5:0]         accessCountQueue_dataIn_hi = {accessCountQueue_enq_bits_3, accessCountQueue_enq_bits_2};
  wire [11:0]        accessCountQueue_dataIn = {accessCountQueue_dataIn_hi, accessCountQueue_dataIn_lo};
  assign accessCountQueue_dataOut_0 = _accessCountQueue_fifo_data_out[2:0];
  assign accessCountQueue_dataOut_1 = _accessCountQueue_fifo_data_out[5:3];
  assign accessCountQueue_dataOut_2 = _accessCountQueue_fifo_data_out[8:6];
  assign accessCountQueue_dataOut_3 = _accessCountQueue_fifo_data_out[11:9];
  wire [2:0]         accessCountQueue_deq_bits_0 = accessCountQueue_dataOut_0;
  wire [2:0]         accessCountQueue_deq_bits_1 = accessCountQueue_dataOut_1;
  wire [2:0]         accessCountQueue_deq_bits_2 = accessCountQueue_dataOut_2;
  wire [2:0]         accessCountQueue_deq_bits_3 = accessCountQueue_dataOut_3;
  wire               accessCountQueue_enq_ready = ~_accessCountQueue_fifo_full;
  wire               accessCountQueue_enq_valid;
  wire               accessCountQueue_deq_ready;
  wire [11:0]        _extendGroupCount_T_1 = {requestCounter, executeIndex};
  wire [11:0]        _executeGroup_T_8 = executeIndexGrowth[0] ? _extendGroupCount_T_1 : 12'h0;
  wire [10:0]        _GEN_141 = _executeGroup_T_8[10:0] | (executeIndexGrowth[1] ? {requestCounter, executeIndex[1]} : 11'h0);
  wire [11:0]        executeGroup = {_executeGroup_T_8[11], _GEN_141[10], _GEN_141[9:0] | (executeIndexGrowth[2] ? requestCounter : 10'h0)};
  wire               vlMisAlign;
  assign vlMisAlign = |(instReg_vl[1:0]);
  wire [11:0]        lastexecuteGroup = instReg_vl[13:2] - {11'h0, ~vlMisAlign};
  wire               isVlBoundary = executeGroup == lastexecuteGroup;
  wire               validExecuteGroup = executeGroup <= lastexecuteGroup;
  wire [3:0]         _maskSplit_vlBoundaryCorrection_T_37 = 4'h1 << instReg_vl[1:0];
  wire [3:0]         _vlBoundaryCorrection_T_5 = _maskSplit_vlBoundaryCorrection_T_37 | {_maskSplit_vlBoundaryCorrection_T_37[2:0], 1'h0};
  wire [3:0]         vlBoundaryCorrection = ~({4{vlMisAlign & isVlBoundary}} & (_vlBoundaryCorrection_T_5 | {_vlBoundaryCorrection_T_5[1:0], 2'h0})) & {4{validExecuteGroup}};
  wire [127:0]       selectReadStageMask_lo_lo_lo_lo_lo_lo = {selectReadStageMask_lo_lo_lo_lo_lo_lo_hi, selectReadStageMask_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]       selectReadStageMask_lo_lo_lo_lo_lo_hi = {selectReadStageMask_lo_lo_lo_lo_lo_hi_hi, selectReadStageMask_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]       selectReadStageMask_lo_lo_lo_lo_lo = {selectReadStageMask_lo_lo_lo_lo_lo_hi, selectReadStageMask_lo_lo_lo_lo_lo_lo};
  wire [127:0]       selectReadStageMask_lo_lo_lo_lo_hi_lo = {selectReadStageMask_lo_lo_lo_lo_hi_lo_hi, selectReadStageMask_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]       selectReadStageMask_lo_lo_lo_lo_hi_hi = {selectReadStageMask_lo_lo_lo_lo_hi_hi_hi, selectReadStageMask_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]       selectReadStageMask_lo_lo_lo_lo_hi = {selectReadStageMask_lo_lo_lo_lo_hi_hi, selectReadStageMask_lo_lo_lo_lo_hi_lo};
  wire [511:0]       selectReadStageMask_lo_lo_lo_lo = {selectReadStageMask_lo_lo_lo_lo_hi, selectReadStageMask_lo_lo_lo_lo_lo};
  wire [127:0]       selectReadStageMask_lo_lo_lo_hi_lo_lo = {selectReadStageMask_lo_lo_lo_hi_lo_lo_hi, selectReadStageMask_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]       selectReadStageMask_lo_lo_lo_hi_lo_hi = {selectReadStageMask_lo_lo_lo_hi_lo_hi_hi, selectReadStageMask_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]       selectReadStageMask_lo_lo_lo_hi_lo = {selectReadStageMask_lo_lo_lo_hi_lo_hi, selectReadStageMask_lo_lo_lo_hi_lo_lo};
  wire [127:0]       selectReadStageMask_lo_lo_lo_hi_hi_lo = {selectReadStageMask_lo_lo_lo_hi_hi_lo_hi, selectReadStageMask_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]       selectReadStageMask_lo_lo_lo_hi_hi_hi = {selectReadStageMask_lo_lo_lo_hi_hi_hi_hi, selectReadStageMask_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]       selectReadStageMask_lo_lo_lo_hi_hi = {selectReadStageMask_lo_lo_lo_hi_hi_hi, selectReadStageMask_lo_lo_lo_hi_hi_lo};
  wire [511:0]       selectReadStageMask_lo_lo_lo_hi = {selectReadStageMask_lo_lo_lo_hi_hi, selectReadStageMask_lo_lo_lo_hi_lo};
  wire [1023:0]      selectReadStageMask_lo_lo_lo = {selectReadStageMask_lo_lo_lo_hi, selectReadStageMask_lo_lo_lo_lo};
  wire [127:0]       selectReadStageMask_lo_lo_hi_lo_lo_lo = {selectReadStageMask_lo_lo_hi_lo_lo_lo_hi, selectReadStageMask_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]       selectReadStageMask_lo_lo_hi_lo_lo_hi = {selectReadStageMask_lo_lo_hi_lo_lo_hi_hi, selectReadStageMask_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]       selectReadStageMask_lo_lo_hi_lo_lo = {selectReadStageMask_lo_lo_hi_lo_lo_hi, selectReadStageMask_lo_lo_hi_lo_lo_lo};
  wire [127:0]       selectReadStageMask_lo_lo_hi_lo_hi_lo = {selectReadStageMask_lo_lo_hi_lo_hi_lo_hi, selectReadStageMask_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]       selectReadStageMask_lo_lo_hi_lo_hi_hi = {selectReadStageMask_lo_lo_hi_lo_hi_hi_hi, selectReadStageMask_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]       selectReadStageMask_lo_lo_hi_lo_hi = {selectReadStageMask_lo_lo_hi_lo_hi_hi, selectReadStageMask_lo_lo_hi_lo_hi_lo};
  wire [511:0]       selectReadStageMask_lo_lo_hi_lo = {selectReadStageMask_lo_lo_hi_lo_hi, selectReadStageMask_lo_lo_hi_lo_lo};
  wire [127:0]       selectReadStageMask_lo_lo_hi_hi_lo_lo = {selectReadStageMask_lo_lo_hi_hi_lo_lo_hi, selectReadStageMask_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]       selectReadStageMask_lo_lo_hi_hi_lo_hi = {selectReadStageMask_lo_lo_hi_hi_lo_hi_hi, selectReadStageMask_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]       selectReadStageMask_lo_lo_hi_hi_lo = {selectReadStageMask_lo_lo_hi_hi_lo_hi, selectReadStageMask_lo_lo_hi_hi_lo_lo};
  wire [127:0]       selectReadStageMask_lo_lo_hi_hi_hi_lo = {selectReadStageMask_lo_lo_hi_hi_hi_lo_hi, selectReadStageMask_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]       selectReadStageMask_lo_lo_hi_hi_hi_hi = {selectReadStageMask_lo_lo_hi_hi_hi_hi_hi, selectReadStageMask_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]       selectReadStageMask_lo_lo_hi_hi_hi = {selectReadStageMask_lo_lo_hi_hi_hi_hi, selectReadStageMask_lo_lo_hi_hi_hi_lo};
  wire [511:0]       selectReadStageMask_lo_lo_hi_hi = {selectReadStageMask_lo_lo_hi_hi_hi, selectReadStageMask_lo_lo_hi_hi_lo};
  wire [1023:0]      selectReadStageMask_lo_lo_hi = {selectReadStageMask_lo_lo_hi_hi, selectReadStageMask_lo_lo_hi_lo};
  wire [2047:0]      selectReadStageMask_lo_lo = {selectReadStageMask_lo_lo_hi, selectReadStageMask_lo_lo_lo};
  wire [127:0]       selectReadStageMask_lo_hi_lo_lo_lo_lo = {selectReadStageMask_lo_hi_lo_lo_lo_lo_hi, selectReadStageMask_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]       selectReadStageMask_lo_hi_lo_lo_lo_hi = {selectReadStageMask_lo_hi_lo_lo_lo_hi_hi, selectReadStageMask_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]       selectReadStageMask_lo_hi_lo_lo_lo = {selectReadStageMask_lo_hi_lo_lo_lo_hi, selectReadStageMask_lo_hi_lo_lo_lo_lo};
  wire [127:0]       selectReadStageMask_lo_hi_lo_lo_hi_lo = {selectReadStageMask_lo_hi_lo_lo_hi_lo_hi, selectReadStageMask_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]       selectReadStageMask_lo_hi_lo_lo_hi_hi = {selectReadStageMask_lo_hi_lo_lo_hi_hi_hi, selectReadStageMask_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]       selectReadStageMask_lo_hi_lo_lo_hi = {selectReadStageMask_lo_hi_lo_lo_hi_hi, selectReadStageMask_lo_hi_lo_lo_hi_lo};
  wire [511:0]       selectReadStageMask_lo_hi_lo_lo = {selectReadStageMask_lo_hi_lo_lo_hi, selectReadStageMask_lo_hi_lo_lo_lo};
  wire [127:0]       selectReadStageMask_lo_hi_lo_hi_lo_lo = {selectReadStageMask_lo_hi_lo_hi_lo_lo_hi, selectReadStageMask_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]       selectReadStageMask_lo_hi_lo_hi_lo_hi = {selectReadStageMask_lo_hi_lo_hi_lo_hi_hi, selectReadStageMask_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]       selectReadStageMask_lo_hi_lo_hi_lo = {selectReadStageMask_lo_hi_lo_hi_lo_hi, selectReadStageMask_lo_hi_lo_hi_lo_lo};
  wire [127:0]       selectReadStageMask_lo_hi_lo_hi_hi_lo = {selectReadStageMask_lo_hi_lo_hi_hi_lo_hi, selectReadStageMask_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]       selectReadStageMask_lo_hi_lo_hi_hi_hi = {selectReadStageMask_lo_hi_lo_hi_hi_hi_hi, selectReadStageMask_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]       selectReadStageMask_lo_hi_lo_hi_hi = {selectReadStageMask_lo_hi_lo_hi_hi_hi, selectReadStageMask_lo_hi_lo_hi_hi_lo};
  wire [511:0]       selectReadStageMask_lo_hi_lo_hi = {selectReadStageMask_lo_hi_lo_hi_hi, selectReadStageMask_lo_hi_lo_hi_lo};
  wire [1023:0]      selectReadStageMask_lo_hi_lo = {selectReadStageMask_lo_hi_lo_hi, selectReadStageMask_lo_hi_lo_lo};
  wire [127:0]       selectReadStageMask_lo_hi_hi_lo_lo_lo = {selectReadStageMask_lo_hi_hi_lo_lo_lo_hi, selectReadStageMask_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]       selectReadStageMask_lo_hi_hi_lo_lo_hi = {selectReadStageMask_lo_hi_hi_lo_lo_hi_hi, selectReadStageMask_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]       selectReadStageMask_lo_hi_hi_lo_lo = {selectReadStageMask_lo_hi_hi_lo_lo_hi, selectReadStageMask_lo_hi_hi_lo_lo_lo};
  wire [127:0]       selectReadStageMask_lo_hi_hi_lo_hi_lo = {selectReadStageMask_lo_hi_hi_lo_hi_lo_hi, selectReadStageMask_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]       selectReadStageMask_lo_hi_hi_lo_hi_hi = {selectReadStageMask_lo_hi_hi_lo_hi_hi_hi, selectReadStageMask_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]       selectReadStageMask_lo_hi_hi_lo_hi = {selectReadStageMask_lo_hi_hi_lo_hi_hi, selectReadStageMask_lo_hi_hi_lo_hi_lo};
  wire [511:0]       selectReadStageMask_lo_hi_hi_lo = {selectReadStageMask_lo_hi_hi_lo_hi, selectReadStageMask_lo_hi_hi_lo_lo};
  wire [127:0]       selectReadStageMask_lo_hi_hi_hi_lo_lo = {selectReadStageMask_lo_hi_hi_hi_lo_lo_hi, selectReadStageMask_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]       selectReadStageMask_lo_hi_hi_hi_lo_hi = {selectReadStageMask_lo_hi_hi_hi_lo_hi_hi, selectReadStageMask_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]       selectReadStageMask_lo_hi_hi_hi_lo = {selectReadStageMask_lo_hi_hi_hi_lo_hi, selectReadStageMask_lo_hi_hi_hi_lo_lo};
  wire [127:0]       selectReadStageMask_lo_hi_hi_hi_hi_lo = {selectReadStageMask_lo_hi_hi_hi_hi_lo_hi, selectReadStageMask_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]       selectReadStageMask_lo_hi_hi_hi_hi_hi = {selectReadStageMask_lo_hi_hi_hi_hi_hi_hi, selectReadStageMask_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]       selectReadStageMask_lo_hi_hi_hi_hi = {selectReadStageMask_lo_hi_hi_hi_hi_hi, selectReadStageMask_lo_hi_hi_hi_hi_lo};
  wire [511:0]       selectReadStageMask_lo_hi_hi_hi = {selectReadStageMask_lo_hi_hi_hi_hi, selectReadStageMask_lo_hi_hi_hi_lo};
  wire [1023:0]      selectReadStageMask_lo_hi_hi = {selectReadStageMask_lo_hi_hi_hi, selectReadStageMask_lo_hi_hi_lo};
  wire [2047:0]      selectReadStageMask_lo_hi = {selectReadStageMask_lo_hi_hi, selectReadStageMask_lo_hi_lo};
  wire [4095:0]      selectReadStageMask_lo = {selectReadStageMask_lo_hi, selectReadStageMask_lo_lo};
  wire [127:0]       selectReadStageMask_hi_lo_lo_lo_lo_lo = {selectReadStageMask_hi_lo_lo_lo_lo_lo_hi, selectReadStageMask_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]       selectReadStageMask_hi_lo_lo_lo_lo_hi = {selectReadStageMask_hi_lo_lo_lo_lo_hi_hi, selectReadStageMask_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]       selectReadStageMask_hi_lo_lo_lo_lo = {selectReadStageMask_hi_lo_lo_lo_lo_hi, selectReadStageMask_hi_lo_lo_lo_lo_lo};
  wire [127:0]       selectReadStageMask_hi_lo_lo_lo_hi_lo = {selectReadStageMask_hi_lo_lo_lo_hi_lo_hi, selectReadStageMask_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]       selectReadStageMask_hi_lo_lo_lo_hi_hi = {selectReadStageMask_hi_lo_lo_lo_hi_hi_hi, selectReadStageMask_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]       selectReadStageMask_hi_lo_lo_lo_hi = {selectReadStageMask_hi_lo_lo_lo_hi_hi, selectReadStageMask_hi_lo_lo_lo_hi_lo};
  wire [511:0]       selectReadStageMask_hi_lo_lo_lo = {selectReadStageMask_hi_lo_lo_lo_hi, selectReadStageMask_hi_lo_lo_lo_lo};
  wire [127:0]       selectReadStageMask_hi_lo_lo_hi_lo_lo = {selectReadStageMask_hi_lo_lo_hi_lo_lo_hi, selectReadStageMask_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]       selectReadStageMask_hi_lo_lo_hi_lo_hi = {selectReadStageMask_hi_lo_lo_hi_lo_hi_hi, selectReadStageMask_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]       selectReadStageMask_hi_lo_lo_hi_lo = {selectReadStageMask_hi_lo_lo_hi_lo_hi, selectReadStageMask_hi_lo_lo_hi_lo_lo};
  wire [127:0]       selectReadStageMask_hi_lo_lo_hi_hi_lo = {selectReadStageMask_hi_lo_lo_hi_hi_lo_hi, selectReadStageMask_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]       selectReadStageMask_hi_lo_lo_hi_hi_hi = {selectReadStageMask_hi_lo_lo_hi_hi_hi_hi, selectReadStageMask_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]       selectReadStageMask_hi_lo_lo_hi_hi = {selectReadStageMask_hi_lo_lo_hi_hi_hi, selectReadStageMask_hi_lo_lo_hi_hi_lo};
  wire [511:0]       selectReadStageMask_hi_lo_lo_hi = {selectReadStageMask_hi_lo_lo_hi_hi, selectReadStageMask_hi_lo_lo_hi_lo};
  wire [1023:0]      selectReadStageMask_hi_lo_lo = {selectReadStageMask_hi_lo_lo_hi, selectReadStageMask_hi_lo_lo_lo};
  wire [127:0]       selectReadStageMask_hi_lo_hi_lo_lo_lo = {selectReadStageMask_hi_lo_hi_lo_lo_lo_hi, selectReadStageMask_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]       selectReadStageMask_hi_lo_hi_lo_lo_hi = {selectReadStageMask_hi_lo_hi_lo_lo_hi_hi, selectReadStageMask_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]       selectReadStageMask_hi_lo_hi_lo_lo = {selectReadStageMask_hi_lo_hi_lo_lo_hi, selectReadStageMask_hi_lo_hi_lo_lo_lo};
  wire [127:0]       selectReadStageMask_hi_lo_hi_lo_hi_lo = {selectReadStageMask_hi_lo_hi_lo_hi_lo_hi, selectReadStageMask_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]       selectReadStageMask_hi_lo_hi_lo_hi_hi = {selectReadStageMask_hi_lo_hi_lo_hi_hi_hi, selectReadStageMask_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]       selectReadStageMask_hi_lo_hi_lo_hi = {selectReadStageMask_hi_lo_hi_lo_hi_hi, selectReadStageMask_hi_lo_hi_lo_hi_lo};
  wire [511:0]       selectReadStageMask_hi_lo_hi_lo = {selectReadStageMask_hi_lo_hi_lo_hi, selectReadStageMask_hi_lo_hi_lo_lo};
  wire [127:0]       selectReadStageMask_hi_lo_hi_hi_lo_lo = {selectReadStageMask_hi_lo_hi_hi_lo_lo_hi, selectReadStageMask_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]       selectReadStageMask_hi_lo_hi_hi_lo_hi = {selectReadStageMask_hi_lo_hi_hi_lo_hi_hi, selectReadStageMask_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]       selectReadStageMask_hi_lo_hi_hi_lo = {selectReadStageMask_hi_lo_hi_hi_lo_hi, selectReadStageMask_hi_lo_hi_hi_lo_lo};
  wire [127:0]       selectReadStageMask_hi_lo_hi_hi_hi_lo = {selectReadStageMask_hi_lo_hi_hi_hi_lo_hi, selectReadStageMask_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]       selectReadStageMask_hi_lo_hi_hi_hi_hi = {selectReadStageMask_hi_lo_hi_hi_hi_hi_hi, selectReadStageMask_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]       selectReadStageMask_hi_lo_hi_hi_hi = {selectReadStageMask_hi_lo_hi_hi_hi_hi, selectReadStageMask_hi_lo_hi_hi_hi_lo};
  wire [511:0]       selectReadStageMask_hi_lo_hi_hi = {selectReadStageMask_hi_lo_hi_hi_hi, selectReadStageMask_hi_lo_hi_hi_lo};
  wire [1023:0]      selectReadStageMask_hi_lo_hi = {selectReadStageMask_hi_lo_hi_hi, selectReadStageMask_hi_lo_hi_lo};
  wire [2047:0]      selectReadStageMask_hi_lo = {selectReadStageMask_hi_lo_hi, selectReadStageMask_hi_lo_lo};
  wire [127:0]       selectReadStageMask_hi_hi_lo_lo_lo_lo = {selectReadStageMask_hi_hi_lo_lo_lo_lo_hi, selectReadStageMask_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]       selectReadStageMask_hi_hi_lo_lo_lo_hi = {selectReadStageMask_hi_hi_lo_lo_lo_hi_hi, selectReadStageMask_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]       selectReadStageMask_hi_hi_lo_lo_lo = {selectReadStageMask_hi_hi_lo_lo_lo_hi, selectReadStageMask_hi_hi_lo_lo_lo_lo};
  wire [127:0]       selectReadStageMask_hi_hi_lo_lo_hi_lo = {selectReadStageMask_hi_hi_lo_lo_hi_lo_hi, selectReadStageMask_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]       selectReadStageMask_hi_hi_lo_lo_hi_hi = {selectReadStageMask_hi_hi_lo_lo_hi_hi_hi, selectReadStageMask_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]       selectReadStageMask_hi_hi_lo_lo_hi = {selectReadStageMask_hi_hi_lo_lo_hi_hi, selectReadStageMask_hi_hi_lo_lo_hi_lo};
  wire [511:0]       selectReadStageMask_hi_hi_lo_lo = {selectReadStageMask_hi_hi_lo_lo_hi, selectReadStageMask_hi_hi_lo_lo_lo};
  wire [127:0]       selectReadStageMask_hi_hi_lo_hi_lo_lo = {selectReadStageMask_hi_hi_lo_hi_lo_lo_hi, selectReadStageMask_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]       selectReadStageMask_hi_hi_lo_hi_lo_hi = {selectReadStageMask_hi_hi_lo_hi_lo_hi_hi, selectReadStageMask_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]       selectReadStageMask_hi_hi_lo_hi_lo = {selectReadStageMask_hi_hi_lo_hi_lo_hi, selectReadStageMask_hi_hi_lo_hi_lo_lo};
  wire [127:0]       selectReadStageMask_hi_hi_lo_hi_hi_lo = {selectReadStageMask_hi_hi_lo_hi_hi_lo_hi, selectReadStageMask_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]       selectReadStageMask_hi_hi_lo_hi_hi_hi = {selectReadStageMask_hi_hi_lo_hi_hi_hi_hi, selectReadStageMask_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]       selectReadStageMask_hi_hi_lo_hi_hi = {selectReadStageMask_hi_hi_lo_hi_hi_hi, selectReadStageMask_hi_hi_lo_hi_hi_lo};
  wire [511:0]       selectReadStageMask_hi_hi_lo_hi = {selectReadStageMask_hi_hi_lo_hi_hi, selectReadStageMask_hi_hi_lo_hi_lo};
  wire [1023:0]      selectReadStageMask_hi_hi_lo = {selectReadStageMask_hi_hi_lo_hi, selectReadStageMask_hi_hi_lo_lo};
  wire [127:0]       selectReadStageMask_hi_hi_hi_lo_lo_lo = {selectReadStageMask_hi_hi_hi_lo_lo_lo_hi, selectReadStageMask_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]       selectReadStageMask_hi_hi_hi_lo_lo_hi = {selectReadStageMask_hi_hi_hi_lo_lo_hi_hi, selectReadStageMask_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]       selectReadStageMask_hi_hi_hi_lo_lo = {selectReadStageMask_hi_hi_hi_lo_lo_hi, selectReadStageMask_hi_hi_hi_lo_lo_lo};
  wire [127:0]       selectReadStageMask_hi_hi_hi_lo_hi_lo = {selectReadStageMask_hi_hi_hi_lo_hi_lo_hi, selectReadStageMask_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]       selectReadStageMask_hi_hi_hi_lo_hi_hi = {selectReadStageMask_hi_hi_hi_lo_hi_hi_hi, selectReadStageMask_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]       selectReadStageMask_hi_hi_hi_lo_hi = {selectReadStageMask_hi_hi_hi_lo_hi_hi, selectReadStageMask_hi_hi_hi_lo_hi_lo};
  wire [511:0]       selectReadStageMask_hi_hi_hi_lo = {selectReadStageMask_hi_hi_hi_lo_hi, selectReadStageMask_hi_hi_hi_lo_lo};
  wire [127:0]       selectReadStageMask_hi_hi_hi_hi_lo_lo = {selectReadStageMask_hi_hi_hi_hi_lo_lo_hi, selectReadStageMask_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]       selectReadStageMask_hi_hi_hi_hi_lo_hi = {selectReadStageMask_hi_hi_hi_hi_lo_hi_hi, selectReadStageMask_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]       selectReadStageMask_hi_hi_hi_hi_lo = {selectReadStageMask_hi_hi_hi_hi_lo_hi, selectReadStageMask_hi_hi_hi_hi_lo_lo};
  wire [127:0]       selectReadStageMask_hi_hi_hi_hi_hi_lo = {selectReadStageMask_hi_hi_hi_hi_hi_lo_hi, selectReadStageMask_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]       selectReadStageMask_hi_hi_hi_hi_hi_hi = {selectReadStageMask_hi_hi_hi_hi_hi_hi_hi, selectReadStageMask_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]       selectReadStageMask_hi_hi_hi_hi_hi = {selectReadStageMask_hi_hi_hi_hi_hi_hi, selectReadStageMask_hi_hi_hi_hi_hi_lo};
  wire [511:0]       selectReadStageMask_hi_hi_hi_hi = {selectReadStageMask_hi_hi_hi_hi_hi, selectReadStageMask_hi_hi_hi_hi_lo};
  wire [1023:0]      selectReadStageMask_hi_hi_hi = {selectReadStageMask_hi_hi_hi_hi, selectReadStageMask_hi_hi_hi_lo};
  wire [2047:0]      selectReadStageMask_hi_hi = {selectReadStageMask_hi_hi_hi, selectReadStageMask_hi_hi_lo};
  wire [4095:0]      selectReadStageMask_hi = {selectReadStageMask_hi_hi, selectReadStageMask_hi_lo};
  wire [2047:0][3:0] _GEN_142 =
    {{selectReadStageMask_hi[4095:4092]},
     {selectReadStageMask_hi[4091:4088]},
     {selectReadStageMask_hi[4087:4084]},
     {selectReadStageMask_hi[4083:4080]},
     {selectReadStageMask_hi[4079:4076]},
     {selectReadStageMask_hi[4075:4072]},
     {selectReadStageMask_hi[4071:4068]},
     {selectReadStageMask_hi[4067:4064]},
     {selectReadStageMask_hi[4063:4060]},
     {selectReadStageMask_hi[4059:4056]},
     {selectReadStageMask_hi[4055:4052]},
     {selectReadStageMask_hi[4051:4048]},
     {selectReadStageMask_hi[4047:4044]},
     {selectReadStageMask_hi[4043:4040]},
     {selectReadStageMask_hi[4039:4036]},
     {selectReadStageMask_hi[4035:4032]},
     {selectReadStageMask_hi[4031:4028]},
     {selectReadStageMask_hi[4027:4024]},
     {selectReadStageMask_hi[4023:4020]},
     {selectReadStageMask_hi[4019:4016]},
     {selectReadStageMask_hi[4015:4012]},
     {selectReadStageMask_hi[4011:4008]},
     {selectReadStageMask_hi[4007:4004]},
     {selectReadStageMask_hi[4003:4000]},
     {selectReadStageMask_hi[3999:3996]},
     {selectReadStageMask_hi[3995:3992]},
     {selectReadStageMask_hi[3991:3988]},
     {selectReadStageMask_hi[3987:3984]},
     {selectReadStageMask_hi[3983:3980]},
     {selectReadStageMask_hi[3979:3976]},
     {selectReadStageMask_hi[3975:3972]},
     {selectReadStageMask_hi[3971:3968]},
     {selectReadStageMask_hi[3967:3964]},
     {selectReadStageMask_hi[3963:3960]},
     {selectReadStageMask_hi[3959:3956]},
     {selectReadStageMask_hi[3955:3952]},
     {selectReadStageMask_hi[3951:3948]},
     {selectReadStageMask_hi[3947:3944]},
     {selectReadStageMask_hi[3943:3940]},
     {selectReadStageMask_hi[3939:3936]},
     {selectReadStageMask_hi[3935:3932]},
     {selectReadStageMask_hi[3931:3928]},
     {selectReadStageMask_hi[3927:3924]},
     {selectReadStageMask_hi[3923:3920]},
     {selectReadStageMask_hi[3919:3916]},
     {selectReadStageMask_hi[3915:3912]},
     {selectReadStageMask_hi[3911:3908]},
     {selectReadStageMask_hi[3907:3904]},
     {selectReadStageMask_hi[3903:3900]},
     {selectReadStageMask_hi[3899:3896]},
     {selectReadStageMask_hi[3895:3892]},
     {selectReadStageMask_hi[3891:3888]},
     {selectReadStageMask_hi[3887:3884]},
     {selectReadStageMask_hi[3883:3880]},
     {selectReadStageMask_hi[3879:3876]},
     {selectReadStageMask_hi[3875:3872]},
     {selectReadStageMask_hi[3871:3868]},
     {selectReadStageMask_hi[3867:3864]},
     {selectReadStageMask_hi[3863:3860]},
     {selectReadStageMask_hi[3859:3856]},
     {selectReadStageMask_hi[3855:3852]},
     {selectReadStageMask_hi[3851:3848]},
     {selectReadStageMask_hi[3847:3844]},
     {selectReadStageMask_hi[3843:3840]},
     {selectReadStageMask_hi[3839:3836]},
     {selectReadStageMask_hi[3835:3832]},
     {selectReadStageMask_hi[3831:3828]},
     {selectReadStageMask_hi[3827:3824]},
     {selectReadStageMask_hi[3823:3820]},
     {selectReadStageMask_hi[3819:3816]},
     {selectReadStageMask_hi[3815:3812]},
     {selectReadStageMask_hi[3811:3808]},
     {selectReadStageMask_hi[3807:3804]},
     {selectReadStageMask_hi[3803:3800]},
     {selectReadStageMask_hi[3799:3796]},
     {selectReadStageMask_hi[3795:3792]},
     {selectReadStageMask_hi[3791:3788]},
     {selectReadStageMask_hi[3787:3784]},
     {selectReadStageMask_hi[3783:3780]},
     {selectReadStageMask_hi[3779:3776]},
     {selectReadStageMask_hi[3775:3772]},
     {selectReadStageMask_hi[3771:3768]},
     {selectReadStageMask_hi[3767:3764]},
     {selectReadStageMask_hi[3763:3760]},
     {selectReadStageMask_hi[3759:3756]},
     {selectReadStageMask_hi[3755:3752]},
     {selectReadStageMask_hi[3751:3748]},
     {selectReadStageMask_hi[3747:3744]},
     {selectReadStageMask_hi[3743:3740]},
     {selectReadStageMask_hi[3739:3736]},
     {selectReadStageMask_hi[3735:3732]},
     {selectReadStageMask_hi[3731:3728]},
     {selectReadStageMask_hi[3727:3724]},
     {selectReadStageMask_hi[3723:3720]},
     {selectReadStageMask_hi[3719:3716]},
     {selectReadStageMask_hi[3715:3712]},
     {selectReadStageMask_hi[3711:3708]},
     {selectReadStageMask_hi[3707:3704]},
     {selectReadStageMask_hi[3703:3700]},
     {selectReadStageMask_hi[3699:3696]},
     {selectReadStageMask_hi[3695:3692]},
     {selectReadStageMask_hi[3691:3688]},
     {selectReadStageMask_hi[3687:3684]},
     {selectReadStageMask_hi[3683:3680]},
     {selectReadStageMask_hi[3679:3676]},
     {selectReadStageMask_hi[3675:3672]},
     {selectReadStageMask_hi[3671:3668]},
     {selectReadStageMask_hi[3667:3664]},
     {selectReadStageMask_hi[3663:3660]},
     {selectReadStageMask_hi[3659:3656]},
     {selectReadStageMask_hi[3655:3652]},
     {selectReadStageMask_hi[3651:3648]},
     {selectReadStageMask_hi[3647:3644]},
     {selectReadStageMask_hi[3643:3640]},
     {selectReadStageMask_hi[3639:3636]},
     {selectReadStageMask_hi[3635:3632]},
     {selectReadStageMask_hi[3631:3628]},
     {selectReadStageMask_hi[3627:3624]},
     {selectReadStageMask_hi[3623:3620]},
     {selectReadStageMask_hi[3619:3616]},
     {selectReadStageMask_hi[3615:3612]},
     {selectReadStageMask_hi[3611:3608]},
     {selectReadStageMask_hi[3607:3604]},
     {selectReadStageMask_hi[3603:3600]},
     {selectReadStageMask_hi[3599:3596]},
     {selectReadStageMask_hi[3595:3592]},
     {selectReadStageMask_hi[3591:3588]},
     {selectReadStageMask_hi[3587:3584]},
     {selectReadStageMask_hi[3583:3580]},
     {selectReadStageMask_hi[3579:3576]},
     {selectReadStageMask_hi[3575:3572]},
     {selectReadStageMask_hi[3571:3568]},
     {selectReadStageMask_hi[3567:3564]},
     {selectReadStageMask_hi[3563:3560]},
     {selectReadStageMask_hi[3559:3556]},
     {selectReadStageMask_hi[3555:3552]},
     {selectReadStageMask_hi[3551:3548]},
     {selectReadStageMask_hi[3547:3544]},
     {selectReadStageMask_hi[3543:3540]},
     {selectReadStageMask_hi[3539:3536]},
     {selectReadStageMask_hi[3535:3532]},
     {selectReadStageMask_hi[3531:3528]},
     {selectReadStageMask_hi[3527:3524]},
     {selectReadStageMask_hi[3523:3520]},
     {selectReadStageMask_hi[3519:3516]},
     {selectReadStageMask_hi[3515:3512]},
     {selectReadStageMask_hi[3511:3508]},
     {selectReadStageMask_hi[3507:3504]},
     {selectReadStageMask_hi[3503:3500]},
     {selectReadStageMask_hi[3499:3496]},
     {selectReadStageMask_hi[3495:3492]},
     {selectReadStageMask_hi[3491:3488]},
     {selectReadStageMask_hi[3487:3484]},
     {selectReadStageMask_hi[3483:3480]},
     {selectReadStageMask_hi[3479:3476]},
     {selectReadStageMask_hi[3475:3472]},
     {selectReadStageMask_hi[3471:3468]},
     {selectReadStageMask_hi[3467:3464]},
     {selectReadStageMask_hi[3463:3460]},
     {selectReadStageMask_hi[3459:3456]},
     {selectReadStageMask_hi[3455:3452]},
     {selectReadStageMask_hi[3451:3448]},
     {selectReadStageMask_hi[3447:3444]},
     {selectReadStageMask_hi[3443:3440]},
     {selectReadStageMask_hi[3439:3436]},
     {selectReadStageMask_hi[3435:3432]},
     {selectReadStageMask_hi[3431:3428]},
     {selectReadStageMask_hi[3427:3424]},
     {selectReadStageMask_hi[3423:3420]},
     {selectReadStageMask_hi[3419:3416]},
     {selectReadStageMask_hi[3415:3412]},
     {selectReadStageMask_hi[3411:3408]},
     {selectReadStageMask_hi[3407:3404]},
     {selectReadStageMask_hi[3403:3400]},
     {selectReadStageMask_hi[3399:3396]},
     {selectReadStageMask_hi[3395:3392]},
     {selectReadStageMask_hi[3391:3388]},
     {selectReadStageMask_hi[3387:3384]},
     {selectReadStageMask_hi[3383:3380]},
     {selectReadStageMask_hi[3379:3376]},
     {selectReadStageMask_hi[3375:3372]},
     {selectReadStageMask_hi[3371:3368]},
     {selectReadStageMask_hi[3367:3364]},
     {selectReadStageMask_hi[3363:3360]},
     {selectReadStageMask_hi[3359:3356]},
     {selectReadStageMask_hi[3355:3352]},
     {selectReadStageMask_hi[3351:3348]},
     {selectReadStageMask_hi[3347:3344]},
     {selectReadStageMask_hi[3343:3340]},
     {selectReadStageMask_hi[3339:3336]},
     {selectReadStageMask_hi[3335:3332]},
     {selectReadStageMask_hi[3331:3328]},
     {selectReadStageMask_hi[3327:3324]},
     {selectReadStageMask_hi[3323:3320]},
     {selectReadStageMask_hi[3319:3316]},
     {selectReadStageMask_hi[3315:3312]},
     {selectReadStageMask_hi[3311:3308]},
     {selectReadStageMask_hi[3307:3304]},
     {selectReadStageMask_hi[3303:3300]},
     {selectReadStageMask_hi[3299:3296]},
     {selectReadStageMask_hi[3295:3292]},
     {selectReadStageMask_hi[3291:3288]},
     {selectReadStageMask_hi[3287:3284]},
     {selectReadStageMask_hi[3283:3280]},
     {selectReadStageMask_hi[3279:3276]},
     {selectReadStageMask_hi[3275:3272]},
     {selectReadStageMask_hi[3271:3268]},
     {selectReadStageMask_hi[3267:3264]},
     {selectReadStageMask_hi[3263:3260]},
     {selectReadStageMask_hi[3259:3256]},
     {selectReadStageMask_hi[3255:3252]},
     {selectReadStageMask_hi[3251:3248]},
     {selectReadStageMask_hi[3247:3244]},
     {selectReadStageMask_hi[3243:3240]},
     {selectReadStageMask_hi[3239:3236]},
     {selectReadStageMask_hi[3235:3232]},
     {selectReadStageMask_hi[3231:3228]},
     {selectReadStageMask_hi[3227:3224]},
     {selectReadStageMask_hi[3223:3220]},
     {selectReadStageMask_hi[3219:3216]},
     {selectReadStageMask_hi[3215:3212]},
     {selectReadStageMask_hi[3211:3208]},
     {selectReadStageMask_hi[3207:3204]},
     {selectReadStageMask_hi[3203:3200]},
     {selectReadStageMask_hi[3199:3196]},
     {selectReadStageMask_hi[3195:3192]},
     {selectReadStageMask_hi[3191:3188]},
     {selectReadStageMask_hi[3187:3184]},
     {selectReadStageMask_hi[3183:3180]},
     {selectReadStageMask_hi[3179:3176]},
     {selectReadStageMask_hi[3175:3172]},
     {selectReadStageMask_hi[3171:3168]},
     {selectReadStageMask_hi[3167:3164]},
     {selectReadStageMask_hi[3163:3160]},
     {selectReadStageMask_hi[3159:3156]},
     {selectReadStageMask_hi[3155:3152]},
     {selectReadStageMask_hi[3151:3148]},
     {selectReadStageMask_hi[3147:3144]},
     {selectReadStageMask_hi[3143:3140]},
     {selectReadStageMask_hi[3139:3136]},
     {selectReadStageMask_hi[3135:3132]},
     {selectReadStageMask_hi[3131:3128]},
     {selectReadStageMask_hi[3127:3124]},
     {selectReadStageMask_hi[3123:3120]},
     {selectReadStageMask_hi[3119:3116]},
     {selectReadStageMask_hi[3115:3112]},
     {selectReadStageMask_hi[3111:3108]},
     {selectReadStageMask_hi[3107:3104]},
     {selectReadStageMask_hi[3103:3100]},
     {selectReadStageMask_hi[3099:3096]},
     {selectReadStageMask_hi[3095:3092]},
     {selectReadStageMask_hi[3091:3088]},
     {selectReadStageMask_hi[3087:3084]},
     {selectReadStageMask_hi[3083:3080]},
     {selectReadStageMask_hi[3079:3076]},
     {selectReadStageMask_hi[3075:3072]},
     {selectReadStageMask_hi[3071:3068]},
     {selectReadStageMask_hi[3067:3064]},
     {selectReadStageMask_hi[3063:3060]},
     {selectReadStageMask_hi[3059:3056]},
     {selectReadStageMask_hi[3055:3052]},
     {selectReadStageMask_hi[3051:3048]},
     {selectReadStageMask_hi[3047:3044]},
     {selectReadStageMask_hi[3043:3040]},
     {selectReadStageMask_hi[3039:3036]},
     {selectReadStageMask_hi[3035:3032]},
     {selectReadStageMask_hi[3031:3028]},
     {selectReadStageMask_hi[3027:3024]},
     {selectReadStageMask_hi[3023:3020]},
     {selectReadStageMask_hi[3019:3016]},
     {selectReadStageMask_hi[3015:3012]},
     {selectReadStageMask_hi[3011:3008]},
     {selectReadStageMask_hi[3007:3004]},
     {selectReadStageMask_hi[3003:3000]},
     {selectReadStageMask_hi[2999:2996]},
     {selectReadStageMask_hi[2995:2992]},
     {selectReadStageMask_hi[2991:2988]},
     {selectReadStageMask_hi[2987:2984]},
     {selectReadStageMask_hi[2983:2980]},
     {selectReadStageMask_hi[2979:2976]},
     {selectReadStageMask_hi[2975:2972]},
     {selectReadStageMask_hi[2971:2968]},
     {selectReadStageMask_hi[2967:2964]},
     {selectReadStageMask_hi[2963:2960]},
     {selectReadStageMask_hi[2959:2956]},
     {selectReadStageMask_hi[2955:2952]},
     {selectReadStageMask_hi[2951:2948]},
     {selectReadStageMask_hi[2947:2944]},
     {selectReadStageMask_hi[2943:2940]},
     {selectReadStageMask_hi[2939:2936]},
     {selectReadStageMask_hi[2935:2932]},
     {selectReadStageMask_hi[2931:2928]},
     {selectReadStageMask_hi[2927:2924]},
     {selectReadStageMask_hi[2923:2920]},
     {selectReadStageMask_hi[2919:2916]},
     {selectReadStageMask_hi[2915:2912]},
     {selectReadStageMask_hi[2911:2908]},
     {selectReadStageMask_hi[2907:2904]},
     {selectReadStageMask_hi[2903:2900]},
     {selectReadStageMask_hi[2899:2896]},
     {selectReadStageMask_hi[2895:2892]},
     {selectReadStageMask_hi[2891:2888]},
     {selectReadStageMask_hi[2887:2884]},
     {selectReadStageMask_hi[2883:2880]},
     {selectReadStageMask_hi[2879:2876]},
     {selectReadStageMask_hi[2875:2872]},
     {selectReadStageMask_hi[2871:2868]},
     {selectReadStageMask_hi[2867:2864]},
     {selectReadStageMask_hi[2863:2860]},
     {selectReadStageMask_hi[2859:2856]},
     {selectReadStageMask_hi[2855:2852]},
     {selectReadStageMask_hi[2851:2848]},
     {selectReadStageMask_hi[2847:2844]},
     {selectReadStageMask_hi[2843:2840]},
     {selectReadStageMask_hi[2839:2836]},
     {selectReadStageMask_hi[2835:2832]},
     {selectReadStageMask_hi[2831:2828]},
     {selectReadStageMask_hi[2827:2824]},
     {selectReadStageMask_hi[2823:2820]},
     {selectReadStageMask_hi[2819:2816]},
     {selectReadStageMask_hi[2815:2812]},
     {selectReadStageMask_hi[2811:2808]},
     {selectReadStageMask_hi[2807:2804]},
     {selectReadStageMask_hi[2803:2800]},
     {selectReadStageMask_hi[2799:2796]},
     {selectReadStageMask_hi[2795:2792]},
     {selectReadStageMask_hi[2791:2788]},
     {selectReadStageMask_hi[2787:2784]},
     {selectReadStageMask_hi[2783:2780]},
     {selectReadStageMask_hi[2779:2776]},
     {selectReadStageMask_hi[2775:2772]},
     {selectReadStageMask_hi[2771:2768]},
     {selectReadStageMask_hi[2767:2764]},
     {selectReadStageMask_hi[2763:2760]},
     {selectReadStageMask_hi[2759:2756]},
     {selectReadStageMask_hi[2755:2752]},
     {selectReadStageMask_hi[2751:2748]},
     {selectReadStageMask_hi[2747:2744]},
     {selectReadStageMask_hi[2743:2740]},
     {selectReadStageMask_hi[2739:2736]},
     {selectReadStageMask_hi[2735:2732]},
     {selectReadStageMask_hi[2731:2728]},
     {selectReadStageMask_hi[2727:2724]},
     {selectReadStageMask_hi[2723:2720]},
     {selectReadStageMask_hi[2719:2716]},
     {selectReadStageMask_hi[2715:2712]},
     {selectReadStageMask_hi[2711:2708]},
     {selectReadStageMask_hi[2707:2704]},
     {selectReadStageMask_hi[2703:2700]},
     {selectReadStageMask_hi[2699:2696]},
     {selectReadStageMask_hi[2695:2692]},
     {selectReadStageMask_hi[2691:2688]},
     {selectReadStageMask_hi[2687:2684]},
     {selectReadStageMask_hi[2683:2680]},
     {selectReadStageMask_hi[2679:2676]},
     {selectReadStageMask_hi[2675:2672]},
     {selectReadStageMask_hi[2671:2668]},
     {selectReadStageMask_hi[2667:2664]},
     {selectReadStageMask_hi[2663:2660]},
     {selectReadStageMask_hi[2659:2656]},
     {selectReadStageMask_hi[2655:2652]},
     {selectReadStageMask_hi[2651:2648]},
     {selectReadStageMask_hi[2647:2644]},
     {selectReadStageMask_hi[2643:2640]},
     {selectReadStageMask_hi[2639:2636]},
     {selectReadStageMask_hi[2635:2632]},
     {selectReadStageMask_hi[2631:2628]},
     {selectReadStageMask_hi[2627:2624]},
     {selectReadStageMask_hi[2623:2620]},
     {selectReadStageMask_hi[2619:2616]},
     {selectReadStageMask_hi[2615:2612]},
     {selectReadStageMask_hi[2611:2608]},
     {selectReadStageMask_hi[2607:2604]},
     {selectReadStageMask_hi[2603:2600]},
     {selectReadStageMask_hi[2599:2596]},
     {selectReadStageMask_hi[2595:2592]},
     {selectReadStageMask_hi[2591:2588]},
     {selectReadStageMask_hi[2587:2584]},
     {selectReadStageMask_hi[2583:2580]},
     {selectReadStageMask_hi[2579:2576]},
     {selectReadStageMask_hi[2575:2572]},
     {selectReadStageMask_hi[2571:2568]},
     {selectReadStageMask_hi[2567:2564]},
     {selectReadStageMask_hi[2563:2560]},
     {selectReadStageMask_hi[2559:2556]},
     {selectReadStageMask_hi[2555:2552]},
     {selectReadStageMask_hi[2551:2548]},
     {selectReadStageMask_hi[2547:2544]},
     {selectReadStageMask_hi[2543:2540]},
     {selectReadStageMask_hi[2539:2536]},
     {selectReadStageMask_hi[2535:2532]},
     {selectReadStageMask_hi[2531:2528]},
     {selectReadStageMask_hi[2527:2524]},
     {selectReadStageMask_hi[2523:2520]},
     {selectReadStageMask_hi[2519:2516]},
     {selectReadStageMask_hi[2515:2512]},
     {selectReadStageMask_hi[2511:2508]},
     {selectReadStageMask_hi[2507:2504]},
     {selectReadStageMask_hi[2503:2500]},
     {selectReadStageMask_hi[2499:2496]},
     {selectReadStageMask_hi[2495:2492]},
     {selectReadStageMask_hi[2491:2488]},
     {selectReadStageMask_hi[2487:2484]},
     {selectReadStageMask_hi[2483:2480]},
     {selectReadStageMask_hi[2479:2476]},
     {selectReadStageMask_hi[2475:2472]},
     {selectReadStageMask_hi[2471:2468]},
     {selectReadStageMask_hi[2467:2464]},
     {selectReadStageMask_hi[2463:2460]},
     {selectReadStageMask_hi[2459:2456]},
     {selectReadStageMask_hi[2455:2452]},
     {selectReadStageMask_hi[2451:2448]},
     {selectReadStageMask_hi[2447:2444]},
     {selectReadStageMask_hi[2443:2440]},
     {selectReadStageMask_hi[2439:2436]},
     {selectReadStageMask_hi[2435:2432]},
     {selectReadStageMask_hi[2431:2428]},
     {selectReadStageMask_hi[2427:2424]},
     {selectReadStageMask_hi[2423:2420]},
     {selectReadStageMask_hi[2419:2416]},
     {selectReadStageMask_hi[2415:2412]},
     {selectReadStageMask_hi[2411:2408]},
     {selectReadStageMask_hi[2407:2404]},
     {selectReadStageMask_hi[2403:2400]},
     {selectReadStageMask_hi[2399:2396]},
     {selectReadStageMask_hi[2395:2392]},
     {selectReadStageMask_hi[2391:2388]},
     {selectReadStageMask_hi[2387:2384]},
     {selectReadStageMask_hi[2383:2380]},
     {selectReadStageMask_hi[2379:2376]},
     {selectReadStageMask_hi[2375:2372]},
     {selectReadStageMask_hi[2371:2368]},
     {selectReadStageMask_hi[2367:2364]},
     {selectReadStageMask_hi[2363:2360]},
     {selectReadStageMask_hi[2359:2356]},
     {selectReadStageMask_hi[2355:2352]},
     {selectReadStageMask_hi[2351:2348]},
     {selectReadStageMask_hi[2347:2344]},
     {selectReadStageMask_hi[2343:2340]},
     {selectReadStageMask_hi[2339:2336]},
     {selectReadStageMask_hi[2335:2332]},
     {selectReadStageMask_hi[2331:2328]},
     {selectReadStageMask_hi[2327:2324]},
     {selectReadStageMask_hi[2323:2320]},
     {selectReadStageMask_hi[2319:2316]},
     {selectReadStageMask_hi[2315:2312]},
     {selectReadStageMask_hi[2311:2308]},
     {selectReadStageMask_hi[2307:2304]},
     {selectReadStageMask_hi[2303:2300]},
     {selectReadStageMask_hi[2299:2296]},
     {selectReadStageMask_hi[2295:2292]},
     {selectReadStageMask_hi[2291:2288]},
     {selectReadStageMask_hi[2287:2284]},
     {selectReadStageMask_hi[2283:2280]},
     {selectReadStageMask_hi[2279:2276]},
     {selectReadStageMask_hi[2275:2272]},
     {selectReadStageMask_hi[2271:2268]},
     {selectReadStageMask_hi[2267:2264]},
     {selectReadStageMask_hi[2263:2260]},
     {selectReadStageMask_hi[2259:2256]},
     {selectReadStageMask_hi[2255:2252]},
     {selectReadStageMask_hi[2251:2248]},
     {selectReadStageMask_hi[2247:2244]},
     {selectReadStageMask_hi[2243:2240]},
     {selectReadStageMask_hi[2239:2236]},
     {selectReadStageMask_hi[2235:2232]},
     {selectReadStageMask_hi[2231:2228]},
     {selectReadStageMask_hi[2227:2224]},
     {selectReadStageMask_hi[2223:2220]},
     {selectReadStageMask_hi[2219:2216]},
     {selectReadStageMask_hi[2215:2212]},
     {selectReadStageMask_hi[2211:2208]},
     {selectReadStageMask_hi[2207:2204]},
     {selectReadStageMask_hi[2203:2200]},
     {selectReadStageMask_hi[2199:2196]},
     {selectReadStageMask_hi[2195:2192]},
     {selectReadStageMask_hi[2191:2188]},
     {selectReadStageMask_hi[2187:2184]},
     {selectReadStageMask_hi[2183:2180]},
     {selectReadStageMask_hi[2179:2176]},
     {selectReadStageMask_hi[2175:2172]},
     {selectReadStageMask_hi[2171:2168]},
     {selectReadStageMask_hi[2167:2164]},
     {selectReadStageMask_hi[2163:2160]},
     {selectReadStageMask_hi[2159:2156]},
     {selectReadStageMask_hi[2155:2152]},
     {selectReadStageMask_hi[2151:2148]},
     {selectReadStageMask_hi[2147:2144]},
     {selectReadStageMask_hi[2143:2140]},
     {selectReadStageMask_hi[2139:2136]},
     {selectReadStageMask_hi[2135:2132]},
     {selectReadStageMask_hi[2131:2128]},
     {selectReadStageMask_hi[2127:2124]},
     {selectReadStageMask_hi[2123:2120]},
     {selectReadStageMask_hi[2119:2116]},
     {selectReadStageMask_hi[2115:2112]},
     {selectReadStageMask_hi[2111:2108]},
     {selectReadStageMask_hi[2107:2104]},
     {selectReadStageMask_hi[2103:2100]},
     {selectReadStageMask_hi[2099:2096]},
     {selectReadStageMask_hi[2095:2092]},
     {selectReadStageMask_hi[2091:2088]},
     {selectReadStageMask_hi[2087:2084]},
     {selectReadStageMask_hi[2083:2080]},
     {selectReadStageMask_hi[2079:2076]},
     {selectReadStageMask_hi[2075:2072]},
     {selectReadStageMask_hi[2071:2068]},
     {selectReadStageMask_hi[2067:2064]},
     {selectReadStageMask_hi[2063:2060]},
     {selectReadStageMask_hi[2059:2056]},
     {selectReadStageMask_hi[2055:2052]},
     {selectReadStageMask_hi[2051:2048]},
     {selectReadStageMask_hi[2047:2044]},
     {selectReadStageMask_hi[2043:2040]},
     {selectReadStageMask_hi[2039:2036]},
     {selectReadStageMask_hi[2035:2032]},
     {selectReadStageMask_hi[2031:2028]},
     {selectReadStageMask_hi[2027:2024]},
     {selectReadStageMask_hi[2023:2020]},
     {selectReadStageMask_hi[2019:2016]},
     {selectReadStageMask_hi[2015:2012]},
     {selectReadStageMask_hi[2011:2008]},
     {selectReadStageMask_hi[2007:2004]},
     {selectReadStageMask_hi[2003:2000]},
     {selectReadStageMask_hi[1999:1996]},
     {selectReadStageMask_hi[1995:1992]},
     {selectReadStageMask_hi[1991:1988]},
     {selectReadStageMask_hi[1987:1984]},
     {selectReadStageMask_hi[1983:1980]},
     {selectReadStageMask_hi[1979:1976]},
     {selectReadStageMask_hi[1975:1972]},
     {selectReadStageMask_hi[1971:1968]},
     {selectReadStageMask_hi[1967:1964]},
     {selectReadStageMask_hi[1963:1960]},
     {selectReadStageMask_hi[1959:1956]},
     {selectReadStageMask_hi[1955:1952]},
     {selectReadStageMask_hi[1951:1948]},
     {selectReadStageMask_hi[1947:1944]},
     {selectReadStageMask_hi[1943:1940]},
     {selectReadStageMask_hi[1939:1936]},
     {selectReadStageMask_hi[1935:1932]},
     {selectReadStageMask_hi[1931:1928]},
     {selectReadStageMask_hi[1927:1924]},
     {selectReadStageMask_hi[1923:1920]},
     {selectReadStageMask_hi[1919:1916]},
     {selectReadStageMask_hi[1915:1912]},
     {selectReadStageMask_hi[1911:1908]},
     {selectReadStageMask_hi[1907:1904]},
     {selectReadStageMask_hi[1903:1900]},
     {selectReadStageMask_hi[1899:1896]},
     {selectReadStageMask_hi[1895:1892]},
     {selectReadStageMask_hi[1891:1888]},
     {selectReadStageMask_hi[1887:1884]},
     {selectReadStageMask_hi[1883:1880]},
     {selectReadStageMask_hi[1879:1876]},
     {selectReadStageMask_hi[1875:1872]},
     {selectReadStageMask_hi[1871:1868]},
     {selectReadStageMask_hi[1867:1864]},
     {selectReadStageMask_hi[1863:1860]},
     {selectReadStageMask_hi[1859:1856]},
     {selectReadStageMask_hi[1855:1852]},
     {selectReadStageMask_hi[1851:1848]},
     {selectReadStageMask_hi[1847:1844]},
     {selectReadStageMask_hi[1843:1840]},
     {selectReadStageMask_hi[1839:1836]},
     {selectReadStageMask_hi[1835:1832]},
     {selectReadStageMask_hi[1831:1828]},
     {selectReadStageMask_hi[1827:1824]},
     {selectReadStageMask_hi[1823:1820]},
     {selectReadStageMask_hi[1819:1816]},
     {selectReadStageMask_hi[1815:1812]},
     {selectReadStageMask_hi[1811:1808]},
     {selectReadStageMask_hi[1807:1804]},
     {selectReadStageMask_hi[1803:1800]},
     {selectReadStageMask_hi[1799:1796]},
     {selectReadStageMask_hi[1795:1792]},
     {selectReadStageMask_hi[1791:1788]},
     {selectReadStageMask_hi[1787:1784]},
     {selectReadStageMask_hi[1783:1780]},
     {selectReadStageMask_hi[1779:1776]},
     {selectReadStageMask_hi[1775:1772]},
     {selectReadStageMask_hi[1771:1768]},
     {selectReadStageMask_hi[1767:1764]},
     {selectReadStageMask_hi[1763:1760]},
     {selectReadStageMask_hi[1759:1756]},
     {selectReadStageMask_hi[1755:1752]},
     {selectReadStageMask_hi[1751:1748]},
     {selectReadStageMask_hi[1747:1744]},
     {selectReadStageMask_hi[1743:1740]},
     {selectReadStageMask_hi[1739:1736]},
     {selectReadStageMask_hi[1735:1732]},
     {selectReadStageMask_hi[1731:1728]},
     {selectReadStageMask_hi[1727:1724]},
     {selectReadStageMask_hi[1723:1720]},
     {selectReadStageMask_hi[1719:1716]},
     {selectReadStageMask_hi[1715:1712]},
     {selectReadStageMask_hi[1711:1708]},
     {selectReadStageMask_hi[1707:1704]},
     {selectReadStageMask_hi[1703:1700]},
     {selectReadStageMask_hi[1699:1696]},
     {selectReadStageMask_hi[1695:1692]},
     {selectReadStageMask_hi[1691:1688]},
     {selectReadStageMask_hi[1687:1684]},
     {selectReadStageMask_hi[1683:1680]},
     {selectReadStageMask_hi[1679:1676]},
     {selectReadStageMask_hi[1675:1672]},
     {selectReadStageMask_hi[1671:1668]},
     {selectReadStageMask_hi[1667:1664]},
     {selectReadStageMask_hi[1663:1660]},
     {selectReadStageMask_hi[1659:1656]},
     {selectReadStageMask_hi[1655:1652]},
     {selectReadStageMask_hi[1651:1648]},
     {selectReadStageMask_hi[1647:1644]},
     {selectReadStageMask_hi[1643:1640]},
     {selectReadStageMask_hi[1639:1636]},
     {selectReadStageMask_hi[1635:1632]},
     {selectReadStageMask_hi[1631:1628]},
     {selectReadStageMask_hi[1627:1624]},
     {selectReadStageMask_hi[1623:1620]},
     {selectReadStageMask_hi[1619:1616]},
     {selectReadStageMask_hi[1615:1612]},
     {selectReadStageMask_hi[1611:1608]},
     {selectReadStageMask_hi[1607:1604]},
     {selectReadStageMask_hi[1603:1600]},
     {selectReadStageMask_hi[1599:1596]},
     {selectReadStageMask_hi[1595:1592]},
     {selectReadStageMask_hi[1591:1588]},
     {selectReadStageMask_hi[1587:1584]},
     {selectReadStageMask_hi[1583:1580]},
     {selectReadStageMask_hi[1579:1576]},
     {selectReadStageMask_hi[1575:1572]},
     {selectReadStageMask_hi[1571:1568]},
     {selectReadStageMask_hi[1567:1564]},
     {selectReadStageMask_hi[1563:1560]},
     {selectReadStageMask_hi[1559:1556]},
     {selectReadStageMask_hi[1555:1552]},
     {selectReadStageMask_hi[1551:1548]},
     {selectReadStageMask_hi[1547:1544]},
     {selectReadStageMask_hi[1543:1540]},
     {selectReadStageMask_hi[1539:1536]},
     {selectReadStageMask_hi[1535:1532]},
     {selectReadStageMask_hi[1531:1528]},
     {selectReadStageMask_hi[1527:1524]},
     {selectReadStageMask_hi[1523:1520]},
     {selectReadStageMask_hi[1519:1516]},
     {selectReadStageMask_hi[1515:1512]},
     {selectReadStageMask_hi[1511:1508]},
     {selectReadStageMask_hi[1507:1504]},
     {selectReadStageMask_hi[1503:1500]},
     {selectReadStageMask_hi[1499:1496]},
     {selectReadStageMask_hi[1495:1492]},
     {selectReadStageMask_hi[1491:1488]},
     {selectReadStageMask_hi[1487:1484]},
     {selectReadStageMask_hi[1483:1480]},
     {selectReadStageMask_hi[1479:1476]},
     {selectReadStageMask_hi[1475:1472]},
     {selectReadStageMask_hi[1471:1468]},
     {selectReadStageMask_hi[1467:1464]},
     {selectReadStageMask_hi[1463:1460]},
     {selectReadStageMask_hi[1459:1456]},
     {selectReadStageMask_hi[1455:1452]},
     {selectReadStageMask_hi[1451:1448]},
     {selectReadStageMask_hi[1447:1444]},
     {selectReadStageMask_hi[1443:1440]},
     {selectReadStageMask_hi[1439:1436]},
     {selectReadStageMask_hi[1435:1432]},
     {selectReadStageMask_hi[1431:1428]},
     {selectReadStageMask_hi[1427:1424]},
     {selectReadStageMask_hi[1423:1420]},
     {selectReadStageMask_hi[1419:1416]},
     {selectReadStageMask_hi[1415:1412]},
     {selectReadStageMask_hi[1411:1408]},
     {selectReadStageMask_hi[1407:1404]},
     {selectReadStageMask_hi[1403:1400]},
     {selectReadStageMask_hi[1399:1396]},
     {selectReadStageMask_hi[1395:1392]},
     {selectReadStageMask_hi[1391:1388]},
     {selectReadStageMask_hi[1387:1384]},
     {selectReadStageMask_hi[1383:1380]},
     {selectReadStageMask_hi[1379:1376]},
     {selectReadStageMask_hi[1375:1372]},
     {selectReadStageMask_hi[1371:1368]},
     {selectReadStageMask_hi[1367:1364]},
     {selectReadStageMask_hi[1363:1360]},
     {selectReadStageMask_hi[1359:1356]},
     {selectReadStageMask_hi[1355:1352]},
     {selectReadStageMask_hi[1351:1348]},
     {selectReadStageMask_hi[1347:1344]},
     {selectReadStageMask_hi[1343:1340]},
     {selectReadStageMask_hi[1339:1336]},
     {selectReadStageMask_hi[1335:1332]},
     {selectReadStageMask_hi[1331:1328]},
     {selectReadStageMask_hi[1327:1324]},
     {selectReadStageMask_hi[1323:1320]},
     {selectReadStageMask_hi[1319:1316]},
     {selectReadStageMask_hi[1315:1312]},
     {selectReadStageMask_hi[1311:1308]},
     {selectReadStageMask_hi[1307:1304]},
     {selectReadStageMask_hi[1303:1300]},
     {selectReadStageMask_hi[1299:1296]},
     {selectReadStageMask_hi[1295:1292]},
     {selectReadStageMask_hi[1291:1288]},
     {selectReadStageMask_hi[1287:1284]},
     {selectReadStageMask_hi[1283:1280]},
     {selectReadStageMask_hi[1279:1276]},
     {selectReadStageMask_hi[1275:1272]},
     {selectReadStageMask_hi[1271:1268]},
     {selectReadStageMask_hi[1267:1264]},
     {selectReadStageMask_hi[1263:1260]},
     {selectReadStageMask_hi[1259:1256]},
     {selectReadStageMask_hi[1255:1252]},
     {selectReadStageMask_hi[1251:1248]},
     {selectReadStageMask_hi[1247:1244]},
     {selectReadStageMask_hi[1243:1240]},
     {selectReadStageMask_hi[1239:1236]},
     {selectReadStageMask_hi[1235:1232]},
     {selectReadStageMask_hi[1231:1228]},
     {selectReadStageMask_hi[1227:1224]},
     {selectReadStageMask_hi[1223:1220]},
     {selectReadStageMask_hi[1219:1216]},
     {selectReadStageMask_hi[1215:1212]},
     {selectReadStageMask_hi[1211:1208]},
     {selectReadStageMask_hi[1207:1204]},
     {selectReadStageMask_hi[1203:1200]},
     {selectReadStageMask_hi[1199:1196]},
     {selectReadStageMask_hi[1195:1192]},
     {selectReadStageMask_hi[1191:1188]},
     {selectReadStageMask_hi[1187:1184]},
     {selectReadStageMask_hi[1183:1180]},
     {selectReadStageMask_hi[1179:1176]},
     {selectReadStageMask_hi[1175:1172]},
     {selectReadStageMask_hi[1171:1168]},
     {selectReadStageMask_hi[1167:1164]},
     {selectReadStageMask_hi[1163:1160]},
     {selectReadStageMask_hi[1159:1156]},
     {selectReadStageMask_hi[1155:1152]},
     {selectReadStageMask_hi[1151:1148]},
     {selectReadStageMask_hi[1147:1144]},
     {selectReadStageMask_hi[1143:1140]},
     {selectReadStageMask_hi[1139:1136]},
     {selectReadStageMask_hi[1135:1132]},
     {selectReadStageMask_hi[1131:1128]},
     {selectReadStageMask_hi[1127:1124]},
     {selectReadStageMask_hi[1123:1120]},
     {selectReadStageMask_hi[1119:1116]},
     {selectReadStageMask_hi[1115:1112]},
     {selectReadStageMask_hi[1111:1108]},
     {selectReadStageMask_hi[1107:1104]},
     {selectReadStageMask_hi[1103:1100]},
     {selectReadStageMask_hi[1099:1096]},
     {selectReadStageMask_hi[1095:1092]},
     {selectReadStageMask_hi[1091:1088]},
     {selectReadStageMask_hi[1087:1084]},
     {selectReadStageMask_hi[1083:1080]},
     {selectReadStageMask_hi[1079:1076]},
     {selectReadStageMask_hi[1075:1072]},
     {selectReadStageMask_hi[1071:1068]},
     {selectReadStageMask_hi[1067:1064]},
     {selectReadStageMask_hi[1063:1060]},
     {selectReadStageMask_hi[1059:1056]},
     {selectReadStageMask_hi[1055:1052]},
     {selectReadStageMask_hi[1051:1048]},
     {selectReadStageMask_hi[1047:1044]},
     {selectReadStageMask_hi[1043:1040]},
     {selectReadStageMask_hi[1039:1036]},
     {selectReadStageMask_hi[1035:1032]},
     {selectReadStageMask_hi[1031:1028]},
     {selectReadStageMask_hi[1027:1024]},
     {selectReadStageMask_hi[1023:1020]},
     {selectReadStageMask_hi[1019:1016]},
     {selectReadStageMask_hi[1015:1012]},
     {selectReadStageMask_hi[1011:1008]},
     {selectReadStageMask_hi[1007:1004]},
     {selectReadStageMask_hi[1003:1000]},
     {selectReadStageMask_hi[999:996]},
     {selectReadStageMask_hi[995:992]},
     {selectReadStageMask_hi[991:988]},
     {selectReadStageMask_hi[987:984]},
     {selectReadStageMask_hi[983:980]},
     {selectReadStageMask_hi[979:976]},
     {selectReadStageMask_hi[975:972]},
     {selectReadStageMask_hi[971:968]},
     {selectReadStageMask_hi[967:964]},
     {selectReadStageMask_hi[963:960]},
     {selectReadStageMask_hi[959:956]},
     {selectReadStageMask_hi[955:952]},
     {selectReadStageMask_hi[951:948]},
     {selectReadStageMask_hi[947:944]},
     {selectReadStageMask_hi[943:940]},
     {selectReadStageMask_hi[939:936]},
     {selectReadStageMask_hi[935:932]},
     {selectReadStageMask_hi[931:928]},
     {selectReadStageMask_hi[927:924]},
     {selectReadStageMask_hi[923:920]},
     {selectReadStageMask_hi[919:916]},
     {selectReadStageMask_hi[915:912]},
     {selectReadStageMask_hi[911:908]},
     {selectReadStageMask_hi[907:904]},
     {selectReadStageMask_hi[903:900]},
     {selectReadStageMask_hi[899:896]},
     {selectReadStageMask_hi[895:892]},
     {selectReadStageMask_hi[891:888]},
     {selectReadStageMask_hi[887:884]},
     {selectReadStageMask_hi[883:880]},
     {selectReadStageMask_hi[879:876]},
     {selectReadStageMask_hi[875:872]},
     {selectReadStageMask_hi[871:868]},
     {selectReadStageMask_hi[867:864]},
     {selectReadStageMask_hi[863:860]},
     {selectReadStageMask_hi[859:856]},
     {selectReadStageMask_hi[855:852]},
     {selectReadStageMask_hi[851:848]},
     {selectReadStageMask_hi[847:844]},
     {selectReadStageMask_hi[843:840]},
     {selectReadStageMask_hi[839:836]},
     {selectReadStageMask_hi[835:832]},
     {selectReadStageMask_hi[831:828]},
     {selectReadStageMask_hi[827:824]},
     {selectReadStageMask_hi[823:820]},
     {selectReadStageMask_hi[819:816]},
     {selectReadStageMask_hi[815:812]},
     {selectReadStageMask_hi[811:808]},
     {selectReadStageMask_hi[807:804]},
     {selectReadStageMask_hi[803:800]},
     {selectReadStageMask_hi[799:796]},
     {selectReadStageMask_hi[795:792]},
     {selectReadStageMask_hi[791:788]},
     {selectReadStageMask_hi[787:784]},
     {selectReadStageMask_hi[783:780]},
     {selectReadStageMask_hi[779:776]},
     {selectReadStageMask_hi[775:772]},
     {selectReadStageMask_hi[771:768]},
     {selectReadStageMask_hi[767:764]},
     {selectReadStageMask_hi[763:760]},
     {selectReadStageMask_hi[759:756]},
     {selectReadStageMask_hi[755:752]},
     {selectReadStageMask_hi[751:748]},
     {selectReadStageMask_hi[747:744]},
     {selectReadStageMask_hi[743:740]},
     {selectReadStageMask_hi[739:736]},
     {selectReadStageMask_hi[735:732]},
     {selectReadStageMask_hi[731:728]},
     {selectReadStageMask_hi[727:724]},
     {selectReadStageMask_hi[723:720]},
     {selectReadStageMask_hi[719:716]},
     {selectReadStageMask_hi[715:712]},
     {selectReadStageMask_hi[711:708]},
     {selectReadStageMask_hi[707:704]},
     {selectReadStageMask_hi[703:700]},
     {selectReadStageMask_hi[699:696]},
     {selectReadStageMask_hi[695:692]},
     {selectReadStageMask_hi[691:688]},
     {selectReadStageMask_hi[687:684]},
     {selectReadStageMask_hi[683:680]},
     {selectReadStageMask_hi[679:676]},
     {selectReadStageMask_hi[675:672]},
     {selectReadStageMask_hi[671:668]},
     {selectReadStageMask_hi[667:664]},
     {selectReadStageMask_hi[663:660]},
     {selectReadStageMask_hi[659:656]},
     {selectReadStageMask_hi[655:652]},
     {selectReadStageMask_hi[651:648]},
     {selectReadStageMask_hi[647:644]},
     {selectReadStageMask_hi[643:640]},
     {selectReadStageMask_hi[639:636]},
     {selectReadStageMask_hi[635:632]},
     {selectReadStageMask_hi[631:628]},
     {selectReadStageMask_hi[627:624]},
     {selectReadStageMask_hi[623:620]},
     {selectReadStageMask_hi[619:616]},
     {selectReadStageMask_hi[615:612]},
     {selectReadStageMask_hi[611:608]},
     {selectReadStageMask_hi[607:604]},
     {selectReadStageMask_hi[603:600]},
     {selectReadStageMask_hi[599:596]},
     {selectReadStageMask_hi[595:592]},
     {selectReadStageMask_hi[591:588]},
     {selectReadStageMask_hi[587:584]},
     {selectReadStageMask_hi[583:580]},
     {selectReadStageMask_hi[579:576]},
     {selectReadStageMask_hi[575:572]},
     {selectReadStageMask_hi[571:568]},
     {selectReadStageMask_hi[567:564]},
     {selectReadStageMask_hi[563:560]},
     {selectReadStageMask_hi[559:556]},
     {selectReadStageMask_hi[555:552]},
     {selectReadStageMask_hi[551:548]},
     {selectReadStageMask_hi[547:544]},
     {selectReadStageMask_hi[543:540]},
     {selectReadStageMask_hi[539:536]},
     {selectReadStageMask_hi[535:532]},
     {selectReadStageMask_hi[531:528]},
     {selectReadStageMask_hi[527:524]},
     {selectReadStageMask_hi[523:520]},
     {selectReadStageMask_hi[519:516]},
     {selectReadStageMask_hi[515:512]},
     {selectReadStageMask_hi[511:508]},
     {selectReadStageMask_hi[507:504]},
     {selectReadStageMask_hi[503:500]},
     {selectReadStageMask_hi[499:496]},
     {selectReadStageMask_hi[495:492]},
     {selectReadStageMask_hi[491:488]},
     {selectReadStageMask_hi[487:484]},
     {selectReadStageMask_hi[483:480]},
     {selectReadStageMask_hi[479:476]},
     {selectReadStageMask_hi[475:472]},
     {selectReadStageMask_hi[471:468]},
     {selectReadStageMask_hi[467:464]},
     {selectReadStageMask_hi[463:460]},
     {selectReadStageMask_hi[459:456]},
     {selectReadStageMask_hi[455:452]},
     {selectReadStageMask_hi[451:448]},
     {selectReadStageMask_hi[447:444]},
     {selectReadStageMask_hi[443:440]},
     {selectReadStageMask_hi[439:436]},
     {selectReadStageMask_hi[435:432]},
     {selectReadStageMask_hi[431:428]},
     {selectReadStageMask_hi[427:424]},
     {selectReadStageMask_hi[423:420]},
     {selectReadStageMask_hi[419:416]},
     {selectReadStageMask_hi[415:412]},
     {selectReadStageMask_hi[411:408]},
     {selectReadStageMask_hi[407:404]},
     {selectReadStageMask_hi[403:400]},
     {selectReadStageMask_hi[399:396]},
     {selectReadStageMask_hi[395:392]},
     {selectReadStageMask_hi[391:388]},
     {selectReadStageMask_hi[387:384]},
     {selectReadStageMask_hi[383:380]},
     {selectReadStageMask_hi[379:376]},
     {selectReadStageMask_hi[375:372]},
     {selectReadStageMask_hi[371:368]},
     {selectReadStageMask_hi[367:364]},
     {selectReadStageMask_hi[363:360]},
     {selectReadStageMask_hi[359:356]},
     {selectReadStageMask_hi[355:352]},
     {selectReadStageMask_hi[351:348]},
     {selectReadStageMask_hi[347:344]},
     {selectReadStageMask_hi[343:340]},
     {selectReadStageMask_hi[339:336]},
     {selectReadStageMask_hi[335:332]},
     {selectReadStageMask_hi[331:328]},
     {selectReadStageMask_hi[327:324]},
     {selectReadStageMask_hi[323:320]},
     {selectReadStageMask_hi[319:316]},
     {selectReadStageMask_hi[315:312]},
     {selectReadStageMask_hi[311:308]},
     {selectReadStageMask_hi[307:304]},
     {selectReadStageMask_hi[303:300]},
     {selectReadStageMask_hi[299:296]},
     {selectReadStageMask_hi[295:292]},
     {selectReadStageMask_hi[291:288]},
     {selectReadStageMask_hi[287:284]},
     {selectReadStageMask_hi[283:280]},
     {selectReadStageMask_hi[279:276]},
     {selectReadStageMask_hi[275:272]},
     {selectReadStageMask_hi[271:268]},
     {selectReadStageMask_hi[267:264]},
     {selectReadStageMask_hi[263:260]},
     {selectReadStageMask_hi[259:256]},
     {selectReadStageMask_hi[255:252]},
     {selectReadStageMask_hi[251:248]},
     {selectReadStageMask_hi[247:244]},
     {selectReadStageMask_hi[243:240]},
     {selectReadStageMask_hi[239:236]},
     {selectReadStageMask_hi[235:232]},
     {selectReadStageMask_hi[231:228]},
     {selectReadStageMask_hi[227:224]},
     {selectReadStageMask_hi[223:220]},
     {selectReadStageMask_hi[219:216]},
     {selectReadStageMask_hi[215:212]},
     {selectReadStageMask_hi[211:208]},
     {selectReadStageMask_hi[207:204]},
     {selectReadStageMask_hi[203:200]},
     {selectReadStageMask_hi[199:196]},
     {selectReadStageMask_hi[195:192]},
     {selectReadStageMask_hi[191:188]},
     {selectReadStageMask_hi[187:184]},
     {selectReadStageMask_hi[183:180]},
     {selectReadStageMask_hi[179:176]},
     {selectReadStageMask_hi[175:172]},
     {selectReadStageMask_hi[171:168]},
     {selectReadStageMask_hi[167:164]},
     {selectReadStageMask_hi[163:160]},
     {selectReadStageMask_hi[159:156]},
     {selectReadStageMask_hi[155:152]},
     {selectReadStageMask_hi[151:148]},
     {selectReadStageMask_hi[147:144]},
     {selectReadStageMask_hi[143:140]},
     {selectReadStageMask_hi[139:136]},
     {selectReadStageMask_hi[135:132]},
     {selectReadStageMask_hi[131:128]},
     {selectReadStageMask_hi[127:124]},
     {selectReadStageMask_hi[123:120]},
     {selectReadStageMask_hi[119:116]},
     {selectReadStageMask_hi[115:112]},
     {selectReadStageMask_hi[111:108]},
     {selectReadStageMask_hi[107:104]},
     {selectReadStageMask_hi[103:100]},
     {selectReadStageMask_hi[99:96]},
     {selectReadStageMask_hi[95:92]},
     {selectReadStageMask_hi[91:88]},
     {selectReadStageMask_hi[87:84]},
     {selectReadStageMask_hi[83:80]},
     {selectReadStageMask_hi[79:76]},
     {selectReadStageMask_hi[75:72]},
     {selectReadStageMask_hi[71:68]},
     {selectReadStageMask_hi[67:64]},
     {selectReadStageMask_hi[63:60]},
     {selectReadStageMask_hi[59:56]},
     {selectReadStageMask_hi[55:52]},
     {selectReadStageMask_hi[51:48]},
     {selectReadStageMask_hi[47:44]},
     {selectReadStageMask_hi[43:40]},
     {selectReadStageMask_hi[39:36]},
     {selectReadStageMask_hi[35:32]},
     {selectReadStageMask_hi[31:28]},
     {selectReadStageMask_hi[27:24]},
     {selectReadStageMask_hi[23:20]},
     {selectReadStageMask_hi[19:16]},
     {selectReadStageMask_hi[15:12]},
     {selectReadStageMask_hi[11:8]},
     {selectReadStageMask_hi[7:4]},
     {selectReadStageMask_hi[3:0]},
     {selectReadStageMask_lo[4095:4092]},
     {selectReadStageMask_lo[4091:4088]},
     {selectReadStageMask_lo[4087:4084]},
     {selectReadStageMask_lo[4083:4080]},
     {selectReadStageMask_lo[4079:4076]},
     {selectReadStageMask_lo[4075:4072]},
     {selectReadStageMask_lo[4071:4068]},
     {selectReadStageMask_lo[4067:4064]},
     {selectReadStageMask_lo[4063:4060]},
     {selectReadStageMask_lo[4059:4056]},
     {selectReadStageMask_lo[4055:4052]},
     {selectReadStageMask_lo[4051:4048]},
     {selectReadStageMask_lo[4047:4044]},
     {selectReadStageMask_lo[4043:4040]},
     {selectReadStageMask_lo[4039:4036]},
     {selectReadStageMask_lo[4035:4032]},
     {selectReadStageMask_lo[4031:4028]},
     {selectReadStageMask_lo[4027:4024]},
     {selectReadStageMask_lo[4023:4020]},
     {selectReadStageMask_lo[4019:4016]},
     {selectReadStageMask_lo[4015:4012]},
     {selectReadStageMask_lo[4011:4008]},
     {selectReadStageMask_lo[4007:4004]},
     {selectReadStageMask_lo[4003:4000]},
     {selectReadStageMask_lo[3999:3996]},
     {selectReadStageMask_lo[3995:3992]},
     {selectReadStageMask_lo[3991:3988]},
     {selectReadStageMask_lo[3987:3984]},
     {selectReadStageMask_lo[3983:3980]},
     {selectReadStageMask_lo[3979:3976]},
     {selectReadStageMask_lo[3975:3972]},
     {selectReadStageMask_lo[3971:3968]},
     {selectReadStageMask_lo[3967:3964]},
     {selectReadStageMask_lo[3963:3960]},
     {selectReadStageMask_lo[3959:3956]},
     {selectReadStageMask_lo[3955:3952]},
     {selectReadStageMask_lo[3951:3948]},
     {selectReadStageMask_lo[3947:3944]},
     {selectReadStageMask_lo[3943:3940]},
     {selectReadStageMask_lo[3939:3936]},
     {selectReadStageMask_lo[3935:3932]},
     {selectReadStageMask_lo[3931:3928]},
     {selectReadStageMask_lo[3927:3924]},
     {selectReadStageMask_lo[3923:3920]},
     {selectReadStageMask_lo[3919:3916]},
     {selectReadStageMask_lo[3915:3912]},
     {selectReadStageMask_lo[3911:3908]},
     {selectReadStageMask_lo[3907:3904]},
     {selectReadStageMask_lo[3903:3900]},
     {selectReadStageMask_lo[3899:3896]},
     {selectReadStageMask_lo[3895:3892]},
     {selectReadStageMask_lo[3891:3888]},
     {selectReadStageMask_lo[3887:3884]},
     {selectReadStageMask_lo[3883:3880]},
     {selectReadStageMask_lo[3879:3876]},
     {selectReadStageMask_lo[3875:3872]},
     {selectReadStageMask_lo[3871:3868]},
     {selectReadStageMask_lo[3867:3864]},
     {selectReadStageMask_lo[3863:3860]},
     {selectReadStageMask_lo[3859:3856]},
     {selectReadStageMask_lo[3855:3852]},
     {selectReadStageMask_lo[3851:3848]},
     {selectReadStageMask_lo[3847:3844]},
     {selectReadStageMask_lo[3843:3840]},
     {selectReadStageMask_lo[3839:3836]},
     {selectReadStageMask_lo[3835:3832]},
     {selectReadStageMask_lo[3831:3828]},
     {selectReadStageMask_lo[3827:3824]},
     {selectReadStageMask_lo[3823:3820]},
     {selectReadStageMask_lo[3819:3816]},
     {selectReadStageMask_lo[3815:3812]},
     {selectReadStageMask_lo[3811:3808]},
     {selectReadStageMask_lo[3807:3804]},
     {selectReadStageMask_lo[3803:3800]},
     {selectReadStageMask_lo[3799:3796]},
     {selectReadStageMask_lo[3795:3792]},
     {selectReadStageMask_lo[3791:3788]},
     {selectReadStageMask_lo[3787:3784]},
     {selectReadStageMask_lo[3783:3780]},
     {selectReadStageMask_lo[3779:3776]},
     {selectReadStageMask_lo[3775:3772]},
     {selectReadStageMask_lo[3771:3768]},
     {selectReadStageMask_lo[3767:3764]},
     {selectReadStageMask_lo[3763:3760]},
     {selectReadStageMask_lo[3759:3756]},
     {selectReadStageMask_lo[3755:3752]},
     {selectReadStageMask_lo[3751:3748]},
     {selectReadStageMask_lo[3747:3744]},
     {selectReadStageMask_lo[3743:3740]},
     {selectReadStageMask_lo[3739:3736]},
     {selectReadStageMask_lo[3735:3732]},
     {selectReadStageMask_lo[3731:3728]},
     {selectReadStageMask_lo[3727:3724]},
     {selectReadStageMask_lo[3723:3720]},
     {selectReadStageMask_lo[3719:3716]},
     {selectReadStageMask_lo[3715:3712]},
     {selectReadStageMask_lo[3711:3708]},
     {selectReadStageMask_lo[3707:3704]},
     {selectReadStageMask_lo[3703:3700]},
     {selectReadStageMask_lo[3699:3696]},
     {selectReadStageMask_lo[3695:3692]},
     {selectReadStageMask_lo[3691:3688]},
     {selectReadStageMask_lo[3687:3684]},
     {selectReadStageMask_lo[3683:3680]},
     {selectReadStageMask_lo[3679:3676]},
     {selectReadStageMask_lo[3675:3672]},
     {selectReadStageMask_lo[3671:3668]},
     {selectReadStageMask_lo[3667:3664]},
     {selectReadStageMask_lo[3663:3660]},
     {selectReadStageMask_lo[3659:3656]},
     {selectReadStageMask_lo[3655:3652]},
     {selectReadStageMask_lo[3651:3648]},
     {selectReadStageMask_lo[3647:3644]},
     {selectReadStageMask_lo[3643:3640]},
     {selectReadStageMask_lo[3639:3636]},
     {selectReadStageMask_lo[3635:3632]},
     {selectReadStageMask_lo[3631:3628]},
     {selectReadStageMask_lo[3627:3624]},
     {selectReadStageMask_lo[3623:3620]},
     {selectReadStageMask_lo[3619:3616]},
     {selectReadStageMask_lo[3615:3612]},
     {selectReadStageMask_lo[3611:3608]},
     {selectReadStageMask_lo[3607:3604]},
     {selectReadStageMask_lo[3603:3600]},
     {selectReadStageMask_lo[3599:3596]},
     {selectReadStageMask_lo[3595:3592]},
     {selectReadStageMask_lo[3591:3588]},
     {selectReadStageMask_lo[3587:3584]},
     {selectReadStageMask_lo[3583:3580]},
     {selectReadStageMask_lo[3579:3576]},
     {selectReadStageMask_lo[3575:3572]},
     {selectReadStageMask_lo[3571:3568]},
     {selectReadStageMask_lo[3567:3564]},
     {selectReadStageMask_lo[3563:3560]},
     {selectReadStageMask_lo[3559:3556]},
     {selectReadStageMask_lo[3555:3552]},
     {selectReadStageMask_lo[3551:3548]},
     {selectReadStageMask_lo[3547:3544]},
     {selectReadStageMask_lo[3543:3540]},
     {selectReadStageMask_lo[3539:3536]},
     {selectReadStageMask_lo[3535:3532]},
     {selectReadStageMask_lo[3531:3528]},
     {selectReadStageMask_lo[3527:3524]},
     {selectReadStageMask_lo[3523:3520]},
     {selectReadStageMask_lo[3519:3516]},
     {selectReadStageMask_lo[3515:3512]},
     {selectReadStageMask_lo[3511:3508]},
     {selectReadStageMask_lo[3507:3504]},
     {selectReadStageMask_lo[3503:3500]},
     {selectReadStageMask_lo[3499:3496]},
     {selectReadStageMask_lo[3495:3492]},
     {selectReadStageMask_lo[3491:3488]},
     {selectReadStageMask_lo[3487:3484]},
     {selectReadStageMask_lo[3483:3480]},
     {selectReadStageMask_lo[3479:3476]},
     {selectReadStageMask_lo[3475:3472]},
     {selectReadStageMask_lo[3471:3468]},
     {selectReadStageMask_lo[3467:3464]},
     {selectReadStageMask_lo[3463:3460]},
     {selectReadStageMask_lo[3459:3456]},
     {selectReadStageMask_lo[3455:3452]},
     {selectReadStageMask_lo[3451:3448]},
     {selectReadStageMask_lo[3447:3444]},
     {selectReadStageMask_lo[3443:3440]},
     {selectReadStageMask_lo[3439:3436]},
     {selectReadStageMask_lo[3435:3432]},
     {selectReadStageMask_lo[3431:3428]},
     {selectReadStageMask_lo[3427:3424]},
     {selectReadStageMask_lo[3423:3420]},
     {selectReadStageMask_lo[3419:3416]},
     {selectReadStageMask_lo[3415:3412]},
     {selectReadStageMask_lo[3411:3408]},
     {selectReadStageMask_lo[3407:3404]},
     {selectReadStageMask_lo[3403:3400]},
     {selectReadStageMask_lo[3399:3396]},
     {selectReadStageMask_lo[3395:3392]},
     {selectReadStageMask_lo[3391:3388]},
     {selectReadStageMask_lo[3387:3384]},
     {selectReadStageMask_lo[3383:3380]},
     {selectReadStageMask_lo[3379:3376]},
     {selectReadStageMask_lo[3375:3372]},
     {selectReadStageMask_lo[3371:3368]},
     {selectReadStageMask_lo[3367:3364]},
     {selectReadStageMask_lo[3363:3360]},
     {selectReadStageMask_lo[3359:3356]},
     {selectReadStageMask_lo[3355:3352]},
     {selectReadStageMask_lo[3351:3348]},
     {selectReadStageMask_lo[3347:3344]},
     {selectReadStageMask_lo[3343:3340]},
     {selectReadStageMask_lo[3339:3336]},
     {selectReadStageMask_lo[3335:3332]},
     {selectReadStageMask_lo[3331:3328]},
     {selectReadStageMask_lo[3327:3324]},
     {selectReadStageMask_lo[3323:3320]},
     {selectReadStageMask_lo[3319:3316]},
     {selectReadStageMask_lo[3315:3312]},
     {selectReadStageMask_lo[3311:3308]},
     {selectReadStageMask_lo[3307:3304]},
     {selectReadStageMask_lo[3303:3300]},
     {selectReadStageMask_lo[3299:3296]},
     {selectReadStageMask_lo[3295:3292]},
     {selectReadStageMask_lo[3291:3288]},
     {selectReadStageMask_lo[3287:3284]},
     {selectReadStageMask_lo[3283:3280]},
     {selectReadStageMask_lo[3279:3276]},
     {selectReadStageMask_lo[3275:3272]},
     {selectReadStageMask_lo[3271:3268]},
     {selectReadStageMask_lo[3267:3264]},
     {selectReadStageMask_lo[3263:3260]},
     {selectReadStageMask_lo[3259:3256]},
     {selectReadStageMask_lo[3255:3252]},
     {selectReadStageMask_lo[3251:3248]},
     {selectReadStageMask_lo[3247:3244]},
     {selectReadStageMask_lo[3243:3240]},
     {selectReadStageMask_lo[3239:3236]},
     {selectReadStageMask_lo[3235:3232]},
     {selectReadStageMask_lo[3231:3228]},
     {selectReadStageMask_lo[3227:3224]},
     {selectReadStageMask_lo[3223:3220]},
     {selectReadStageMask_lo[3219:3216]},
     {selectReadStageMask_lo[3215:3212]},
     {selectReadStageMask_lo[3211:3208]},
     {selectReadStageMask_lo[3207:3204]},
     {selectReadStageMask_lo[3203:3200]},
     {selectReadStageMask_lo[3199:3196]},
     {selectReadStageMask_lo[3195:3192]},
     {selectReadStageMask_lo[3191:3188]},
     {selectReadStageMask_lo[3187:3184]},
     {selectReadStageMask_lo[3183:3180]},
     {selectReadStageMask_lo[3179:3176]},
     {selectReadStageMask_lo[3175:3172]},
     {selectReadStageMask_lo[3171:3168]},
     {selectReadStageMask_lo[3167:3164]},
     {selectReadStageMask_lo[3163:3160]},
     {selectReadStageMask_lo[3159:3156]},
     {selectReadStageMask_lo[3155:3152]},
     {selectReadStageMask_lo[3151:3148]},
     {selectReadStageMask_lo[3147:3144]},
     {selectReadStageMask_lo[3143:3140]},
     {selectReadStageMask_lo[3139:3136]},
     {selectReadStageMask_lo[3135:3132]},
     {selectReadStageMask_lo[3131:3128]},
     {selectReadStageMask_lo[3127:3124]},
     {selectReadStageMask_lo[3123:3120]},
     {selectReadStageMask_lo[3119:3116]},
     {selectReadStageMask_lo[3115:3112]},
     {selectReadStageMask_lo[3111:3108]},
     {selectReadStageMask_lo[3107:3104]},
     {selectReadStageMask_lo[3103:3100]},
     {selectReadStageMask_lo[3099:3096]},
     {selectReadStageMask_lo[3095:3092]},
     {selectReadStageMask_lo[3091:3088]},
     {selectReadStageMask_lo[3087:3084]},
     {selectReadStageMask_lo[3083:3080]},
     {selectReadStageMask_lo[3079:3076]},
     {selectReadStageMask_lo[3075:3072]},
     {selectReadStageMask_lo[3071:3068]},
     {selectReadStageMask_lo[3067:3064]},
     {selectReadStageMask_lo[3063:3060]},
     {selectReadStageMask_lo[3059:3056]},
     {selectReadStageMask_lo[3055:3052]},
     {selectReadStageMask_lo[3051:3048]},
     {selectReadStageMask_lo[3047:3044]},
     {selectReadStageMask_lo[3043:3040]},
     {selectReadStageMask_lo[3039:3036]},
     {selectReadStageMask_lo[3035:3032]},
     {selectReadStageMask_lo[3031:3028]},
     {selectReadStageMask_lo[3027:3024]},
     {selectReadStageMask_lo[3023:3020]},
     {selectReadStageMask_lo[3019:3016]},
     {selectReadStageMask_lo[3015:3012]},
     {selectReadStageMask_lo[3011:3008]},
     {selectReadStageMask_lo[3007:3004]},
     {selectReadStageMask_lo[3003:3000]},
     {selectReadStageMask_lo[2999:2996]},
     {selectReadStageMask_lo[2995:2992]},
     {selectReadStageMask_lo[2991:2988]},
     {selectReadStageMask_lo[2987:2984]},
     {selectReadStageMask_lo[2983:2980]},
     {selectReadStageMask_lo[2979:2976]},
     {selectReadStageMask_lo[2975:2972]},
     {selectReadStageMask_lo[2971:2968]},
     {selectReadStageMask_lo[2967:2964]},
     {selectReadStageMask_lo[2963:2960]},
     {selectReadStageMask_lo[2959:2956]},
     {selectReadStageMask_lo[2955:2952]},
     {selectReadStageMask_lo[2951:2948]},
     {selectReadStageMask_lo[2947:2944]},
     {selectReadStageMask_lo[2943:2940]},
     {selectReadStageMask_lo[2939:2936]},
     {selectReadStageMask_lo[2935:2932]},
     {selectReadStageMask_lo[2931:2928]},
     {selectReadStageMask_lo[2927:2924]},
     {selectReadStageMask_lo[2923:2920]},
     {selectReadStageMask_lo[2919:2916]},
     {selectReadStageMask_lo[2915:2912]},
     {selectReadStageMask_lo[2911:2908]},
     {selectReadStageMask_lo[2907:2904]},
     {selectReadStageMask_lo[2903:2900]},
     {selectReadStageMask_lo[2899:2896]},
     {selectReadStageMask_lo[2895:2892]},
     {selectReadStageMask_lo[2891:2888]},
     {selectReadStageMask_lo[2887:2884]},
     {selectReadStageMask_lo[2883:2880]},
     {selectReadStageMask_lo[2879:2876]},
     {selectReadStageMask_lo[2875:2872]},
     {selectReadStageMask_lo[2871:2868]},
     {selectReadStageMask_lo[2867:2864]},
     {selectReadStageMask_lo[2863:2860]},
     {selectReadStageMask_lo[2859:2856]},
     {selectReadStageMask_lo[2855:2852]},
     {selectReadStageMask_lo[2851:2848]},
     {selectReadStageMask_lo[2847:2844]},
     {selectReadStageMask_lo[2843:2840]},
     {selectReadStageMask_lo[2839:2836]},
     {selectReadStageMask_lo[2835:2832]},
     {selectReadStageMask_lo[2831:2828]},
     {selectReadStageMask_lo[2827:2824]},
     {selectReadStageMask_lo[2823:2820]},
     {selectReadStageMask_lo[2819:2816]},
     {selectReadStageMask_lo[2815:2812]},
     {selectReadStageMask_lo[2811:2808]},
     {selectReadStageMask_lo[2807:2804]},
     {selectReadStageMask_lo[2803:2800]},
     {selectReadStageMask_lo[2799:2796]},
     {selectReadStageMask_lo[2795:2792]},
     {selectReadStageMask_lo[2791:2788]},
     {selectReadStageMask_lo[2787:2784]},
     {selectReadStageMask_lo[2783:2780]},
     {selectReadStageMask_lo[2779:2776]},
     {selectReadStageMask_lo[2775:2772]},
     {selectReadStageMask_lo[2771:2768]},
     {selectReadStageMask_lo[2767:2764]},
     {selectReadStageMask_lo[2763:2760]},
     {selectReadStageMask_lo[2759:2756]},
     {selectReadStageMask_lo[2755:2752]},
     {selectReadStageMask_lo[2751:2748]},
     {selectReadStageMask_lo[2747:2744]},
     {selectReadStageMask_lo[2743:2740]},
     {selectReadStageMask_lo[2739:2736]},
     {selectReadStageMask_lo[2735:2732]},
     {selectReadStageMask_lo[2731:2728]},
     {selectReadStageMask_lo[2727:2724]},
     {selectReadStageMask_lo[2723:2720]},
     {selectReadStageMask_lo[2719:2716]},
     {selectReadStageMask_lo[2715:2712]},
     {selectReadStageMask_lo[2711:2708]},
     {selectReadStageMask_lo[2707:2704]},
     {selectReadStageMask_lo[2703:2700]},
     {selectReadStageMask_lo[2699:2696]},
     {selectReadStageMask_lo[2695:2692]},
     {selectReadStageMask_lo[2691:2688]},
     {selectReadStageMask_lo[2687:2684]},
     {selectReadStageMask_lo[2683:2680]},
     {selectReadStageMask_lo[2679:2676]},
     {selectReadStageMask_lo[2675:2672]},
     {selectReadStageMask_lo[2671:2668]},
     {selectReadStageMask_lo[2667:2664]},
     {selectReadStageMask_lo[2663:2660]},
     {selectReadStageMask_lo[2659:2656]},
     {selectReadStageMask_lo[2655:2652]},
     {selectReadStageMask_lo[2651:2648]},
     {selectReadStageMask_lo[2647:2644]},
     {selectReadStageMask_lo[2643:2640]},
     {selectReadStageMask_lo[2639:2636]},
     {selectReadStageMask_lo[2635:2632]},
     {selectReadStageMask_lo[2631:2628]},
     {selectReadStageMask_lo[2627:2624]},
     {selectReadStageMask_lo[2623:2620]},
     {selectReadStageMask_lo[2619:2616]},
     {selectReadStageMask_lo[2615:2612]},
     {selectReadStageMask_lo[2611:2608]},
     {selectReadStageMask_lo[2607:2604]},
     {selectReadStageMask_lo[2603:2600]},
     {selectReadStageMask_lo[2599:2596]},
     {selectReadStageMask_lo[2595:2592]},
     {selectReadStageMask_lo[2591:2588]},
     {selectReadStageMask_lo[2587:2584]},
     {selectReadStageMask_lo[2583:2580]},
     {selectReadStageMask_lo[2579:2576]},
     {selectReadStageMask_lo[2575:2572]},
     {selectReadStageMask_lo[2571:2568]},
     {selectReadStageMask_lo[2567:2564]},
     {selectReadStageMask_lo[2563:2560]},
     {selectReadStageMask_lo[2559:2556]},
     {selectReadStageMask_lo[2555:2552]},
     {selectReadStageMask_lo[2551:2548]},
     {selectReadStageMask_lo[2547:2544]},
     {selectReadStageMask_lo[2543:2540]},
     {selectReadStageMask_lo[2539:2536]},
     {selectReadStageMask_lo[2535:2532]},
     {selectReadStageMask_lo[2531:2528]},
     {selectReadStageMask_lo[2527:2524]},
     {selectReadStageMask_lo[2523:2520]},
     {selectReadStageMask_lo[2519:2516]},
     {selectReadStageMask_lo[2515:2512]},
     {selectReadStageMask_lo[2511:2508]},
     {selectReadStageMask_lo[2507:2504]},
     {selectReadStageMask_lo[2503:2500]},
     {selectReadStageMask_lo[2499:2496]},
     {selectReadStageMask_lo[2495:2492]},
     {selectReadStageMask_lo[2491:2488]},
     {selectReadStageMask_lo[2487:2484]},
     {selectReadStageMask_lo[2483:2480]},
     {selectReadStageMask_lo[2479:2476]},
     {selectReadStageMask_lo[2475:2472]},
     {selectReadStageMask_lo[2471:2468]},
     {selectReadStageMask_lo[2467:2464]},
     {selectReadStageMask_lo[2463:2460]},
     {selectReadStageMask_lo[2459:2456]},
     {selectReadStageMask_lo[2455:2452]},
     {selectReadStageMask_lo[2451:2448]},
     {selectReadStageMask_lo[2447:2444]},
     {selectReadStageMask_lo[2443:2440]},
     {selectReadStageMask_lo[2439:2436]},
     {selectReadStageMask_lo[2435:2432]},
     {selectReadStageMask_lo[2431:2428]},
     {selectReadStageMask_lo[2427:2424]},
     {selectReadStageMask_lo[2423:2420]},
     {selectReadStageMask_lo[2419:2416]},
     {selectReadStageMask_lo[2415:2412]},
     {selectReadStageMask_lo[2411:2408]},
     {selectReadStageMask_lo[2407:2404]},
     {selectReadStageMask_lo[2403:2400]},
     {selectReadStageMask_lo[2399:2396]},
     {selectReadStageMask_lo[2395:2392]},
     {selectReadStageMask_lo[2391:2388]},
     {selectReadStageMask_lo[2387:2384]},
     {selectReadStageMask_lo[2383:2380]},
     {selectReadStageMask_lo[2379:2376]},
     {selectReadStageMask_lo[2375:2372]},
     {selectReadStageMask_lo[2371:2368]},
     {selectReadStageMask_lo[2367:2364]},
     {selectReadStageMask_lo[2363:2360]},
     {selectReadStageMask_lo[2359:2356]},
     {selectReadStageMask_lo[2355:2352]},
     {selectReadStageMask_lo[2351:2348]},
     {selectReadStageMask_lo[2347:2344]},
     {selectReadStageMask_lo[2343:2340]},
     {selectReadStageMask_lo[2339:2336]},
     {selectReadStageMask_lo[2335:2332]},
     {selectReadStageMask_lo[2331:2328]},
     {selectReadStageMask_lo[2327:2324]},
     {selectReadStageMask_lo[2323:2320]},
     {selectReadStageMask_lo[2319:2316]},
     {selectReadStageMask_lo[2315:2312]},
     {selectReadStageMask_lo[2311:2308]},
     {selectReadStageMask_lo[2307:2304]},
     {selectReadStageMask_lo[2303:2300]},
     {selectReadStageMask_lo[2299:2296]},
     {selectReadStageMask_lo[2295:2292]},
     {selectReadStageMask_lo[2291:2288]},
     {selectReadStageMask_lo[2287:2284]},
     {selectReadStageMask_lo[2283:2280]},
     {selectReadStageMask_lo[2279:2276]},
     {selectReadStageMask_lo[2275:2272]},
     {selectReadStageMask_lo[2271:2268]},
     {selectReadStageMask_lo[2267:2264]},
     {selectReadStageMask_lo[2263:2260]},
     {selectReadStageMask_lo[2259:2256]},
     {selectReadStageMask_lo[2255:2252]},
     {selectReadStageMask_lo[2251:2248]},
     {selectReadStageMask_lo[2247:2244]},
     {selectReadStageMask_lo[2243:2240]},
     {selectReadStageMask_lo[2239:2236]},
     {selectReadStageMask_lo[2235:2232]},
     {selectReadStageMask_lo[2231:2228]},
     {selectReadStageMask_lo[2227:2224]},
     {selectReadStageMask_lo[2223:2220]},
     {selectReadStageMask_lo[2219:2216]},
     {selectReadStageMask_lo[2215:2212]},
     {selectReadStageMask_lo[2211:2208]},
     {selectReadStageMask_lo[2207:2204]},
     {selectReadStageMask_lo[2203:2200]},
     {selectReadStageMask_lo[2199:2196]},
     {selectReadStageMask_lo[2195:2192]},
     {selectReadStageMask_lo[2191:2188]},
     {selectReadStageMask_lo[2187:2184]},
     {selectReadStageMask_lo[2183:2180]},
     {selectReadStageMask_lo[2179:2176]},
     {selectReadStageMask_lo[2175:2172]},
     {selectReadStageMask_lo[2171:2168]},
     {selectReadStageMask_lo[2167:2164]},
     {selectReadStageMask_lo[2163:2160]},
     {selectReadStageMask_lo[2159:2156]},
     {selectReadStageMask_lo[2155:2152]},
     {selectReadStageMask_lo[2151:2148]},
     {selectReadStageMask_lo[2147:2144]},
     {selectReadStageMask_lo[2143:2140]},
     {selectReadStageMask_lo[2139:2136]},
     {selectReadStageMask_lo[2135:2132]},
     {selectReadStageMask_lo[2131:2128]},
     {selectReadStageMask_lo[2127:2124]},
     {selectReadStageMask_lo[2123:2120]},
     {selectReadStageMask_lo[2119:2116]},
     {selectReadStageMask_lo[2115:2112]},
     {selectReadStageMask_lo[2111:2108]},
     {selectReadStageMask_lo[2107:2104]},
     {selectReadStageMask_lo[2103:2100]},
     {selectReadStageMask_lo[2099:2096]},
     {selectReadStageMask_lo[2095:2092]},
     {selectReadStageMask_lo[2091:2088]},
     {selectReadStageMask_lo[2087:2084]},
     {selectReadStageMask_lo[2083:2080]},
     {selectReadStageMask_lo[2079:2076]},
     {selectReadStageMask_lo[2075:2072]},
     {selectReadStageMask_lo[2071:2068]},
     {selectReadStageMask_lo[2067:2064]},
     {selectReadStageMask_lo[2063:2060]},
     {selectReadStageMask_lo[2059:2056]},
     {selectReadStageMask_lo[2055:2052]},
     {selectReadStageMask_lo[2051:2048]},
     {selectReadStageMask_lo[2047:2044]},
     {selectReadStageMask_lo[2043:2040]},
     {selectReadStageMask_lo[2039:2036]},
     {selectReadStageMask_lo[2035:2032]},
     {selectReadStageMask_lo[2031:2028]},
     {selectReadStageMask_lo[2027:2024]},
     {selectReadStageMask_lo[2023:2020]},
     {selectReadStageMask_lo[2019:2016]},
     {selectReadStageMask_lo[2015:2012]},
     {selectReadStageMask_lo[2011:2008]},
     {selectReadStageMask_lo[2007:2004]},
     {selectReadStageMask_lo[2003:2000]},
     {selectReadStageMask_lo[1999:1996]},
     {selectReadStageMask_lo[1995:1992]},
     {selectReadStageMask_lo[1991:1988]},
     {selectReadStageMask_lo[1987:1984]},
     {selectReadStageMask_lo[1983:1980]},
     {selectReadStageMask_lo[1979:1976]},
     {selectReadStageMask_lo[1975:1972]},
     {selectReadStageMask_lo[1971:1968]},
     {selectReadStageMask_lo[1967:1964]},
     {selectReadStageMask_lo[1963:1960]},
     {selectReadStageMask_lo[1959:1956]},
     {selectReadStageMask_lo[1955:1952]},
     {selectReadStageMask_lo[1951:1948]},
     {selectReadStageMask_lo[1947:1944]},
     {selectReadStageMask_lo[1943:1940]},
     {selectReadStageMask_lo[1939:1936]},
     {selectReadStageMask_lo[1935:1932]},
     {selectReadStageMask_lo[1931:1928]},
     {selectReadStageMask_lo[1927:1924]},
     {selectReadStageMask_lo[1923:1920]},
     {selectReadStageMask_lo[1919:1916]},
     {selectReadStageMask_lo[1915:1912]},
     {selectReadStageMask_lo[1911:1908]},
     {selectReadStageMask_lo[1907:1904]},
     {selectReadStageMask_lo[1903:1900]},
     {selectReadStageMask_lo[1899:1896]},
     {selectReadStageMask_lo[1895:1892]},
     {selectReadStageMask_lo[1891:1888]},
     {selectReadStageMask_lo[1887:1884]},
     {selectReadStageMask_lo[1883:1880]},
     {selectReadStageMask_lo[1879:1876]},
     {selectReadStageMask_lo[1875:1872]},
     {selectReadStageMask_lo[1871:1868]},
     {selectReadStageMask_lo[1867:1864]},
     {selectReadStageMask_lo[1863:1860]},
     {selectReadStageMask_lo[1859:1856]},
     {selectReadStageMask_lo[1855:1852]},
     {selectReadStageMask_lo[1851:1848]},
     {selectReadStageMask_lo[1847:1844]},
     {selectReadStageMask_lo[1843:1840]},
     {selectReadStageMask_lo[1839:1836]},
     {selectReadStageMask_lo[1835:1832]},
     {selectReadStageMask_lo[1831:1828]},
     {selectReadStageMask_lo[1827:1824]},
     {selectReadStageMask_lo[1823:1820]},
     {selectReadStageMask_lo[1819:1816]},
     {selectReadStageMask_lo[1815:1812]},
     {selectReadStageMask_lo[1811:1808]},
     {selectReadStageMask_lo[1807:1804]},
     {selectReadStageMask_lo[1803:1800]},
     {selectReadStageMask_lo[1799:1796]},
     {selectReadStageMask_lo[1795:1792]},
     {selectReadStageMask_lo[1791:1788]},
     {selectReadStageMask_lo[1787:1784]},
     {selectReadStageMask_lo[1783:1780]},
     {selectReadStageMask_lo[1779:1776]},
     {selectReadStageMask_lo[1775:1772]},
     {selectReadStageMask_lo[1771:1768]},
     {selectReadStageMask_lo[1767:1764]},
     {selectReadStageMask_lo[1763:1760]},
     {selectReadStageMask_lo[1759:1756]},
     {selectReadStageMask_lo[1755:1752]},
     {selectReadStageMask_lo[1751:1748]},
     {selectReadStageMask_lo[1747:1744]},
     {selectReadStageMask_lo[1743:1740]},
     {selectReadStageMask_lo[1739:1736]},
     {selectReadStageMask_lo[1735:1732]},
     {selectReadStageMask_lo[1731:1728]},
     {selectReadStageMask_lo[1727:1724]},
     {selectReadStageMask_lo[1723:1720]},
     {selectReadStageMask_lo[1719:1716]},
     {selectReadStageMask_lo[1715:1712]},
     {selectReadStageMask_lo[1711:1708]},
     {selectReadStageMask_lo[1707:1704]},
     {selectReadStageMask_lo[1703:1700]},
     {selectReadStageMask_lo[1699:1696]},
     {selectReadStageMask_lo[1695:1692]},
     {selectReadStageMask_lo[1691:1688]},
     {selectReadStageMask_lo[1687:1684]},
     {selectReadStageMask_lo[1683:1680]},
     {selectReadStageMask_lo[1679:1676]},
     {selectReadStageMask_lo[1675:1672]},
     {selectReadStageMask_lo[1671:1668]},
     {selectReadStageMask_lo[1667:1664]},
     {selectReadStageMask_lo[1663:1660]},
     {selectReadStageMask_lo[1659:1656]},
     {selectReadStageMask_lo[1655:1652]},
     {selectReadStageMask_lo[1651:1648]},
     {selectReadStageMask_lo[1647:1644]},
     {selectReadStageMask_lo[1643:1640]},
     {selectReadStageMask_lo[1639:1636]},
     {selectReadStageMask_lo[1635:1632]},
     {selectReadStageMask_lo[1631:1628]},
     {selectReadStageMask_lo[1627:1624]},
     {selectReadStageMask_lo[1623:1620]},
     {selectReadStageMask_lo[1619:1616]},
     {selectReadStageMask_lo[1615:1612]},
     {selectReadStageMask_lo[1611:1608]},
     {selectReadStageMask_lo[1607:1604]},
     {selectReadStageMask_lo[1603:1600]},
     {selectReadStageMask_lo[1599:1596]},
     {selectReadStageMask_lo[1595:1592]},
     {selectReadStageMask_lo[1591:1588]},
     {selectReadStageMask_lo[1587:1584]},
     {selectReadStageMask_lo[1583:1580]},
     {selectReadStageMask_lo[1579:1576]},
     {selectReadStageMask_lo[1575:1572]},
     {selectReadStageMask_lo[1571:1568]},
     {selectReadStageMask_lo[1567:1564]},
     {selectReadStageMask_lo[1563:1560]},
     {selectReadStageMask_lo[1559:1556]},
     {selectReadStageMask_lo[1555:1552]},
     {selectReadStageMask_lo[1551:1548]},
     {selectReadStageMask_lo[1547:1544]},
     {selectReadStageMask_lo[1543:1540]},
     {selectReadStageMask_lo[1539:1536]},
     {selectReadStageMask_lo[1535:1532]},
     {selectReadStageMask_lo[1531:1528]},
     {selectReadStageMask_lo[1527:1524]},
     {selectReadStageMask_lo[1523:1520]},
     {selectReadStageMask_lo[1519:1516]},
     {selectReadStageMask_lo[1515:1512]},
     {selectReadStageMask_lo[1511:1508]},
     {selectReadStageMask_lo[1507:1504]},
     {selectReadStageMask_lo[1503:1500]},
     {selectReadStageMask_lo[1499:1496]},
     {selectReadStageMask_lo[1495:1492]},
     {selectReadStageMask_lo[1491:1488]},
     {selectReadStageMask_lo[1487:1484]},
     {selectReadStageMask_lo[1483:1480]},
     {selectReadStageMask_lo[1479:1476]},
     {selectReadStageMask_lo[1475:1472]},
     {selectReadStageMask_lo[1471:1468]},
     {selectReadStageMask_lo[1467:1464]},
     {selectReadStageMask_lo[1463:1460]},
     {selectReadStageMask_lo[1459:1456]},
     {selectReadStageMask_lo[1455:1452]},
     {selectReadStageMask_lo[1451:1448]},
     {selectReadStageMask_lo[1447:1444]},
     {selectReadStageMask_lo[1443:1440]},
     {selectReadStageMask_lo[1439:1436]},
     {selectReadStageMask_lo[1435:1432]},
     {selectReadStageMask_lo[1431:1428]},
     {selectReadStageMask_lo[1427:1424]},
     {selectReadStageMask_lo[1423:1420]},
     {selectReadStageMask_lo[1419:1416]},
     {selectReadStageMask_lo[1415:1412]},
     {selectReadStageMask_lo[1411:1408]},
     {selectReadStageMask_lo[1407:1404]},
     {selectReadStageMask_lo[1403:1400]},
     {selectReadStageMask_lo[1399:1396]},
     {selectReadStageMask_lo[1395:1392]},
     {selectReadStageMask_lo[1391:1388]},
     {selectReadStageMask_lo[1387:1384]},
     {selectReadStageMask_lo[1383:1380]},
     {selectReadStageMask_lo[1379:1376]},
     {selectReadStageMask_lo[1375:1372]},
     {selectReadStageMask_lo[1371:1368]},
     {selectReadStageMask_lo[1367:1364]},
     {selectReadStageMask_lo[1363:1360]},
     {selectReadStageMask_lo[1359:1356]},
     {selectReadStageMask_lo[1355:1352]},
     {selectReadStageMask_lo[1351:1348]},
     {selectReadStageMask_lo[1347:1344]},
     {selectReadStageMask_lo[1343:1340]},
     {selectReadStageMask_lo[1339:1336]},
     {selectReadStageMask_lo[1335:1332]},
     {selectReadStageMask_lo[1331:1328]},
     {selectReadStageMask_lo[1327:1324]},
     {selectReadStageMask_lo[1323:1320]},
     {selectReadStageMask_lo[1319:1316]},
     {selectReadStageMask_lo[1315:1312]},
     {selectReadStageMask_lo[1311:1308]},
     {selectReadStageMask_lo[1307:1304]},
     {selectReadStageMask_lo[1303:1300]},
     {selectReadStageMask_lo[1299:1296]},
     {selectReadStageMask_lo[1295:1292]},
     {selectReadStageMask_lo[1291:1288]},
     {selectReadStageMask_lo[1287:1284]},
     {selectReadStageMask_lo[1283:1280]},
     {selectReadStageMask_lo[1279:1276]},
     {selectReadStageMask_lo[1275:1272]},
     {selectReadStageMask_lo[1271:1268]},
     {selectReadStageMask_lo[1267:1264]},
     {selectReadStageMask_lo[1263:1260]},
     {selectReadStageMask_lo[1259:1256]},
     {selectReadStageMask_lo[1255:1252]},
     {selectReadStageMask_lo[1251:1248]},
     {selectReadStageMask_lo[1247:1244]},
     {selectReadStageMask_lo[1243:1240]},
     {selectReadStageMask_lo[1239:1236]},
     {selectReadStageMask_lo[1235:1232]},
     {selectReadStageMask_lo[1231:1228]},
     {selectReadStageMask_lo[1227:1224]},
     {selectReadStageMask_lo[1223:1220]},
     {selectReadStageMask_lo[1219:1216]},
     {selectReadStageMask_lo[1215:1212]},
     {selectReadStageMask_lo[1211:1208]},
     {selectReadStageMask_lo[1207:1204]},
     {selectReadStageMask_lo[1203:1200]},
     {selectReadStageMask_lo[1199:1196]},
     {selectReadStageMask_lo[1195:1192]},
     {selectReadStageMask_lo[1191:1188]},
     {selectReadStageMask_lo[1187:1184]},
     {selectReadStageMask_lo[1183:1180]},
     {selectReadStageMask_lo[1179:1176]},
     {selectReadStageMask_lo[1175:1172]},
     {selectReadStageMask_lo[1171:1168]},
     {selectReadStageMask_lo[1167:1164]},
     {selectReadStageMask_lo[1163:1160]},
     {selectReadStageMask_lo[1159:1156]},
     {selectReadStageMask_lo[1155:1152]},
     {selectReadStageMask_lo[1151:1148]},
     {selectReadStageMask_lo[1147:1144]},
     {selectReadStageMask_lo[1143:1140]},
     {selectReadStageMask_lo[1139:1136]},
     {selectReadStageMask_lo[1135:1132]},
     {selectReadStageMask_lo[1131:1128]},
     {selectReadStageMask_lo[1127:1124]},
     {selectReadStageMask_lo[1123:1120]},
     {selectReadStageMask_lo[1119:1116]},
     {selectReadStageMask_lo[1115:1112]},
     {selectReadStageMask_lo[1111:1108]},
     {selectReadStageMask_lo[1107:1104]},
     {selectReadStageMask_lo[1103:1100]},
     {selectReadStageMask_lo[1099:1096]},
     {selectReadStageMask_lo[1095:1092]},
     {selectReadStageMask_lo[1091:1088]},
     {selectReadStageMask_lo[1087:1084]},
     {selectReadStageMask_lo[1083:1080]},
     {selectReadStageMask_lo[1079:1076]},
     {selectReadStageMask_lo[1075:1072]},
     {selectReadStageMask_lo[1071:1068]},
     {selectReadStageMask_lo[1067:1064]},
     {selectReadStageMask_lo[1063:1060]},
     {selectReadStageMask_lo[1059:1056]},
     {selectReadStageMask_lo[1055:1052]},
     {selectReadStageMask_lo[1051:1048]},
     {selectReadStageMask_lo[1047:1044]},
     {selectReadStageMask_lo[1043:1040]},
     {selectReadStageMask_lo[1039:1036]},
     {selectReadStageMask_lo[1035:1032]},
     {selectReadStageMask_lo[1031:1028]},
     {selectReadStageMask_lo[1027:1024]},
     {selectReadStageMask_lo[1023:1020]},
     {selectReadStageMask_lo[1019:1016]},
     {selectReadStageMask_lo[1015:1012]},
     {selectReadStageMask_lo[1011:1008]},
     {selectReadStageMask_lo[1007:1004]},
     {selectReadStageMask_lo[1003:1000]},
     {selectReadStageMask_lo[999:996]},
     {selectReadStageMask_lo[995:992]},
     {selectReadStageMask_lo[991:988]},
     {selectReadStageMask_lo[987:984]},
     {selectReadStageMask_lo[983:980]},
     {selectReadStageMask_lo[979:976]},
     {selectReadStageMask_lo[975:972]},
     {selectReadStageMask_lo[971:968]},
     {selectReadStageMask_lo[967:964]},
     {selectReadStageMask_lo[963:960]},
     {selectReadStageMask_lo[959:956]},
     {selectReadStageMask_lo[955:952]},
     {selectReadStageMask_lo[951:948]},
     {selectReadStageMask_lo[947:944]},
     {selectReadStageMask_lo[943:940]},
     {selectReadStageMask_lo[939:936]},
     {selectReadStageMask_lo[935:932]},
     {selectReadStageMask_lo[931:928]},
     {selectReadStageMask_lo[927:924]},
     {selectReadStageMask_lo[923:920]},
     {selectReadStageMask_lo[919:916]},
     {selectReadStageMask_lo[915:912]},
     {selectReadStageMask_lo[911:908]},
     {selectReadStageMask_lo[907:904]},
     {selectReadStageMask_lo[903:900]},
     {selectReadStageMask_lo[899:896]},
     {selectReadStageMask_lo[895:892]},
     {selectReadStageMask_lo[891:888]},
     {selectReadStageMask_lo[887:884]},
     {selectReadStageMask_lo[883:880]},
     {selectReadStageMask_lo[879:876]},
     {selectReadStageMask_lo[875:872]},
     {selectReadStageMask_lo[871:868]},
     {selectReadStageMask_lo[867:864]},
     {selectReadStageMask_lo[863:860]},
     {selectReadStageMask_lo[859:856]},
     {selectReadStageMask_lo[855:852]},
     {selectReadStageMask_lo[851:848]},
     {selectReadStageMask_lo[847:844]},
     {selectReadStageMask_lo[843:840]},
     {selectReadStageMask_lo[839:836]},
     {selectReadStageMask_lo[835:832]},
     {selectReadStageMask_lo[831:828]},
     {selectReadStageMask_lo[827:824]},
     {selectReadStageMask_lo[823:820]},
     {selectReadStageMask_lo[819:816]},
     {selectReadStageMask_lo[815:812]},
     {selectReadStageMask_lo[811:808]},
     {selectReadStageMask_lo[807:804]},
     {selectReadStageMask_lo[803:800]},
     {selectReadStageMask_lo[799:796]},
     {selectReadStageMask_lo[795:792]},
     {selectReadStageMask_lo[791:788]},
     {selectReadStageMask_lo[787:784]},
     {selectReadStageMask_lo[783:780]},
     {selectReadStageMask_lo[779:776]},
     {selectReadStageMask_lo[775:772]},
     {selectReadStageMask_lo[771:768]},
     {selectReadStageMask_lo[767:764]},
     {selectReadStageMask_lo[763:760]},
     {selectReadStageMask_lo[759:756]},
     {selectReadStageMask_lo[755:752]},
     {selectReadStageMask_lo[751:748]},
     {selectReadStageMask_lo[747:744]},
     {selectReadStageMask_lo[743:740]},
     {selectReadStageMask_lo[739:736]},
     {selectReadStageMask_lo[735:732]},
     {selectReadStageMask_lo[731:728]},
     {selectReadStageMask_lo[727:724]},
     {selectReadStageMask_lo[723:720]},
     {selectReadStageMask_lo[719:716]},
     {selectReadStageMask_lo[715:712]},
     {selectReadStageMask_lo[711:708]},
     {selectReadStageMask_lo[707:704]},
     {selectReadStageMask_lo[703:700]},
     {selectReadStageMask_lo[699:696]},
     {selectReadStageMask_lo[695:692]},
     {selectReadStageMask_lo[691:688]},
     {selectReadStageMask_lo[687:684]},
     {selectReadStageMask_lo[683:680]},
     {selectReadStageMask_lo[679:676]},
     {selectReadStageMask_lo[675:672]},
     {selectReadStageMask_lo[671:668]},
     {selectReadStageMask_lo[667:664]},
     {selectReadStageMask_lo[663:660]},
     {selectReadStageMask_lo[659:656]},
     {selectReadStageMask_lo[655:652]},
     {selectReadStageMask_lo[651:648]},
     {selectReadStageMask_lo[647:644]},
     {selectReadStageMask_lo[643:640]},
     {selectReadStageMask_lo[639:636]},
     {selectReadStageMask_lo[635:632]},
     {selectReadStageMask_lo[631:628]},
     {selectReadStageMask_lo[627:624]},
     {selectReadStageMask_lo[623:620]},
     {selectReadStageMask_lo[619:616]},
     {selectReadStageMask_lo[615:612]},
     {selectReadStageMask_lo[611:608]},
     {selectReadStageMask_lo[607:604]},
     {selectReadStageMask_lo[603:600]},
     {selectReadStageMask_lo[599:596]},
     {selectReadStageMask_lo[595:592]},
     {selectReadStageMask_lo[591:588]},
     {selectReadStageMask_lo[587:584]},
     {selectReadStageMask_lo[583:580]},
     {selectReadStageMask_lo[579:576]},
     {selectReadStageMask_lo[575:572]},
     {selectReadStageMask_lo[571:568]},
     {selectReadStageMask_lo[567:564]},
     {selectReadStageMask_lo[563:560]},
     {selectReadStageMask_lo[559:556]},
     {selectReadStageMask_lo[555:552]},
     {selectReadStageMask_lo[551:548]},
     {selectReadStageMask_lo[547:544]},
     {selectReadStageMask_lo[543:540]},
     {selectReadStageMask_lo[539:536]},
     {selectReadStageMask_lo[535:532]},
     {selectReadStageMask_lo[531:528]},
     {selectReadStageMask_lo[527:524]},
     {selectReadStageMask_lo[523:520]},
     {selectReadStageMask_lo[519:516]},
     {selectReadStageMask_lo[515:512]},
     {selectReadStageMask_lo[511:508]},
     {selectReadStageMask_lo[507:504]},
     {selectReadStageMask_lo[503:500]},
     {selectReadStageMask_lo[499:496]},
     {selectReadStageMask_lo[495:492]},
     {selectReadStageMask_lo[491:488]},
     {selectReadStageMask_lo[487:484]},
     {selectReadStageMask_lo[483:480]},
     {selectReadStageMask_lo[479:476]},
     {selectReadStageMask_lo[475:472]},
     {selectReadStageMask_lo[471:468]},
     {selectReadStageMask_lo[467:464]},
     {selectReadStageMask_lo[463:460]},
     {selectReadStageMask_lo[459:456]},
     {selectReadStageMask_lo[455:452]},
     {selectReadStageMask_lo[451:448]},
     {selectReadStageMask_lo[447:444]},
     {selectReadStageMask_lo[443:440]},
     {selectReadStageMask_lo[439:436]},
     {selectReadStageMask_lo[435:432]},
     {selectReadStageMask_lo[431:428]},
     {selectReadStageMask_lo[427:424]},
     {selectReadStageMask_lo[423:420]},
     {selectReadStageMask_lo[419:416]},
     {selectReadStageMask_lo[415:412]},
     {selectReadStageMask_lo[411:408]},
     {selectReadStageMask_lo[407:404]},
     {selectReadStageMask_lo[403:400]},
     {selectReadStageMask_lo[399:396]},
     {selectReadStageMask_lo[395:392]},
     {selectReadStageMask_lo[391:388]},
     {selectReadStageMask_lo[387:384]},
     {selectReadStageMask_lo[383:380]},
     {selectReadStageMask_lo[379:376]},
     {selectReadStageMask_lo[375:372]},
     {selectReadStageMask_lo[371:368]},
     {selectReadStageMask_lo[367:364]},
     {selectReadStageMask_lo[363:360]},
     {selectReadStageMask_lo[359:356]},
     {selectReadStageMask_lo[355:352]},
     {selectReadStageMask_lo[351:348]},
     {selectReadStageMask_lo[347:344]},
     {selectReadStageMask_lo[343:340]},
     {selectReadStageMask_lo[339:336]},
     {selectReadStageMask_lo[335:332]},
     {selectReadStageMask_lo[331:328]},
     {selectReadStageMask_lo[327:324]},
     {selectReadStageMask_lo[323:320]},
     {selectReadStageMask_lo[319:316]},
     {selectReadStageMask_lo[315:312]},
     {selectReadStageMask_lo[311:308]},
     {selectReadStageMask_lo[307:304]},
     {selectReadStageMask_lo[303:300]},
     {selectReadStageMask_lo[299:296]},
     {selectReadStageMask_lo[295:292]},
     {selectReadStageMask_lo[291:288]},
     {selectReadStageMask_lo[287:284]},
     {selectReadStageMask_lo[283:280]},
     {selectReadStageMask_lo[279:276]},
     {selectReadStageMask_lo[275:272]},
     {selectReadStageMask_lo[271:268]},
     {selectReadStageMask_lo[267:264]},
     {selectReadStageMask_lo[263:260]},
     {selectReadStageMask_lo[259:256]},
     {selectReadStageMask_lo[255:252]},
     {selectReadStageMask_lo[251:248]},
     {selectReadStageMask_lo[247:244]},
     {selectReadStageMask_lo[243:240]},
     {selectReadStageMask_lo[239:236]},
     {selectReadStageMask_lo[235:232]},
     {selectReadStageMask_lo[231:228]},
     {selectReadStageMask_lo[227:224]},
     {selectReadStageMask_lo[223:220]},
     {selectReadStageMask_lo[219:216]},
     {selectReadStageMask_lo[215:212]},
     {selectReadStageMask_lo[211:208]},
     {selectReadStageMask_lo[207:204]},
     {selectReadStageMask_lo[203:200]},
     {selectReadStageMask_lo[199:196]},
     {selectReadStageMask_lo[195:192]},
     {selectReadStageMask_lo[191:188]},
     {selectReadStageMask_lo[187:184]},
     {selectReadStageMask_lo[183:180]},
     {selectReadStageMask_lo[179:176]},
     {selectReadStageMask_lo[175:172]},
     {selectReadStageMask_lo[171:168]},
     {selectReadStageMask_lo[167:164]},
     {selectReadStageMask_lo[163:160]},
     {selectReadStageMask_lo[159:156]},
     {selectReadStageMask_lo[155:152]},
     {selectReadStageMask_lo[151:148]},
     {selectReadStageMask_lo[147:144]},
     {selectReadStageMask_lo[143:140]},
     {selectReadStageMask_lo[139:136]},
     {selectReadStageMask_lo[135:132]},
     {selectReadStageMask_lo[131:128]},
     {selectReadStageMask_lo[127:124]},
     {selectReadStageMask_lo[123:120]},
     {selectReadStageMask_lo[119:116]},
     {selectReadStageMask_lo[115:112]},
     {selectReadStageMask_lo[111:108]},
     {selectReadStageMask_lo[107:104]},
     {selectReadStageMask_lo[103:100]},
     {selectReadStageMask_lo[99:96]},
     {selectReadStageMask_lo[95:92]},
     {selectReadStageMask_lo[91:88]},
     {selectReadStageMask_lo[87:84]},
     {selectReadStageMask_lo[83:80]},
     {selectReadStageMask_lo[79:76]},
     {selectReadStageMask_lo[75:72]},
     {selectReadStageMask_lo[71:68]},
     {selectReadStageMask_lo[67:64]},
     {selectReadStageMask_lo[63:60]},
     {selectReadStageMask_lo[59:56]},
     {selectReadStageMask_lo[55:52]},
     {selectReadStageMask_lo[51:48]},
     {selectReadStageMask_lo[47:44]},
     {selectReadStageMask_lo[43:40]},
     {selectReadStageMask_lo[39:36]},
     {selectReadStageMask_lo[35:32]},
     {selectReadStageMask_lo[31:28]},
     {selectReadStageMask_lo[27:24]},
     {selectReadStageMask_lo[23:20]},
     {selectReadStageMask_lo[19:16]},
     {selectReadStageMask_lo[15:12]},
     {selectReadStageMask_lo[11:8]},
     {selectReadStageMask_lo[7:4]},
     {selectReadStageMask_lo[3:0]}};
  wire [3:0]         readMaskCorrection = (instReg_maskType ? _GEN_142[executeGroup[10:0]] : 4'hF) & vlBoundaryCorrection;
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_lo_lo_lo = {maskSplit_maskSelect_lo_lo_lo_lo_lo_lo_hi, maskSplit_maskSelect_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_lo_lo_hi = {maskSplit_maskSelect_lo_lo_lo_lo_lo_hi_hi, maskSplit_maskSelect_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]       maskSplit_maskSelect_lo_lo_lo_lo_lo = {maskSplit_maskSelect_lo_lo_lo_lo_lo_hi, maskSplit_maskSelect_lo_lo_lo_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_lo_hi_lo = {maskSplit_maskSelect_lo_lo_lo_lo_hi_lo_hi, maskSplit_maskSelect_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_lo_hi_hi = {maskSplit_maskSelect_lo_lo_lo_lo_hi_hi_hi, maskSplit_maskSelect_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]       maskSplit_maskSelect_lo_lo_lo_lo_hi = {maskSplit_maskSelect_lo_lo_lo_lo_hi_hi, maskSplit_maskSelect_lo_lo_lo_lo_hi_lo};
  wire [511:0]       maskSplit_maskSelect_lo_lo_lo_lo = {maskSplit_maskSelect_lo_lo_lo_lo_hi, maskSplit_maskSelect_lo_lo_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_hi_lo_lo = {maskSplit_maskSelect_lo_lo_lo_hi_lo_lo_hi, maskSplit_maskSelect_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_hi_lo_hi = {maskSplit_maskSelect_lo_lo_lo_hi_lo_hi_hi, maskSplit_maskSelect_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]       maskSplit_maskSelect_lo_lo_lo_hi_lo = {maskSplit_maskSelect_lo_lo_lo_hi_lo_hi, maskSplit_maskSelect_lo_lo_lo_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_hi_hi_lo = {maskSplit_maskSelect_lo_lo_lo_hi_hi_lo_hi, maskSplit_maskSelect_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_hi_hi_hi = {maskSplit_maskSelect_lo_lo_lo_hi_hi_hi_hi, maskSplit_maskSelect_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]       maskSplit_maskSelect_lo_lo_lo_hi_hi = {maskSplit_maskSelect_lo_lo_lo_hi_hi_hi, maskSplit_maskSelect_lo_lo_lo_hi_hi_lo};
  wire [511:0]       maskSplit_maskSelect_lo_lo_lo_hi = {maskSplit_maskSelect_lo_lo_lo_hi_hi, maskSplit_maskSelect_lo_lo_lo_hi_lo};
  wire [1023:0]      maskSplit_maskSelect_lo_lo_lo = {maskSplit_maskSelect_lo_lo_lo_hi, maskSplit_maskSelect_lo_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_lo_lo_lo = {maskSplit_maskSelect_lo_lo_hi_lo_lo_lo_hi, maskSplit_maskSelect_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_lo_lo_hi = {maskSplit_maskSelect_lo_lo_hi_lo_lo_hi_hi, maskSplit_maskSelect_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]       maskSplit_maskSelect_lo_lo_hi_lo_lo = {maskSplit_maskSelect_lo_lo_hi_lo_lo_hi, maskSplit_maskSelect_lo_lo_hi_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_lo_hi_lo = {maskSplit_maskSelect_lo_lo_hi_lo_hi_lo_hi, maskSplit_maskSelect_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_lo_hi_hi = {maskSplit_maskSelect_lo_lo_hi_lo_hi_hi_hi, maskSplit_maskSelect_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]       maskSplit_maskSelect_lo_lo_hi_lo_hi = {maskSplit_maskSelect_lo_lo_hi_lo_hi_hi, maskSplit_maskSelect_lo_lo_hi_lo_hi_lo};
  wire [511:0]       maskSplit_maskSelect_lo_lo_hi_lo = {maskSplit_maskSelect_lo_lo_hi_lo_hi, maskSplit_maskSelect_lo_lo_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_hi_lo_lo = {maskSplit_maskSelect_lo_lo_hi_hi_lo_lo_hi, maskSplit_maskSelect_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_hi_lo_hi = {maskSplit_maskSelect_lo_lo_hi_hi_lo_hi_hi, maskSplit_maskSelect_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]       maskSplit_maskSelect_lo_lo_hi_hi_lo = {maskSplit_maskSelect_lo_lo_hi_hi_lo_hi, maskSplit_maskSelect_lo_lo_hi_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_hi_hi_lo = {maskSplit_maskSelect_lo_lo_hi_hi_hi_lo_hi, maskSplit_maskSelect_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_hi_hi_hi = {maskSplit_maskSelect_lo_lo_hi_hi_hi_hi_hi, maskSplit_maskSelect_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]       maskSplit_maskSelect_lo_lo_hi_hi_hi = {maskSplit_maskSelect_lo_lo_hi_hi_hi_hi, maskSplit_maskSelect_lo_lo_hi_hi_hi_lo};
  wire [511:0]       maskSplit_maskSelect_lo_lo_hi_hi = {maskSplit_maskSelect_lo_lo_hi_hi_hi, maskSplit_maskSelect_lo_lo_hi_hi_lo};
  wire [1023:0]      maskSplit_maskSelect_lo_lo_hi = {maskSplit_maskSelect_lo_lo_hi_hi, maskSplit_maskSelect_lo_lo_hi_lo};
  wire [2047:0]      maskSplit_maskSelect_lo_lo = {maskSplit_maskSelect_lo_lo_hi, maskSplit_maskSelect_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_lo_lo_lo = {maskSplit_maskSelect_lo_hi_lo_lo_lo_lo_hi, maskSplit_maskSelect_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_lo_lo_hi = {maskSplit_maskSelect_lo_hi_lo_lo_lo_hi_hi, maskSplit_maskSelect_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]       maskSplit_maskSelect_lo_hi_lo_lo_lo = {maskSplit_maskSelect_lo_hi_lo_lo_lo_hi, maskSplit_maskSelect_lo_hi_lo_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_lo_hi_lo = {maskSplit_maskSelect_lo_hi_lo_lo_hi_lo_hi, maskSplit_maskSelect_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_lo_hi_hi = {maskSplit_maskSelect_lo_hi_lo_lo_hi_hi_hi, maskSplit_maskSelect_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]       maskSplit_maskSelect_lo_hi_lo_lo_hi = {maskSplit_maskSelect_lo_hi_lo_lo_hi_hi, maskSplit_maskSelect_lo_hi_lo_lo_hi_lo};
  wire [511:0]       maskSplit_maskSelect_lo_hi_lo_lo = {maskSplit_maskSelect_lo_hi_lo_lo_hi, maskSplit_maskSelect_lo_hi_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_hi_lo_lo = {maskSplit_maskSelect_lo_hi_lo_hi_lo_lo_hi, maskSplit_maskSelect_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_hi_lo_hi = {maskSplit_maskSelect_lo_hi_lo_hi_lo_hi_hi, maskSplit_maskSelect_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]       maskSplit_maskSelect_lo_hi_lo_hi_lo = {maskSplit_maskSelect_lo_hi_lo_hi_lo_hi, maskSplit_maskSelect_lo_hi_lo_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_hi_hi_lo = {maskSplit_maskSelect_lo_hi_lo_hi_hi_lo_hi, maskSplit_maskSelect_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_hi_hi_hi = {maskSplit_maskSelect_lo_hi_lo_hi_hi_hi_hi, maskSplit_maskSelect_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]       maskSplit_maskSelect_lo_hi_lo_hi_hi = {maskSplit_maskSelect_lo_hi_lo_hi_hi_hi, maskSplit_maskSelect_lo_hi_lo_hi_hi_lo};
  wire [511:0]       maskSplit_maskSelect_lo_hi_lo_hi = {maskSplit_maskSelect_lo_hi_lo_hi_hi, maskSplit_maskSelect_lo_hi_lo_hi_lo};
  wire [1023:0]      maskSplit_maskSelect_lo_hi_lo = {maskSplit_maskSelect_lo_hi_lo_hi, maskSplit_maskSelect_lo_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_lo_lo_lo = {maskSplit_maskSelect_lo_hi_hi_lo_lo_lo_hi, maskSplit_maskSelect_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_lo_lo_hi = {maskSplit_maskSelect_lo_hi_hi_lo_lo_hi_hi, maskSplit_maskSelect_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]       maskSplit_maskSelect_lo_hi_hi_lo_lo = {maskSplit_maskSelect_lo_hi_hi_lo_lo_hi, maskSplit_maskSelect_lo_hi_hi_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_lo_hi_lo = {maskSplit_maskSelect_lo_hi_hi_lo_hi_lo_hi, maskSplit_maskSelect_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_lo_hi_hi = {maskSplit_maskSelect_lo_hi_hi_lo_hi_hi_hi, maskSplit_maskSelect_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]       maskSplit_maskSelect_lo_hi_hi_lo_hi = {maskSplit_maskSelect_lo_hi_hi_lo_hi_hi, maskSplit_maskSelect_lo_hi_hi_lo_hi_lo};
  wire [511:0]       maskSplit_maskSelect_lo_hi_hi_lo = {maskSplit_maskSelect_lo_hi_hi_lo_hi, maskSplit_maskSelect_lo_hi_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_hi_lo_lo = {maskSplit_maskSelect_lo_hi_hi_hi_lo_lo_hi, maskSplit_maskSelect_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_hi_lo_hi = {maskSplit_maskSelect_lo_hi_hi_hi_lo_hi_hi, maskSplit_maskSelect_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]       maskSplit_maskSelect_lo_hi_hi_hi_lo = {maskSplit_maskSelect_lo_hi_hi_hi_lo_hi, maskSplit_maskSelect_lo_hi_hi_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_hi_hi_lo = {maskSplit_maskSelect_lo_hi_hi_hi_hi_lo_hi, maskSplit_maskSelect_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_hi_hi_hi = {maskSplit_maskSelect_lo_hi_hi_hi_hi_hi_hi, maskSplit_maskSelect_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]       maskSplit_maskSelect_lo_hi_hi_hi_hi = {maskSplit_maskSelect_lo_hi_hi_hi_hi_hi, maskSplit_maskSelect_lo_hi_hi_hi_hi_lo};
  wire [511:0]       maskSplit_maskSelect_lo_hi_hi_hi = {maskSplit_maskSelect_lo_hi_hi_hi_hi, maskSplit_maskSelect_lo_hi_hi_hi_lo};
  wire [1023:0]      maskSplit_maskSelect_lo_hi_hi = {maskSplit_maskSelect_lo_hi_hi_hi, maskSplit_maskSelect_lo_hi_hi_lo};
  wire [2047:0]      maskSplit_maskSelect_lo_hi = {maskSplit_maskSelect_lo_hi_hi, maskSplit_maskSelect_lo_hi_lo};
  wire [4095:0]      maskSplit_maskSelect_lo = {maskSplit_maskSelect_lo_hi, maskSplit_maskSelect_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_lo_lo_lo = {maskSplit_maskSelect_hi_lo_lo_lo_lo_lo_hi, maskSplit_maskSelect_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_lo_lo_hi = {maskSplit_maskSelect_hi_lo_lo_lo_lo_hi_hi, maskSplit_maskSelect_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]       maskSplit_maskSelect_hi_lo_lo_lo_lo = {maskSplit_maskSelect_hi_lo_lo_lo_lo_hi, maskSplit_maskSelect_hi_lo_lo_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_lo_hi_lo = {maskSplit_maskSelect_hi_lo_lo_lo_hi_lo_hi, maskSplit_maskSelect_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_lo_hi_hi = {maskSplit_maskSelect_hi_lo_lo_lo_hi_hi_hi, maskSplit_maskSelect_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]       maskSplit_maskSelect_hi_lo_lo_lo_hi = {maskSplit_maskSelect_hi_lo_lo_lo_hi_hi, maskSplit_maskSelect_hi_lo_lo_lo_hi_lo};
  wire [511:0]       maskSplit_maskSelect_hi_lo_lo_lo = {maskSplit_maskSelect_hi_lo_lo_lo_hi, maskSplit_maskSelect_hi_lo_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_hi_lo_lo = {maskSplit_maskSelect_hi_lo_lo_hi_lo_lo_hi, maskSplit_maskSelect_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_hi_lo_hi = {maskSplit_maskSelect_hi_lo_lo_hi_lo_hi_hi, maskSplit_maskSelect_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]       maskSplit_maskSelect_hi_lo_lo_hi_lo = {maskSplit_maskSelect_hi_lo_lo_hi_lo_hi, maskSplit_maskSelect_hi_lo_lo_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_hi_hi_lo = {maskSplit_maskSelect_hi_lo_lo_hi_hi_lo_hi, maskSplit_maskSelect_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_hi_hi_hi = {maskSplit_maskSelect_hi_lo_lo_hi_hi_hi_hi, maskSplit_maskSelect_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]       maskSplit_maskSelect_hi_lo_lo_hi_hi = {maskSplit_maskSelect_hi_lo_lo_hi_hi_hi, maskSplit_maskSelect_hi_lo_lo_hi_hi_lo};
  wire [511:0]       maskSplit_maskSelect_hi_lo_lo_hi = {maskSplit_maskSelect_hi_lo_lo_hi_hi, maskSplit_maskSelect_hi_lo_lo_hi_lo};
  wire [1023:0]      maskSplit_maskSelect_hi_lo_lo = {maskSplit_maskSelect_hi_lo_lo_hi, maskSplit_maskSelect_hi_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_lo_lo_lo = {maskSplit_maskSelect_hi_lo_hi_lo_lo_lo_hi, maskSplit_maskSelect_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_lo_lo_hi = {maskSplit_maskSelect_hi_lo_hi_lo_lo_hi_hi, maskSplit_maskSelect_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]       maskSplit_maskSelect_hi_lo_hi_lo_lo = {maskSplit_maskSelect_hi_lo_hi_lo_lo_hi, maskSplit_maskSelect_hi_lo_hi_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_lo_hi_lo = {maskSplit_maskSelect_hi_lo_hi_lo_hi_lo_hi, maskSplit_maskSelect_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_lo_hi_hi = {maskSplit_maskSelect_hi_lo_hi_lo_hi_hi_hi, maskSplit_maskSelect_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]       maskSplit_maskSelect_hi_lo_hi_lo_hi = {maskSplit_maskSelect_hi_lo_hi_lo_hi_hi, maskSplit_maskSelect_hi_lo_hi_lo_hi_lo};
  wire [511:0]       maskSplit_maskSelect_hi_lo_hi_lo = {maskSplit_maskSelect_hi_lo_hi_lo_hi, maskSplit_maskSelect_hi_lo_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_hi_lo_lo = {maskSplit_maskSelect_hi_lo_hi_hi_lo_lo_hi, maskSplit_maskSelect_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_hi_lo_hi = {maskSplit_maskSelect_hi_lo_hi_hi_lo_hi_hi, maskSplit_maskSelect_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]       maskSplit_maskSelect_hi_lo_hi_hi_lo = {maskSplit_maskSelect_hi_lo_hi_hi_lo_hi, maskSplit_maskSelect_hi_lo_hi_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_hi_hi_lo = {maskSplit_maskSelect_hi_lo_hi_hi_hi_lo_hi, maskSplit_maskSelect_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_hi_hi_hi = {maskSplit_maskSelect_hi_lo_hi_hi_hi_hi_hi, maskSplit_maskSelect_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]       maskSplit_maskSelect_hi_lo_hi_hi_hi = {maskSplit_maskSelect_hi_lo_hi_hi_hi_hi, maskSplit_maskSelect_hi_lo_hi_hi_hi_lo};
  wire [511:0]       maskSplit_maskSelect_hi_lo_hi_hi = {maskSplit_maskSelect_hi_lo_hi_hi_hi, maskSplit_maskSelect_hi_lo_hi_hi_lo};
  wire [1023:0]      maskSplit_maskSelect_hi_lo_hi = {maskSplit_maskSelect_hi_lo_hi_hi, maskSplit_maskSelect_hi_lo_hi_lo};
  wire [2047:0]      maskSplit_maskSelect_hi_lo = {maskSplit_maskSelect_hi_lo_hi, maskSplit_maskSelect_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_lo_lo_lo = {maskSplit_maskSelect_hi_hi_lo_lo_lo_lo_hi, maskSplit_maskSelect_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_lo_lo_hi = {maskSplit_maskSelect_hi_hi_lo_lo_lo_hi_hi, maskSplit_maskSelect_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]       maskSplit_maskSelect_hi_hi_lo_lo_lo = {maskSplit_maskSelect_hi_hi_lo_lo_lo_hi, maskSplit_maskSelect_hi_hi_lo_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_lo_hi_lo = {maskSplit_maskSelect_hi_hi_lo_lo_hi_lo_hi, maskSplit_maskSelect_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_lo_hi_hi = {maskSplit_maskSelect_hi_hi_lo_lo_hi_hi_hi, maskSplit_maskSelect_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]       maskSplit_maskSelect_hi_hi_lo_lo_hi = {maskSplit_maskSelect_hi_hi_lo_lo_hi_hi, maskSplit_maskSelect_hi_hi_lo_lo_hi_lo};
  wire [511:0]       maskSplit_maskSelect_hi_hi_lo_lo = {maskSplit_maskSelect_hi_hi_lo_lo_hi, maskSplit_maskSelect_hi_hi_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_hi_lo_lo = {maskSplit_maskSelect_hi_hi_lo_hi_lo_lo_hi, maskSplit_maskSelect_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_hi_lo_hi = {maskSplit_maskSelect_hi_hi_lo_hi_lo_hi_hi, maskSplit_maskSelect_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]       maskSplit_maskSelect_hi_hi_lo_hi_lo = {maskSplit_maskSelect_hi_hi_lo_hi_lo_hi, maskSplit_maskSelect_hi_hi_lo_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_hi_hi_lo = {maskSplit_maskSelect_hi_hi_lo_hi_hi_lo_hi, maskSplit_maskSelect_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_hi_hi_hi = {maskSplit_maskSelect_hi_hi_lo_hi_hi_hi_hi, maskSplit_maskSelect_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]       maskSplit_maskSelect_hi_hi_lo_hi_hi = {maskSplit_maskSelect_hi_hi_lo_hi_hi_hi, maskSplit_maskSelect_hi_hi_lo_hi_hi_lo};
  wire [511:0]       maskSplit_maskSelect_hi_hi_lo_hi = {maskSplit_maskSelect_hi_hi_lo_hi_hi, maskSplit_maskSelect_hi_hi_lo_hi_lo};
  wire [1023:0]      maskSplit_maskSelect_hi_hi_lo = {maskSplit_maskSelect_hi_hi_lo_hi, maskSplit_maskSelect_hi_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_lo_lo_lo = {maskSplit_maskSelect_hi_hi_hi_lo_lo_lo_hi, maskSplit_maskSelect_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_lo_lo_hi = {maskSplit_maskSelect_hi_hi_hi_lo_lo_hi_hi, maskSplit_maskSelect_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]       maskSplit_maskSelect_hi_hi_hi_lo_lo = {maskSplit_maskSelect_hi_hi_hi_lo_lo_hi, maskSplit_maskSelect_hi_hi_hi_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_lo_hi_lo = {maskSplit_maskSelect_hi_hi_hi_lo_hi_lo_hi, maskSplit_maskSelect_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_lo_hi_hi = {maskSplit_maskSelect_hi_hi_hi_lo_hi_hi_hi, maskSplit_maskSelect_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]       maskSplit_maskSelect_hi_hi_hi_lo_hi = {maskSplit_maskSelect_hi_hi_hi_lo_hi_hi, maskSplit_maskSelect_hi_hi_hi_lo_hi_lo};
  wire [511:0]       maskSplit_maskSelect_hi_hi_hi_lo = {maskSplit_maskSelect_hi_hi_hi_lo_hi, maskSplit_maskSelect_hi_hi_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_hi_lo_lo = {maskSplit_maskSelect_hi_hi_hi_hi_lo_lo_hi, maskSplit_maskSelect_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_hi_lo_hi = {maskSplit_maskSelect_hi_hi_hi_hi_lo_hi_hi, maskSplit_maskSelect_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]       maskSplit_maskSelect_hi_hi_hi_hi_lo = {maskSplit_maskSelect_hi_hi_hi_hi_lo_hi, maskSplit_maskSelect_hi_hi_hi_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_hi_hi_lo = {maskSplit_maskSelect_hi_hi_hi_hi_hi_lo_hi, maskSplit_maskSelect_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_hi_hi_hi = {maskSplit_maskSelect_hi_hi_hi_hi_hi_hi_hi, maskSplit_maskSelect_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]       maskSplit_maskSelect_hi_hi_hi_hi_hi = {maskSplit_maskSelect_hi_hi_hi_hi_hi_hi, maskSplit_maskSelect_hi_hi_hi_hi_hi_lo};
  wire [511:0]       maskSplit_maskSelect_hi_hi_hi_hi = {maskSplit_maskSelect_hi_hi_hi_hi_hi, maskSplit_maskSelect_hi_hi_hi_hi_lo};
  wire [1023:0]      maskSplit_maskSelect_hi_hi_hi = {maskSplit_maskSelect_hi_hi_hi_hi, maskSplit_maskSelect_hi_hi_hi_lo};
  wire [2047:0]      maskSplit_maskSelect_hi_hi = {maskSplit_maskSelect_hi_hi_hi, maskSplit_maskSelect_hi_hi_lo};
  wire [4095:0]      maskSplit_maskSelect_hi = {maskSplit_maskSelect_hi_hi, maskSplit_maskSelect_hi_lo};
  wire [9:0]         executeGroupCounter;
  wire               maskSplit_vlMisAlign = |(instReg_vl[3:0]);
  wire [9:0]         maskSplit_lastexecuteGroup = instReg_vl[13:4] - {9'h0, ~maskSplit_vlMisAlign};
  wire               maskSplit_isVlBoundary = executeGroupCounter == maskSplit_lastexecuteGroup;
  wire               maskSplit_validExecuteGroup = executeGroupCounter <= maskSplit_lastexecuteGroup;
  wire [15:0]        _maskSplit_vlBoundaryCorrection_T_2 = 16'h1 << instReg_vl[3:0];
  wire [15:0]        _maskSplit_vlBoundaryCorrection_T_5 = _maskSplit_vlBoundaryCorrection_T_2 | {_maskSplit_vlBoundaryCorrection_T_2[14:0], 1'h0};
  wire [15:0]        _maskSplit_vlBoundaryCorrection_T_8 = _maskSplit_vlBoundaryCorrection_T_5 | {_maskSplit_vlBoundaryCorrection_T_5[13:0], 2'h0};
  wire [15:0]        _maskSplit_vlBoundaryCorrection_T_11 = _maskSplit_vlBoundaryCorrection_T_8 | {_maskSplit_vlBoundaryCorrection_T_8[11:0], 4'h0};
  wire [15:0]        maskSplit_vlBoundaryCorrection = ~({16{maskSplit_vlMisAlign & maskSplit_isVlBoundary}} & (_maskSplit_vlBoundaryCorrection_T_11 | {_maskSplit_vlBoundaryCorrection_T_11[7:0], 8'h0})) & {16{maskSplit_validExecuteGroup}};
  wire [511:0][15:0] _GEN_143 =
    {{maskSplit_maskSelect_hi[4095:4080]},
     {maskSplit_maskSelect_hi[4079:4064]},
     {maskSplit_maskSelect_hi[4063:4048]},
     {maskSplit_maskSelect_hi[4047:4032]},
     {maskSplit_maskSelect_hi[4031:4016]},
     {maskSplit_maskSelect_hi[4015:4000]},
     {maskSplit_maskSelect_hi[3999:3984]},
     {maskSplit_maskSelect_hi[3983:3968]},
     {maskSplit_maskSelect_hi[3967:3952]},
     {maskSplit_maskSelect_hi[3951:3936]},
     {maskSplit_maskSelect_hi[3935:3920]},
     {maskSplit_maskSelect_hi[3919:3904]},
     {maskSplit_maskSelect_hi[3903:3888]},
     {maskSplit_maskSelect_hi[3887:3872]},
     {maskSplit_maskSelect_hi[3871:3856]},
     {maskSplit_maskSelect_hi[3855:3840]},
     {maskSplit_maskSelect_hi[3839:3824]},
     {maskSplit_maskSelect_hi[3823:3808]},
     {maskSplit_maskSelect_hi[3807:3792]},
     {maskSplit_maskSelect_hi[3791:3776]},
     {maskSplit_maskSelect_hi[3775:3760]},
     {maskSplit_maskSelect_hi[3759:3744]},
     {maskSplit_maskSelect_hi[3743:3728]},
     {maskSplit_maskSelect_hi[3727:3712]},
     {maskSplit_maskSelect_hi[3711:3696]},
     {maskSplit_maskSelect_hi[3695:3680]},
     {maskSplit_maskSelect_hi[3679:3664]},
     {maskSplit_maskSelect_hi[3663:3648]},
     {maskSplit_maskSelect_hi[3647:3632]},
     {maskSplit_maskSelect_hi[3631:3616]},
     {maskSplit_maskSelect_hi[3615:3600]},
     {maskSplit_maskSelect_hi[3599:3584]},
     {maskSplit_maskSelect_hi[3583:3568]},
     {maskSplit_maskSelect_hi[3567:3552]},
     {maskSplit_maskSelect_hi[3551:3536]},
     {maskSplit_maskSelect_hi[3535:3520]},
     {maskSplit_maskSelect_hi[3519:3504]},
     {maskSplit_maskSelect_hi[3503:3488]},
     {maskSplit_maskSelect_hi[3487:3472]},
     {maskSplit_maskSelect_hi[3471:3456]},
     {maskSplit_maskSelect_hi[3455:3440]},
     {maskSplit_maskSelect_hi[3439:3424]},
     {maskSplit_maskSelect_hi[3423:3408]},
     {maskSplit_maskSelect_hi[3407:3392]},
     {maskSplit_maskSelect_hi[3391:3376]},
     {maskSplit_maskSelect_hi[3375:3360]},
     {maskSplit_maskSelect_hi[3359:3344]},
     {maskSplit_maskSelect_hi[3343:3328]},
     {maskSplit_maskSelect_hi[3327:3312]},
     {maskSplit_maskSelect_hi[3311:3296]},
     {maskSplit_maskSelect_hi[3295:3280]},
     {maskSplit_maskSelect_hi[3279:3264]},
     {maskSplit_maskSelect_hi[3263:3248]},
     {maskSplit_maskSelect_hi[3247:3232]},
     {maskSplit_maskSelect_hi[3231:3216]},
     {maskSplit_maskSelect_hi[3215:3200]},
     {maskSplit_maskSelect_hi[3199:3184]},
     {maskSplit_maskSelect_hi[3183:3168]},
     {maskSplit_maskSelect_hi[3167:3152]},
     {maskSplit_maskSelect_hi[3151:3136]},
     {maskSplit_maskSelect_hi[3135:3120]},
     {maskSplit_maskSelect_hi[3119:3104]},
     {maskSplit_maskSelect_hi[3103:3088]},
     {maskSplit_maskSelect_hi[3087:3072]},
     {maskSplit_maskSelect_hi[3071:3056]},
     {maskSplit_maskSelect_hi[3055:3040]},
     {maskSplit_maskSelect_hi[3039:3024]},
     {maskSplit_maskSelect_hi[3023:3008]},
     {maskSplit_maskSelect_hi[3007:2992]},
     {maskSplit_maskSelect_hi[2991:2976]},
     {maskSplit_maskSelect_hi[2975:2960]},
     {maskSplit_maskSelect_hi[2959:2944]},
     {maskSplit_maskSelect_hi[2943:2928]},
     {maskSplit_maskSelect_hi[2927:2912]},
     {maskSplit_maskSelect_hi[2911:2896]},
     {maskSplit_maskSelect_hi[2895:2880]},
     {maskSplit_maskSelect_hi[2879:2864]},
     {maskSplit_maskSelect_hi[2863:2848]},
     {maskSplit_maskSelect_hi[2847:2832]},
     {maskSplit_maskSelect_hi[2831:2816]},
     {maskSplit_maskSelect_hi[2815:2800]},
     {maskSplit_maskSelect_hi[2799:2784]},
     {maskSplit_maskSelect_hi[2783:2768]},
     {maskSplit_maskSelect_hi[2767:2752]},
     {maskSplit_maskSelect_hi[2751:2736]},
     {maskSplit_maskSelect_hi[2735:2720]},
     {maskSplit_maskSelect_hi[2719:2704]},
     {maskSplit_maskSelect_hi[2703:2688]},
     {maskSplit_maskSelect_hi[2687:2672]},
     {maskSplit_maskSelect_hi[2671:2656]},
     {maskSplit_maskSelect_hi[2655:2640]},
     {maskSplit_maskSelect_hi[2639:2624]},
     {maskSplit_maskSelect_hi[2623:2608]},
     {maskSplit_maskSelect_hi[2607:2592]},
     {maskSplit_maskSelect_hi[2591:2576]},
     {maskSplit_maskSelect_hi[2575:2560]},
     {maskSplit_maskSelect_hi[2559:2544]},
     {maskSplit_maskSelect_hi[2543:2528]},
     {maskSplit_maskSelect_hi[2527:2512]},
     {maskSplit_maskSelect_hi[2511:2496]},
     {maskSplit_maskSelect_hi[2495:2480]},
     {maskSplit_maskSelect_hi[2479:2464]},
     {maskSplit_maskSelect_hi[2463:2448]},
     {maskSplit_maskSelect_hi[2447:2432]},
     {maskSplit_maskSelect_hi[2431:2416]},
     {maskSplit_maskSelect_hi[2415:2400]},
     {maskSplit_maskSelect_hi[2399:2384]},
     {maskSplit_maskSelect_hi[2383:2368]},
     {maskSplit_maskSelect_hi[2367:2352]},
     {maskSplit_maskSelect_hi[2351:2336]},
     {maskSplit_maskSelect_hi[2335:2320]},
     {maskSplit_maskSelect_hi[2319:2304]},
     {maskSplit_maskSelect_hi[2303:2288]},
     {maskSplit_maskSelect_hi[2287:2272]},
     {maskSplit_maskSelect_hi[2271:2256]},
     {maskSplit_maskSelect_hi[2255:2240]},
     {maskSplit_maskSelect_hi[2239:2224]},
     {maskSplit_maskSelect_hi[2223:2208]},
     {maskSplit_maskSelect_hi[2207:2192]},
     {maskSplit_maskSelect_hi[2191:2176]},
     {maskSplit_maskSelect_hi[2175:2160]},
     {maskSplit_maskSelect_hi[2159:2144]},
     {maskSplit_maskSelect_hi[2143:2128]},
     {maskSplit_maskSelect_hi[2127:2112]},
     {maskSplit_maskSelect_hi[2111:2096]},
     {maskSplit_maskSelect_hi[2095:2080]},
     {maskSplit_maskSelect_hi[2079:2064]},
     {maskSplit_maskSelect_hi[2063:2048]},
     {maskSplit_maskSelect_hi[2047:2032]},
     {maskSplit_maskSelect_hi[2031:2016]},
     {maskSplit_maskSelect_hi[2015:2000]},
     {maskSplit_maskSelect_hi[1999:1984]},
     {maskSplit_maskSelect_hi[1983:1968]},
     {maskSplit_maskSelect_hi[1967:1952]},
     {maskSplit_maskSelect_hi[1951:1936]},
     {maskSplit_maskSelect_hi[1935:1920]},
     {maskSplit_maskSelect_hi[1919:1904]},
     {maskSplit_maskSelect_hi[1903:1888]},
     {maskSplit_maskSelect_hi[1887:1872]},
     {maskSplit_maskSelect_hi[1871:1856]},
     {maskSplit_maskSelect_hi[1855:1840]},
     {maskSplit_maskSelect_hi[1839:1824]},
     {maskSplit_maskSelect_hi[1823:1808]},
     {maskSplit_maskSelect_hi[1807:1792]},
     {maskSplit_maskSelect_hi[1791:1776]},
     {maskSplit_maskSelect_hi[1775:1760]},
     {maskSplit_maskSelect_hi[1759:1744]},
     {maskSplit_maskSelect_hi[1743:1728]},
     {maskSplit_maskSelect_hi[1727:1712]},
     {maskSplit_maskSelect_hi[1711:1696]},
     {maskSplit_maskSelect_hi[1695:1680]},
     {maskSplit_maskSelect_hi[1679:1664]},
     {maskSplit_maskSelect_hi[1663:1648]},
     {maskSplit_maskSelect_hi[1647:1632]},
     {maskSplit_maskSelect_hi[1631:1616]},
     {maskSplit_maskSelect_hi[1615:1600]},
     {maskSplit_maskSelect_hi[1599:1584]},
     {maskSplit_maskSelect_hi[1583:1568]},
     {maskSplit_maskSelect_hi[1567:1552]},
     {maskSplit_maskSelect_hi[1551:1536]},
     {maskSplit_maskSelect_hi[1535:1520]},
     {maskSplit_maskSelect_hi[1519:1504]},
     {maskSplit_maskSelect_hi[1503:1488]},
     {maskSplit_maskSelect_hi[1487:1472]},
     {maskSplit_maskSelect_hi[1471:1456]},
     {maskSplit_maskSelect_hi[1455:1440]},
     {maskSplit_maskSelect_hi[1439:1424]},
     {maskSplit_maskSelect_hi[1423:1408]},
     {maskSplit_maskSelect_hi[1407:1392]},
     {maskSplit_maskSelect_hi[1391:1376]},
     {maskSplit_maskSelect_hi[1375:1360]},
     {maskSplit_maskSelect_hi[1359:1344]},
     {maskSplit_maskSelect_hi[1343:1328]},
     {maskSplit_maskSelect_hi[1327:1312]},
     {maskSplit_maskSelect_hi[1311:1296]},
     {maskSplit_maskSelect_hi[1295:1280]},
     {maskSplit_maskSelect_hi[1279:1264]},
     {maskSplit_maskSelect_hi[1263:1248]},
     {maskSplit_maskSelect_hi[1247:1232]},
     {maskSplit_maskSelect_hi[1231:1216]},
     {maskSplit_maskSelect_hi[1215:1200]},
     {maskSplit_maskSelect_hi[1199:1184]},
     {maskSplit_maskSelect_hi[1183:1168]},
     {maskSplit_maskSelect_hi[1167:1152]},
     {maskSplit_maskSelect_hi[1151:1136]},
     {maskSplit_maskSelect_hi[1135:1120]},
     {maskSplit_maskSelect_hi[1119:1104]},
     {maskSplit_maskSelect_hi[1103:1088]},
     {maskSplit_maskSelect_hi[1087:1072]},
     {maskSplit_maskSelect_hi[1071:1056]},
     {maskSplit_maskSelect_hi[1055:1040]},
     {maskSplit_maskSelect_hi[1039:1024]},
     {maskSplit_maskSelect_hi[1023:1008]},
     {maskSplit_maskSelect_hi[1007:992]},
     {maskSplit_maskSelect_hi[991:976]},
     {maskSplit_maskSelect_hi[975:960]},
     {maskSplit_maskSelect_hi[959:944]},
     {maskSplit_maskSelect_hi[943:928]},
     {maskSplit_maskSelect_hi[927:912]},
     {maskSplit_maskSelect_hi[911:896]},
     {maskSplit_maskSelect_hi[895:880]},
     {maskSplit_maskSelect_hi[879:864]},
     {maskSplit_maskSelect_hi[863:848]},
     {maskSplit_maskSelect_hi[847:832]},
     {maskSplit_maskSelect_hi[831:816]},
     {maskSplit_maskSelect_hi[815:800]},
     {maskSplit_maskSelect_hi[799:784]},
     {maskSplit_maskSelect_hi[783:768]},
     {maskSplit_maskSelect_hi[767:752]},
     {maskSplit_maskSelect_hi[751:736]},
     {maskSplit_maskSelect_hi[735:720]},
     {maskSplit_maskSelect_hi[719:704]},
     {maskSplit_maskSelect_hi[703:688]},
     {maskSplit_maskSelect_hi[687:672]},
     {maskSplit_maskSelect_hi[671:656]},
     {maskSplit_maskSelect_hi[655:640]},
     {maskSplit_maskSelect_hi[639:624]},
     {maskSplit_maskSelect_hi[623:608]},
     {maskSplit_maskSelect_hi[607:592]},
     {maskSplit_maskSelect_hi[591:576]},
     {maskSplit_maskSelect_hi[575:560]},
     {maskSplit_maskSelect_hi[559:544]},
     {maskSplit_maskSelect_hi[543:528]},
     {maskSplit_maskSelect_hi[527:512]},
     {maskSplit_maskSelect_hi[511:496]},
     {maskSplit_maskSelect_hi[495:480]},
     {maskSplit_maskSelect_hi[479:464]},
     {maskSplit_maskSelect_hi[463:448]},
     {maskSplit_maskSelect_hi[447:432]},
     {maskSplit_maskSelect_hi[431:416]},
     {maskSplit_maskSelect_hi[415:400]},
     {maskSplit_maskSelect_hi[399:384]},
     {maskSplit_maskSelect_hi[383:368]},
     {maskSplit_maskSelect_hi[367:352]},
     {maskSplit_maskSelect_hi[351:336]},
     {maskSplit_maskSelect_hi[335:320]},
     {maskSplit_maskSelect_hi[319:304]},
     {maskSplit_maskSelect_hi[303:288]},
     {maskSplit_maskSelect_hi[287:272]},
     {maskSplit_maskSelect_hi[271:256]},
     {maskSplit_maskSelect_hi[255:240]},
     {maskSplit_maskSelect_hi[239:224]},
     {maskSplit_maskSelect_hi[223:208]},
     {maskSplit_maskSelect_hi[207:192]},
     {maskSplit_maskSelect_hi[191:176]},
     {maskSplit_maskSelect_hi[175:160]},
     {maskSplit_maskSelect_hi[159:144]},
     {maskSplit_maskSelect_hi[143:128]},
     {maskSplit_maskSelect_hi[127:112]},
     {maskSplit_maskSelect_hi[111:96]},
     {maskSplit_maskSelect_hi[95:80]},
     {maskSplit_maskSelect_hi[79:64]},
     {maskSplit_maskSelect_hi[63:48]},
     {maskSplit_maskSelect_hi[47:32]},
     {maskSplit_maskSelect_hi[31:16]},
     {maskSplit_maskSelect_hi[15:0]},
     {maskSplit_maskSelect_lo[4095:4080]},
     {maskSplit_maskSelect_lo[4079:4064]},
     {maskSplit_maskSelect_lo[4063:4048]},
     {maskSplit_maskSelect_lo[4047:4032]},
     {maskSplit_maskSelect_lo[4031:4016]},
     {maskSplit_maskSelect_lo[4015:4000]},
     {maskSplit_maskSelect_lo[3999:3984]},
     {maskSplit_maskSelect_lo[3983:3968]},
     {maskSplit_maskSelect_lo[3967:3952]},
     {maskSplit_maskSelect_lo[3951:3936]},
     {maskSplit_maskSelect_lo[3935:3920]},
     {maskSplit_maskSelect_lo[3919:3904]},
     {maskSplit_maskSelect_lo[3903:3888]},
     {maskSplit_maskSelect_lo[3887:3872]},
     {maskSplit_maskSelect_lo[3871:3856]},
     {maskSplit_maskSelect_lo[3855:3840]},
     {maskSplit_maskSelect_lo[3839:3824]},
     {maskSplit_maskSelect_lo[3823:3808]},
     {maskSplit_maskSelect_lo[3807:3792]},
     {maskSplit_maskSelect_lo[3791:3776]},
     {maskSplit_maskSelect_lo[3775:3760]},
     {maskSplit_maskSelect_lo[3759:3744]},
     {maskSplit_maskSelect_lo[3743:3728]},
     {maskSplit_maskSelect_lo[3727:3712]},
     {maskSplit_maskSelect_lo[3711:3696]},
     {maskSplit_maskSelect_lo[3695:3680]},
     {maskSplit_maskSelect_lo[3679:3664]},
     {maskSplit_maskSelect_lo[3663:3648]},
     {maskSplit_maskSelect_lo[3647:3632]},
     {maskSplit_maskSelect_lo[3631:3616]},
     {maskSplit_maskSelect_lo[3615:3600]},
     {maskSplit_maskSelect_lo[3599:3584]},
     {maskSplit_maskSelect_lo[3583:3568]},
     {maskSplit_maskSelect_lo[3567:3552]},
     {maskSplit_maskSelect_lo[3551:3536]},
     {maskSplit_maskSelect_lo[3535:3520]},
     {maskSplit_maskSelect_lo[3519:3504]},
     {maskSplit_maskSelect_lo[3503:3488]},
     {maskSplit_maskSelect_lo[3487:3472]},
     {maskSplit_maskSelect_lo[3471:3456]},
     {maskSplit_maskSelect_lo[3455:3440]},
     {maskSplit_maskSelect_lo[3439:3424]},
     {maskSplit_maskSelect_lo[3423:3408]},
     {maskSplit_maskSelect_lo[3407:3392]},
     {maskSplit_maskSelect_lo[3391:3376]},
     {maskSplit_maskSelect_lo[3375:3360]},
     {maskSplit_maskSelect_lo[3359:3344]},
     {maskSplit_maskSelect_lo[3343:3328]},
     {maskSplit_maskSelect_lo[3327:3312]},
     {maskSplit_maskSelect_lo[3311:3296]},
     {maskSplit_maskSelect_lo[3295:3280]},
     {maskSplit_maskSelect_lo[3279:3264]},
     {maskSplit_maskSelect_lo[3263:3248]},
     {maskSplit_maskSelect_lo[3247:3232]},
     {maskSplit_maskSelect_lo[3231:3216]},
     {maskSplit_maskSelect_lo[3215:3200]},
     {maskSplit_maskSelect_lo[3199:3184]},
     {maskSplit_maskSelect_lo[3183:3168]},
     {maskSplit_maskSelect_lo[3167:3152]},
     {maskSplit_maskSelect_lo[3151:3136]},
     {maskSplit_maskSelect_lo[3135:3120]},
     {maskSplit_maskSelect_lo[3119:3104]},
     {maskSplit_maskSelect_lo[3103:3088]},
     {maskSplit_maskSelect_lo[3087:3072]},
     {maskSplit_maskSelect_lo[3071:3056]},
     {maskSplit_maskSelect_lo[3055:3040]},
     {maskSplit_maskSelect_lo[3039:3024]},
     {maskSplit_maskSelect_lo[3023:3008]},
     {maskSplit_maskSelect_lo[3007:2992]},
     {maskSplit_maskSelect_lo[2991:2976]},
     {maskSplit_maskSelect_lo[2975:2960]},
     {maskSplit_maskSelect_lo[2959:2944]},
     {maskSplit_maskSelect_lo[2943:2928]},
     {maskSplit_maskSelect_lo[2927:2912]},
     {maskSplit_maskSelect_lo[2911:2896]},
     {maskSplit_maskSelect_lo[2895:2880]},
     {maskSplit_maskSelect_lo[2879:2864]},
     {maskSplit_maskSelect_lo[2863:2848]},
     {maskSplit_maskSelect_lo[2847:2832]},
     {maskSplit_maskSelect_lo[2831:2816]},
     {maskSplit_maskSelect_lo[2815:2800]},
     {maskSplit_maskSelect_lo[2799:2784]},
     {maskSplit_maskSelect_lo[2783:2768]},
     {maskSplit_maskSelect_lo[2767:2752]},
     {maskSplit_maskSelect_lo[2751:2736]},
     {maskSplit_maskSelect_lo[2735:2720]},
     {maskSplit_maskSelect_lo[2719:2704]},
     {maskSplit_maskSelect_lo[2703:2688]},
     {maskSplit_maskSelect_lo[2687:2672]},
     {maskSplit_maskSelect_lo[2671:2656]},
     {maskSplit_maskSelect_lo[2655:2640]},
     {maskSplit_maskSelect_lo[2639:2624]},
     {maskSplit_maskSelect_lo[2623:2608]},
     {maskSplit_maskSelect_lo[2607:2592]},
     {maskSplit_maskSelect_lo[2591:2576]},
     {maskSplit_maskSelect_lo[2575:2560]},
     {maskSplit_maskSelect_lo[2559:2544]},
     {maskSplit_maskSelect_lo[2543:2528]},
     {maskSplit_maskSelect_lo[2527:2512]},
     {maskSplit_maskSelect_lo[2511:2496]},
     {maskSplit_maskSelect_lo[2495:2480]},
     {maskSplit_maskSelect_lo[2479:2464]},
     {maskSplit_maskSelect_lo[2463:2448]},
     {maskSplit_maskSelect_lo[2447:2432]},
     {maskSplit_maskSelect_lo[2431:2416]},
     {maskSplit_maskSelect_lo[2415:2400]},
     {maskSplit_maskSelect_lo[2399:2384]},
     {maskSplit_maskSelect_lo[2383:2368]},
     {maskSplit_maskSelect_lo[2367:2352]},
     {maskSplit_maskSelect_lo[2351:2336]},
     {maskSplit_maskSelect_lo[2335:2320]},
     {maskSplit_maskSelect_lo[2319:2304]},
     {maskSplit_maskSelect_lo[2303:2288]},
     {maskSplit_maskSelect_lo[2287:2272]},
     {maskSplit_maskSelect_lo[2271:2256]},
     {maskSplit_maskSelect_lo[2255:2240]},
     {maskSplit_maskSelect_lo[2239:2224]},
     {maskSplit_maskSelect_lo[2223:2208]},
     {maskSplit_maskSelect_lo[2207:2192]},
     {maskSplit_maskSelect_lo[2191:2176]},
     {maskSplit_maskSelect_lo[2175:2160]},
     {maskSplit_maskSelect_lo[2159:2144]},
     {maskSplit_maskSelect_lo[2143:2128]},
     {maskSplit_maskSelect_lo[2127:2112]},
     {maskSplit_maskSelect_lo[2111:2096]},
     {maskSplit_maskSelect_lo[2095:2080]},
     {maskSplit_maskSelect_lo[2079:2064]},
     {maskSplit_maskSelect_lo[2063:2048]},
     {maskSplit_maskSelect_lo[2047:2032]},
     {maskSplit_maskSelect_lo[2031:2016]},
     {maskSplit_maskSelect_lo[2015:2000]},
     {maskSplit_maskSelect_lo[1999:1984]},
     {maskSplit_maskSelect_lo[1983:1968]},
     {maskSplit_maskSelect_lo[1967:1952]},
     {maskSplit_maskSelect_lo[1951:1936]},
     {maskSplit_maskSelect_lo[1935:1920]},
     {maskSplit_maskSelect_lo[1919:1904]},
     {maskSplit_maskSelect_lo[1903:1888]},
     {maskSplit_maskSelect_lo[1887:1872]},
     {maskSplit_maskSelect_lo[1871:1856]},
     {maskSplit_maskSelect_lo[1855:1840]},
     {maskSplit_maskSelect_lo[1839:1824]},
     {maskSplit_maskSelect_lo[1823:1808]},
     {maskSplit_maskSelect_lo[1807:1792]},
     {maskSplit_maskSelect_lo[1791:1776]},
     {maskSplit_maskSelect_lo[1775:1760]},
     {maskSplit_maskSelect_lo[1759:1744]},
     {maskSplit_maskSelect_lo[1743:1728]},
     {maskSplit_maskSelect_lo[1727:1712]},
     {maskSplit_maskSelect_lo[1711:1696]},
     {maskSplit_maskSelect_lo[1695:1680]},
     {maskSplit_maskSelect_lo[1679:1664]},
     {maskSplit_maskSelect_lo[1663:1648]},
     {maskSplit_maskSelect_lo[1647:1632]},
     {maskSplit_maskSelect_lo[1631:1616]},
     {maskSplit_maskSelect_lo[1615:1600]},
     {maskSplit_maskSelect_lo[1599:1584]},
     {maskSplit_maskSelect_lo[1583:1568]},
     {maskSplit_maskSelect_lo[1567:1552]},
     {maskSplit_maskSelect_lo[1551:1536]},
     {maskSplit_maskSelect_lo[1535:1520]},
     {maskSplit_maskSelect_lo[1519:1504]},
     {maskSplit_maskSelect_lo[1503:1488]},
     {maskSplit_maskSelect_lo[1487:1472]},
     {maskSplit_maskSelect_lo[1471:1456]},
     {maskSplit_maskSelect_lo[1455:1440]},
     {maskSplit_maskSelect_lo[1439:1424]},
     {maskSplit_maskSelect_lo[1423:1408]},
     {maskSplit_maskSelect_lo[1407:1392]},
     {maskSplit_maskSelect_lo[1391:1376]},
     {maskSplit_maskSelect_lo[1375:1360]},
     {maskSplit_maskSelect_lo[1359:1344]},
     {maskSplit_maskSelect_lo[1343:1328]},
     {maskSplit_maskSelect_lo[1327:1312]},
     {maskSplit_maskSelect_lo[1311:1296]},
     {maskSplit_maskSelect_lo[1295:1280]},
     {maskSplit_maskSelect_lo[1279:1264]},
     {maskSplit_maskSelect_lo[1263:1248]},
     {maskSplit_maskSelect_lo[1247:1232]},
     {maskSplit_maskSelect_lo[1231:1216]},
     {maskSplit_maskSelect_lo[1215:1200]},
     {maskSplit_maskSelect_lo[1199:1184]},
     {maskSplit_maskSelect_lo[1183:1168]},
     {maskSplit_maskSelect_lo[1167:1152]},
     {maskSplit_maskSelect_lo[1151:1136]},
     {maskSplit_maskSelect_lo[1135:1120]},
     {maskSplit_maskSelect_lo[1119:1104]},
     {maskSplit_maskSelect_lo[1103:1088]},
     {maskSplit_maskSelect_lo[1087:1072]},
     {maskSplit_maskSelect_lo[1071:1056]},
     {maskSplit_maskSelect_lo[1055:1040]},
     {maskSplit_maskSelect_lo[1039:1024]},
     {maskSplit_maskSelect_lo[1023:1008]},
     {maskSplit_maskSelect_lo[1007:992]},
     {maskSplit_maskSelect_lo[991:976]},
     {maskSplit_maskSelect_lo[975:960]},
     {maskSplit_maskSelect_lo[959:944]},
     {maskSplit_maskSelect_lo[943:928]},
     {maskSplit_maskSelect_lo[927:912]},
     {maskSplit_maskSelect_lo[911:896]},
     {maskSplit_maskSelect_lo[895:880]},
     {maskSplit_maskSelect_lo[879:864]},
     {maskSplit_maskSelect_lo[863:848]},
     {maskSplit_maskSelect_lo[847:832]},
     {maskSplit_maskSelect_lo[831:816]},
     {maskSplit_maskSelect_lo[815:800]},
     {maskSplit_maskSelect_lo[799:784]},
     {maskSplit_maskSelect_lo[783:768]},
     {maskSplit_maskSelect_lo[767:752]},
     {maskSplit_maskSelect_lo[751:736]},
     {maskSplit_maskSelect_lo[735:720]},
     {maskSplit_maskSelect_lo[719:704]},
     {maskSplit_maskSelect_lo[703:688]},
     {maskSplit_maskSelect_lo[687:672]},
     {maskSplit_maskSelect_lo[671:656]},
     {maskSplit_maskSelect_lo[655:640]},
     {maskSplit_maskSelect_lo[639:624]},
     {maskSplit_maskSelect_lo[623:608]},
     {maskSplit_maskSelect_lo[607:592]},
     {maskSplit_maskSelect_lo[591:576]},
     {maskSplit_maskSelect_lo[575:560]},
     {maskSplit_maskSelect_lo[559:544]},
     {maskSplit_maskSelect_lo[543:528]},
     {maskSplit_maskSelect_lo[527:512]},
     {maskSplit_maskSelect_lo[511:496]},
     {maskSplit_maskSelect_lo[495:480]},
     {maskSplit_maskSelect_lo[479:464]},
     {maskSplit_maskSelect_lo[463:448]},
     {maskSplit_maskSelect_lo[447:432]},
     {maskSplit_maskSelect_lo[431:416]},
     {maskSplit_maskSelect_lo[415:400]},
     {maskSplit_maskSelect_lo[399:384]},
     {maskSplit_maskSelect_lo[383:368]},
     {maskSplit_maskSelect_lo[367:352]},
     {maskSplit_maskSelect_lo[351:336]},
     {maskSplit_maskSelect_lo[335:320]},
     {maskSplit_maskSelect_lo[319:304]},
     {maskSplit_maskSelect_lo[303:288]},
     {maskSplit_maskSelect_lo[287:272]},
     {maskSplit_maskSelect_lo[271:256]},
     {maskSplit_maskSelect_lo[255:240]},
     {maskSplit_maskSelect_lo[239:224]},
     {maskSplit_maskSelect_lo[223:208]},
     {maskSplit_maskSelect_lo[207:192]},
     {maskSplit_maskSelect_lo[191:176]},
     {maskSplit_maskSelect_lo[175:160]},
     {maskSplit_maskSelect_lo[159:144]},
     {maskSplit_maskSelect_lo[143:128]},
     {maskSplit_maskSelect_lo[127:112]},
     {maskSplit_maskSelect_lo[111:96]},
     {maskSplit_maskSelect_lo[95:80]},
     {maskSplit_maskSelect_lo[79:64]},
     {maskSplit_maskSelect_lo[63:48]},
     {maskSplit_maskSelect_lo[47:32]},
     {maskSplit_maskSelect_lo[31:16]},
     {maskSplit_maskSelect_lo[15:0]}};
  wire [15:0]        maskSplit_0_2 = (instReg_maskType ? _GEN_143[executeGroupCounter[8:0]] : 16'hFFFF) & maskSplit_vlBoundaryCorrection;
  wire [1:0]         maskSplit_byteMask_lo_lo_lo = maskSplit_0_2[1:0];
  wire [1:0]         maskSplit_byteMask_lo_lo_hi = maskSplit_0_2[3:2];
  wire [3:0]         maskSplit_byteMask_lo_lo = {maskSplit_byteMask_lo_lo_hi, maskSplit_byteMask_lo_lo_lo};
  wire [1:0]         maskSplit_byteMask_lo_hi_lo = maskSplit_0_2[5:4];
  wire [1:0]         maskSplit_byteMask_lo_hi_hi = maskSplit_0_2[7:6];
  wire [3:0]         maskSplit_byteMask_lo_hi = {maskSplit_byteMask_lo_hi_hi, maskSplit_byteMask_lo_hi_lo};
  wire [7:0]         maskSplit_byteMask_lo = {maskSplit_byteMask_lo_hi, maskSplit_byteMask_lo_lo};
  wire [1:0]         maskSplit_byteMask_hi_lo_lo = maskSplit_0_2[9:8];
  wire [1:0]         maskSplit_byteMask_hi_lo_hi = maskSplit_0_2[11:10];
  wire [3:0]         maskSplit_byteMask_hi_lo = {maskSplit_byteMask_hi_lo_hi, maskSplit_byteMask_hi_lo_lo};
  wire [1:0]         maskSplit_byteMask_hi_hi_lo = maskSplit_0_2[13:12];
  wire [1:0]         maskSplit_byteMask_hi_hi_hi = maskSplit_0_2[15:14];
  wire [3:0]         maskSplit_byteMask_hi_hi = {maskSplit_byteMask_hi_hi_hi, maskSplit_byteMask_hi_hi_lo};
  wire [7:0]         maskSplit_byteMask_hi = {maskSplit_byteMask_hi_hi, maskSplit_byteMask_hi_lo};
  wire [15:0]        maskSplit_0_1 = {maskSplit_byteMask_hi, maskSplit_byteMask_lo};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_lo_lo_lo_1 = {maskSplit_maskSelect_lo_lo_lo_lo_lo_lo_hi_1, maskSplit_maskSelect_lo_lo_lo_lo_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_lo_lo_hi_1 = {maskSplit_maskSelect_lo_lo_lo_lo_lo_hi_hi_1, maskSplit_maskSelect_lo_lo_lo_lo_lo_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_lo_lo_lo_lo_lo_1 = {maskSplit_maskSelect_lo_lo_lo_lo_lo_hi_1, maskSplit_maskSelect_lo_lo_lo_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_lo_hi_lo_1 = {maskSplit_maskSelect_lo_lo_lo_lo_hi_lo_hi_1, maskSplit_maskSelect_lo_lo_lo_lo_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_lo_hi_hi_1 = {maskSplit_maskSelect_lo_lo_lo_lo_hi_hi_hi_1, maskSplit_maskSelect_lo_lo_lo_lo_hi_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_lo_lo_lo_lo_hi_1 = {maskSplit_maskSelect_lo_lo_lo_lo_hi_hi_1, maskSplit_maskSelect_lo_lo_lo_lo_hi_lo_1};
  wire [511:0]       maskSplit_maskSelect_lo_lo_lo_lo_1 = {maskSplit_maskSelect_lo_lo_lo_lo_hi_1, maskSplit_maskSelect_lo_lo_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_hi_lo_lo_1 = {maskSplit_maskSelect_lo_lo_lo_hi_lo_lo_hi_1, maskSplit_maskSelect_lo_lo_lo_hi_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_hi_lo_hi_1 = {maskSplit_maskSelect_lo_lo_lo_hi_lo_hi_hi_1, maskSplit_maskSelect_lo_lo_lo_hi_lo_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_lo_lo_lo_hi_lo_1 = {maskSplit_maskSelect_lo_lo_lo_hi_lo_hi_1, maskSplit_maskSelect_lo_lo_lo_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_hi_hi_lo_1 = {maskSplit_maskSelect_lo_lo_lo_hi_hi_lo_hi_1, maskSplit_maskSelect_lo_lo_lo_hi_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_hi_hi_hi_1 = {maskSplit_maskSelect_lo_lo_lo_hi_hi_hi_hi_1, maskSplit_maskSelect_lo_lo_lo_hi_hi_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_lo_lo_lo_hi_hi_1 = {maskSplit_maskSelect_lo_lo_lo_hi_hi_hi_1, maskSplit_maskSelect_lo_lo_lo_hi_hi_lo_1};
  wire [511:0]       maskSplit_maskSelect_lo_lo_lo_hi_1 = {maskSplit_maskSelect_lo_lo_lo_hi_hi_1, maskSplit_maskSelect_lo_lo_lo_hi_lo_1};
  wire [1023:0]      maskSplit_maskSelect_lo_lo_lo_1 = {maskSplit_maskSelect_lo_lo_lo_hi_1, maskSplit_maskSelect_lo_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_lo_lo_lo_1 = {maskSplit_maskSelect_lo_lo_hi_lo_lo_lo_hi_1, maskSplit_maskSelect_lo_lo_hi_lo_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_lo_lo_hi_1 = {maskSplit_maskSelect_lo_lo_hi_lo_lo_hi_hi_1, maskSplit_maskSelect_lo_lo_hi_lo_lo_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_lo_lo_hi_lo_lo_1 = {maskSplit_maskSelect_lo_lo_hi_lo_lo_hi_1, maskSplit_maskSelect_lo_lo_hi_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_lo_hi_lo_1 = {maskSplit_maskSelect_lo_lo_hi_lo_hi_lo_hi_1, maskSplit_maskSelect_lo_lo_hi_lo_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_lo_hi_hi_1 = {maskSplit_maskSelect_lo_lo_hi_lo_hi_hi_hi_1, maskSplit_maskSelect_lo_lo_hi_lo_hi_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_lo_lo_hi_lo_hi_1 = {maskSplit_maskSelect_lo_lo_hi_lo_hi_hi_1, maskSplit_maskSelect_lo_lo_hi_lo_hi_lo_1};
  wire [511:0]       maskSplit_maskSelect_lo_lo_hi_lo_1 = {maskSplit_maskSelect_lo_lo_hi_lo_hi_1, maskSplit_maskSelect_lo_lo_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_hi_lo_lo_1 = {maskSplit_maskSelect_lo_lo_hi_hi_lo_lo_hi_1, maskSplit_maskSelect_lo_lo_hi_hi_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_hi_lo_hi_1 = {maskSplit_maskSelect_lo_lo_hi_hi_lo_hi_hi_1, maskSplit_maskSelect_lo_lo_hi_hi_lo_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_lo_lo_hi_hi_lo_1 = {maskSplit_maskSelect_lo_lo_hi_hi_lo_hi_1, maskSplit_maskSelect_lo_lo_hi_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_hi_hi_lo_1 = {maskSplit_maskSelect_lo_lo_hi_hi_hi_lo_hi_1, maskSplit_maskSelect_lo_lo_hi_hi_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_hi_hi_hi_1 = {maskSplit_maskSelect_lo_lo_hi_hi_hi_hi_hi_1, maskSplit_maskSelect_lo_lo_hi_hi_hi_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_lo_lo_hi_hi_hi_1 = {maskSplit_maskSelect_lo_lo_hi_hi_hi_hi_1, maskSplit_maskSelect_lo_lo_hi_hi_hi_lo_1};
  wire [511:0]       maskSplit_maskSelect_lo_lo_hi_hi_1 = {maskSplit_maskSelect_lo_lo_hi_hi_hi_1, maskSplit_maskSelect_lo_lo_hi_hi_lo_1};
  wire [1023:0]      maskSplit_maskSelect_lo_lo_hi_1 = {maskSplit_maskSelect_lo_lo_hi_hi_1, maskSplit_maskSelect_lo_lo_hi_lo_1};
  wire [2047:0]      maskSplit_maskSelect_lo_lo_1 = {maskSplit_maskSelect_lo_lo_hi_1, maskSplit_maskSelect_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_lo_lo_lo_1 = {maskSplit_maskSelect_lo_hi_lo_lo_lo_lo_hi_1, maskSplit_maskSelect_lo_hi_lo_lo_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_lo_lo_hi_1 = {maskSplit_maskSelect_lo_hi_lo_lo_lo_hi_hi_1, maskSplit_maskSelect_lo_hi_lo_lo_lo_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_lo_hi_lo_lo_lo_1 = {maskSplit_maskSelect_lo_hi_lo_lo_lo_hi_1, maskSplit_maskSelect_lo_hi_lo_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_lo_hi_lo_1 = {maskSplit_maskSelect_lo_hi_lo_lo_hi_lo_hi_1, maskSplit_maskSelect_lo_hi_lo_lo_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_lo_hi_hi_1 = {maskSplit_maskSelect_lo_hi_lo_lo_hi_hi_hi_1, maskSplit_maskSelect_lo_hi_lo_lo_hi_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_lo_hi_lo_lo_hi_1 = {maskSplit_maskSelect_lo_hi_lo_lo_hi_hi_1, maskSplit_maskSelect_lo_hi_lo_lo_hi_lo_1};
  wire [511:0]       maskSplit_maskSelect_lo_hi_lo_lo_1 = {maskSplit_maskSelect_lo_hi_lo_lo_hi_1, maskSplit_maskSelect_lo_hi_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_hi_lo_lo_1 = {maskSplit_maskSelect_lo_hi_lo_hi_lo_lo_hi_1, maskSplit_maskSelect_lo_hi_lo_hi_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_hi_lo_hi_1 = {maskSplit_maskSelect_lo_hi_lo_hi_lo_hi_hi_1, maskSplit_maskSelect_lo_hi_lo_hi_lo_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_lo_hi_lo_hi_lo_1 = {maskSplit_maskSelect_lo_hi_lo_hi_lo_hi_1, maskSplit_maskSelect_lo_hi_lo_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_hi_hi_lo_1 = {maskSplit_maskSelect_lo_hi_lo_hi_hi_lo_hi_1, maskSplit_maskSelect_lo_hi_lo_hi_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_hi_hi_hi_1 = {maskSplit_maskSelect_lo_hi_lo_hi_hi_hi_hi_1, maskSplit_maskSelect_lo_hi_lo_hi_hi_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_lo_hi_lo_hi_hi_1 = {maskSplit_maskSelect_lo_hi_lo_hi_hi_hi_1, maskSplit_maskSelect_lo_hi_lo_hi_hi_lo_1};
  wire [511:0]       maskSplit_maskSelect_lo_hi_lo_hi_1 = {maskSplit_maskSelect_lo_hi_lo_hi_hi_1, maskSplit_maskSelect_lo_hi_lo_hi_lo_1};
  wire [1023:0]      maskSplit_maskSelect_lo_hi_lo_1 = {maskSplit_maskSelect_lo_hi_lo_hi_1, maskSplit_maskSelect_lo_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_lo_lo_lo_1 = {maskSplit_maskSelect_lo_hi_hi_lo_lo_lo_hi_1, maskSplit_maskSelect_lo_hi_hi_lo_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_lo_lo_hi_1 = {maskSplit_maskSelect_lo_hi_hi_lo_lo_hi_hi_1, maskSplit_maskSelect_lo_hi_hi_lo_lo_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_lo_hi_hi_lo_lo_1 = {maskSplit_maskSelect_lo_hi_hi_lo_lo_hi_1, maskSplit_maskSelect_lo_hi_hi_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_lo_hi_lo_1 = {maskSplit_maskSelect_lo_hi_hi_lo_hi_lo_hi_1, maskSplit_maskSelect_lo_hi_hi_lo_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_lo_hi_hi_1 = {maskSplit_maskSelect_lo_hi_hi_lo_hi_hi_hi_1, maskSplit_maskSelect_lo_hi_hi_lo_hi_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_lo_hi_hi_lo_hi_1 = {maskSplit_maskSelect_lo_hi_hi_lo_hi_hi_1, maskSplit_maskSelect_lo_hi_hi_lo_hi_lo_1};
  wire [511:0]       maskSplit_maskSelect_lo_hi_hi_lo_1 = {maskSplit_maskSelect_lo_hi_hi_lo_hi_1, maskSplit_maskSelect_lo_hi_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_hi_lo_lo_1 = {maskSplit_maskSelect_lo_hi_hi_hi_lo_lo_hi_1, maskSplit_maskSelect_lo_hi_hi_hi_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_hi_lo_hi_1 = {maskSplit_maskSelect_lo_hi_hi_hi_lo_hi_hi_1, maskSplit_maskSelect_lo_hi_hi_hi_lo_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_lo_hi_hi_hi_lo_1 = {maskSplit_maskSelect_lo_hi_hi_hi_lo_hi_1, maskSplit_maskSelect_lo_hi_hi_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_hi_hi_lo_1 = {maskSplit_maskSelect_lo_hi_hi_hi_hi_lo_hi_1, maskSplit_maskSelect_lo_hi_hi_hi_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_hi_hi_hi_1 = {maskSplit_maskSelect_lo_hi_hi_hi_hi_hi_hi_1, maskSplit_maskSelect_lo_hi_hi_hi_hi_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_lo_hi_hi_hi_hi_1 = {maskSplit_maskSelect_lo_hi_hi_hi_hi_hi_1, maskSplit_maskSelect_lo_hi_hi_hi_hi_lo_1};
  wire [511:0]       maskSplit_maskSelect_lo_hi_hi_hi_1 = {maskSplit_maskSelect_lo_hi_hi_hi_hi_1, maskSplit_maskSelect_lo_hi_hi_hi_lo_1};
  wire [1023:0]      maskSplit_maskSelect_lo_hi_hi_1 = {maskSplit_maskSelect_lo_hi_hi_hi_1, maskSplit_maskSelect_lo_hi_hi_lo_1};
  wire [2047:0]      maskSplit_maskSelect_lo_hi_1 = {maskSplit_maskSelect_lo_hi_hi_1, maskSplit_maskSelect_lo_hi_lo_1};
  wire [4095:0]      maskSplit_maskSelect_lo_1 = {maskSplit_maskSelect_lo_hi_1, maskSplit_maskSelect_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_lo_lo_lo_1 = {maskSplit_maskSelect_hi_lo_lo_lo_lo_lo_hi_1, maskSplit_maskSelect_hi_lo_lo_lo_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_lo_lo_hi_1 = {maskSplit_maskSelect_hi_lo_lo_lo_lo_hi_hi_1, maskSplit_maskSelect_hi_lo_lo_lo_lo_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_hi_lo_lo_lo_lo_1 = {maskSplit_maskSelect_hi_lo_lo_lo_lo_hi_1, maskSplit_maskSelect_hi_lo_lo_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_lo_hi_lo_1 = {maskSplit_maskSelect_hi_lo_lo_lo_hi_lo_hi_1, maskSplit_maskSelect_hi_lo_lo_lo_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_lo_hi_hi_1 = {maskSplit_maskSelect_hi_lo_lo_lo_hi_hi_hi_1, maskSplit_maskSelect_hi_lo_lo_lo_hi_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_hi_lo_lo_lo_hi_1 = {maskSplit_maskSelect_hi_lo_lo_lo_hi_hi_1, maskSplit_maskSelect_hi_lo_lo_lo_hi_lo_1};
  wire [511:0]       maskSplit_maskSelect_hi_lo_lo_lo_1 = {maskSplit_maskSelect_hi_lo_lo_lo_hi_1, maskSplit_maskSelect_hi_lo_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_hi_lo_lo_1 = {maskSplit_maskSelect_hi_lo_lo_hi_lo_lo_hi_1, maskSplit_maskSelect_hi_lo_lo_hi_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_hi_lo_hi_1 = {maskSplit_maskSelect_hi_lo_lo_hi_lo_hi_hi_1, maskSplit_maskSelect_hi_lo_lo_hi_lo_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_hi_lo_lo_hi_lo_1 = {maskSplit_maskSelect_hi_lo_lo_hi_lo_hi_1, maskSplit_maskSelect_hi_lo_lo_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_hi_hi_lo_1 = {maskSplit_maskSelect_hi_lo_lo_hi_hi_lo_hi_1, maskSplit_maskSelect_hi_lo_lo_hi_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_hi_hi_hi_1 = {maskSplit_maskSelect_hi_lo_lo_hi_hi_hi_hi_1, maskSplit_maskSelect_hi_lo_lo_hi_hi_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_hi_lo_lo_hi_hi_1 = {maskSplit_maskSelect_hi_lo_lo_hi_hi_hi_1, maskSplit_maskSelect_hi_lo_lo_hi_hi_lo_1};
  wire [511:0]       maskSplit_maskSelect_hi_lo_lo_hi_1 = {maskSplit_maskSelect_hi_lo_lo_hi_hi_1, maskSplit_maskSelect_hi_lo_lo_hi_lo_1};
  wire [1023:0]      maskSplit_maskSelect_hi_lo_lo_1 = {maskSplit_maskSelect_hi_lo_lo_hi_1, maskSplit_maskSelect_hi_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_lo_lo_lo_1 = {maskSplit_maskSelect_hi_lo_hi_lo_lo_lo_hi_1, maskSplit_maskSelect_hi_lo_hi_lo_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_lo_lo_hi_1 = {maskSplit_maskSelect_hi_lo_hi_lo_lo_hi_hi_1, maskSplit_maskSelect_hi_lo_hi_lo_lo_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_hi_lo_hi_lo_lo_1 = {maskSplit_maskSelect_hi_lo_hi_lo_lo_hi_1, maskSplit_maskSelect_hi_lo_hi_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_lo_hi_lo_1 = {maskSplit_maskSelect_hi_lo_hi_lo_hi_lo_hi_1, maskSplit_maskSelect_hi_lo_hi_lo_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_lo_hi_hi_1 = {maskSplit_maskSelect_hi_lo_hi_lo_hi_hi_hi_1, maskSplit_maskSelect_hi_lo_hi_lo_hi_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_hi_lo_hi_lo_hi_1 = {maskSplit_maskSelect_hi_lo_hi_lo_hi_hi_1, maskSplit_maskSelect_hi_lo_hi_lo_hi_lo_1};
  wire [511:0]       maskSplit_maskSelect_hi_lo_hi_lo_1 = {maskSplit_maskSelect_hi_lo_hi_lo_hi_1, maskSplit_maskSelect_hi_lo_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_hi_lo_lo_1 = {maskSplit_maskSelect_hi_lo_hi_hi_lo_lo_hi_1, maskSplit_maskSelect_hi_lo_hi_hi_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_hi_lo_hi_1 = {maskSplit_maskSelect_hi_lo_hi_hi_lo_hi_hi_1, maskSplit_maskSelect_hi_lo_hi_hi_lo_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_hi_lo_hi_hi_lo_1 = {maskSplit_maskSelect_hi_lo_hi_hi_lo_hi_1, maskSplit_maskSelect_hi_lo_hi_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_hi_hi_lo_1 = {maskSplit_maskSelect_hi_lo_hi_hi_hi_lo_hi_1, maskSplit_maskSelect_hi_lo_hi_hi_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_hi_hi_hi_1 = {maskSplit_maskSelect_hi_lo_hi_hi_hi_hi_hi_1, maskSplit_maskSelect_hi_lo_hi_hi_hi_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_hi_lo_hi_hi_hi_1 = {maskSplit_maskSelect_hi_lo_hi_hi_hi_hi_1, maskSplit_maskSelect_hi_lo_hi_hi_hi_lo_1};
  wire [511:0]       maskSplit_maskSelect_hi_lo_hi_hi_1 = {maskSplit_maskSelect_hi_lo_hi_hi_hi_1, maskSplit_maskSelect_hi_lo_hi_hi_lo_1};
  wire [1023:0]      maskSplit_maskSelect_hi_lo_hi_1 = {maskSplit_maskSelect_hi_lo_hi_hi_1, maskSplit_maskSelect_hi_lo_hi_lo_1};
  wire [2047:0]      maskSplit_maskSelect_hi_lo_1 = {maskSplit_maskSelect_hi_lo_hi_1, maskSplit_maskSelect_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_lo_lo_lo_1 = {maskSplit_maskSelect_hi_hi_lo_lo_lo_lo_hi_1, maskSplit_maskSelect_hi_hi_lo_lo_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_lo_lo_hi_1 = {maskSplit_maskSelect_hi_hi_lo_lo_lo_hi_hi_1, maskSplit_maskSelect_hi_hi_lo_lo_lo_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_hi_hi_lo_lo_lo_1 = {maskSplit_maskSelect_hi_hi_lo_lo_lo_hi_1, maskSplit_maskSelect_hi_hi_lo_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_lo_hi_lo_1 = {maskSplit_maskSelect_hi_hi_lo_lo_hi_lo_hi_1, maskSplit_maskSelect_hi_hi_lo_lo_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_lo_hi_hi_1 = {maskSplit_maskSelect_hi_hi_lo_lo_hi_hi_hi_1, maskSplit_maskSelect_hi_hi_lo_lo_hi_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_hi_hi_lo_lo_hi_1 = {maskSplit_maskSelect_hi_hi_lo_lo_hi_hi_1, maskSplit_maskSelect_hi_hi_lo_lo_hi_lo_1};
  wire [511:0]       maskSplit_maskSelect_hi_hi_lo_lo_1 = {maskSplit_maskSelect_hi_hi_lo_lo_hi_1, maskSplit_maskSelect_hi_hi_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_hi_lo_lo_1 = {maskSplit_maskSelect_hi_hi_lo_hi_lo_lo_hi_1, maskSplit_maskSelect_hi_hi_lo_hi_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_hi_lo_hi_1 = {maskSplit_maskSelect_hi_hi_lo_hi_lo_hi_hi_1, maskSplit_maskSelect_hi_hi_lo_hi_lo_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_hi_hi_lo_hi_lo_1 = {maskSplit_maskSelect_hi_hi_lo_hi_lo_hi_1, maskSplit_maskSelect_hi_hi_lo_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_hi_hi_lo_1 = {maskSplit_maskSelect_hi_hi_lo_hi_hi_lo_hi_1, maskSplit_maskSelect_hi_hi_lo_hi_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_hi_hi_hi_1 = {maskSplit_maskSelect_hi_hi_lo_hi_hi_hi_hi_1, maskSplit_maskSelect_hi_hi_lo_hi_hi_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_hi_hi_lo_hi_hi_1 = {maskSplit_maskSelect_hi_hi_lo_hi_hi_hi_1, maskSplit_maskSelect_hi_hi_lo_hi_hi_lo_1};
  wire [511:0]       maskSplit_maskSelect_hi_hi_lo_hi_1 = {maskSplit_maskSelect_hi_hi_lo_hi_hi_1, maskSplit_maskSelect_hi_hi_lo_hi_lo_1};
  wire [1023:0]      maskSplit_maskSelect_hi_hi_lo_1 = {maskSplit_maskSelect_hi_hi_lo_hi_1, maskSplit_maskSelect_hi_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_lo_lo_lo_1 = {maskSplit_maskSelect_hi_hi_hi_lo_lo_lo_hi_1, maskSplit_maskSelect_hi_hi_hi_lo_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_lo_lo_hi_1 = {maskSplit_maskSelect_hi_hi_hi_lo_lo_hi_hi_1, maskSplit_maskSelect_hi_hi_hi_lo_lo_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_hi_hi_hi_lo_lo_1 = {maskSplit_maskSelect_hi_hi_hi_lo_lo_hi_1, maskSplit_maskSelect_hi_hi_hi_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_lo_hi_lo_1 = {maskSplit_maskSelect_hi_hi_hi_lo_hi_lo_hi_1, maskSplit_maskSelect_hi_hi_hi_lo_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_lo_hi_hi_1 = {maskSplit_maskSelect_hi_hi_hi_lo_hi_hi_hi_1, maskSplit_maskSelect_hi_hi_hi_lo_hi_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_hi_hi_hi_lo_hi_1 = {maskSplit_maskSelect_hi_hi_hi_lo_hi_hi_1, maskSplit_maskSelect_hi_hi_hi_lo_hi_lo_1};
  wire [511:0]       maskSplit_maskSelect_hi_hi_hi_lo_1 = {maskSplit_maskSelect_hi_hi_hi_lo_hi_1, maskSplit_maskSelect_hi_hi_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_hi_lo_lo_1 = {maskSplit_maskSelect_hi_hi_hi_hi_lo_lo_hi_1, maskSplit_maskSelect_hi_hi_hi_hi_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_hi_lo_hi_1 = {maskSplit_maskSelect_hi_hi_hi_hi_lo_hi_hi_1, maskSplit_maskSelect_hi_hi_hi_hi_lo_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_hi_hi_hi_hi_lo_1 = {maskSplit_maskSelect_hi_hi_hi_hi_lo_hi_1, maskSplit_maskSelect_hi_hi_hi_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_hi_hi_lo_1 = {maskSplit_maskSelect_hi_hi_hi_hi_hi_lo_hi_1, maskSplit_maskSelect_hi_hi_hi_hi_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_hi_hi_hi_1 = {maskSplit_maskSelect_hi_hi_hi_hi_hi_hi_hi_1, maskSplit_maskSelect_hi_hi_hi_hi_hi_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_hi_hi_hi_hi_hi_1 = {maskSplit_maskSelect_hi_hi_hi_hi_hi_hi_1, maskSplit_maskSelect_hi_hi_hi_hi_hi_lo_1};
  wire [511:0]       maskSplit_maskSelect_hi_hi_hi_hi_1 = {maskSplit_maskSelect_hi_hi_hi_hi_hi_1, maskSplit_maskSelect_hi_hi_hi_hi_lo_1};
  wire [1023:0]      maskSplit_maskSelect_hi_hi_hi_1 = {maskSplit_maskSelect_hi_hi_hi_hi_1, maskSplit_maskSelect_hi_hi_hi_lo_1};
  wire [2047:0]      maskSplit_maskSelect_hi_hi_1 = {maskSplit_maskSelect_hi_hi_hi_1, maskSplit_maskSelect_hi_hi_lo_1};
  wire [4095:0]      maskSplit_maskSelect_hi_1 = {maskSplit_maskSelect_hi_hi_1, maskSplit_maskSelect_hi_lo_1};
  wire               maskSplit_vlMisAlign_1 = |(instReg_vl[2:0]);
  wire [10:0]        maskSplit_lastexecuteGroup_1 = instReg_vl[13:3] - {10'h0, ~maskSplit_vlMisAlign_1};
  wire [10:0]        _GEN_144 = {1'h0, executeGroupCounter};
  wire               maskSplit_isVlBoundary_1 = _GEN_144 == maskSplit_lastexecuteGroup_1;
  wire               maskSplit_validExecuteGroup_1 = _GEN_144 <= maskSplit_lastexecuteGroup_1;
  wire [7:0]         _maskSplit_vlBoundaryCorrection_T_21 = 8'h1 << instReg_vl[2:0];
  wire [7:0]         _maskSplit_vlBoundaryCorrection_T_24 = _maskSplit_vlBoundaryCorrection_T_21 | {_maskSplit_vlBoundaryCorrection_T_21[6:0], 1'h0};
  wire [7:0]         _maskSplit_vlBoundaryCorrection_T_27 = _maskSplit_vlBoundaryCorrection_T_24 | {_maskSplit_vlBoundaryCorrection_T_24[5:0], 2'h0};
  wire [7:0]         maskSplit_vlBoundaryCorrection_1 =
    ~({8{maskSplit_vlMisAlign_1 & maskSplit_isVlBoundary_1}} & (_maskSplit_vlBoundaryCorrection_T_27 | {_maskSplit_vlBoundaryCorrection_T_27[3:0], 4'h0})) & {8{maskSplit_validExecuteGroup_1}};
  wire [1023:0][7:0] _GEN_145 =
    {{maskSplit_maskSelect_hi_1[4095:4088]},
     {maskSplit_maskSelect_hi_1[4087:4080]},
     {maskSplit_maskSelect_hi_1[4079:4072]},
     {maskSplit_maskSelect_hi_1[4071:4064]},
     {maskSplit_maskSelect_hi_1[4063:4056]},
     {maskSplit_maskSelect_hi_1[4055:4048]},
     {maskSplit_maskSelect_hi_1[4047:4040]},
     {maskSplit_maskSelect_hi_1[4039:4032]},
     {maskSplit_maskSelect_hi_1[4031:4024]},
     {maskSplit_maskSelect_hi_1[4023:4016]},
     {maskSplit_maskSelect_hi_1[4015:4008]},
     {maskSplit_maskSelect_hi_1[4007:4000]},
     {maskSplit_maskSelect_hi_1[3999:3992]},
     {maskSplit_maskSelect_hi_1[3991:3984]},
     {maskSplit_maskSelect_hi_1[3983:3976]},
     {maskSplit_maskSelect_hi_1[3975:3968]},
     {maskSplit_maskSelect_hi_1[3967:3960]},
     {maskSplit_maskSelect_hi_1[3959:3952]},
     {maskSplit_maskSelect_hi_1[3951:3944]},
     {maskSplit_maskSelect_hi_1[3943:3936]},
     {maskSplit_maskSelect_hi_1[3935:3928]},
     {maskSplit_maskSelect_hi_1[3927:3920]},
     {maskSplit_maskSelect_hi_1[3919:3912]},
     {maskSplit_maskSelect_hi_1[3911:3904]},
     {maskSplit_maskSelect_hi_1[3903:3896]},
     {maskSplit_maskSelect_hi_1[3895:3888]},
     {maskSplit_maskSelect_hi_1[3887:3880]},
     {maskSplit_maskSelect_hi_1[3879:3872]},
     {maskSplit_maskSelect_hi_1[3871:3864]},
     {maskSplit_maskSelect_hi_1[3863:3856]},
     {maskSplit_maskSelect_hi_1[3855:3848]},
     {maskSplit_maskSelect_hi_1[3847:3840]},
     {maskSplit_maskSelect_hi_1[3839:3832]},
     {maskSplit_maskSelect_hi_1[3831:3824]},
     {maskSplit_maskSelect_hi_1[3823:3816]},
     {maskSplit_maskSelect_hi_1[3815:3808]},
     {maskSplit_maskSelect_hi_1[3807:3800]},
     {maskSplit_maskSelect_hi_1[3799:3792]},
     {maskSplit_maskSelect_hi_1[3791:3784]},
     {maskSplit_maskSelect_hi_1[3783:3776]},
     {maskSplit_maskSelect_hi_1[3775:3768]},
     {maskSplit_maskSelect_hi_1[3767:3760]},
     {maskSplit_maskSelect_hi_1[3759:3752]},
     {maskSplit_maskSelect_hi_1[3751:3744]},
     {maskSplit_maskSelect_hi_1[3743:3736]},
     {maskSplit_maskSelect_hi_1[3735:3728]},
     {maskSplit_maskSelect_hi_1[3727:3720]},
     {maskSplit_maskSelect_hi_1[3719:3712]},
     {maskSplit_maskSelect_hi_1[3711:3704]},
     {maskSplit_maskSelect_hi_1[3703:3696]},
     {maskSplit_maskSelect_hi_1[3695:3688]},
     {maskSplit_maskSelect_hi_1[3687:3680]},
     {maskSplit_maskSelect_hi_1[3679:3672]},
     {maskSplit_maskSelect_hi_1[3671:3664]},
     {maskSplit_maskSelect_hi_1[3663:3656]},
     {maskSplit_maskSelect_hi_1[3655:3648]},
     {maskSplit_maskSelect_hi_1[3647:3640]},
     {maskSplit_maskSelect_hi_1[3639:3632]},
     {maskSplit_maskSelect_hi_1[3631:3624]},
     {maskSplit_maskSelect_hi_1[3623:3616]},
     {maskSplit_maskSelect_hi_1[3615:3608]},
     {maskSplit_maskSelect_hi_1[3607:3600]},
     {maskSplit_maskSelect_hi_1[3599:3592]},
     {maskSplit_maskSelect_hi_1[3591:3584]},
     {maskSplit_maskSelect_hi_1[3583:3576]},
     {maskSplit_maskSelect_hi_1[3575:3568]},
     {maskSplit_maskSelect_hi_1[3567:3560]},
     {maskSplit_maskSelect_hi_1[3559:3552]},
     {maskSplit_maskSelect_hi_1[3551:3544]},
     {maskSplit_maskSelect_hi_1[3543:3536]},
     {maskSplit_maskSelect_hi_1[3535:3528]},
     {maskSplit_maskSelect_hi_1[3527:3520]},
     {maskSplit_maskSelect_hi_1[3519:3512]},
     {maskSplit_maskSelect_hi_1[3511:3504]},
     {maskSplit_maskSelect_hi_1[3503:3496]},
     {maskSplit_maskSelect_hi_1[3495:3488]},
     {maskSplit_maskSelect_hi_1[3487:3480]},
     {maskSplit_maskSelect_hi_1[3479:3472]},
     {maskSplit_maskSelect_hi_1[3471:3464]},
     {maskSplit_maskSelect_hi_1[3463:3456]},
     {maskSplit_maskSelect_hi_1[3455:3448]},
     {maskSplit_maskSelect_hi_1[3447:3440]},
     {maskSplit_maskSelect_hi_1[3439:3432]},
     {maskSplit_maskSelect_hi_1[3431:3424]},
     {maskSplit_maskSelect_hi_1[3423:3416]},
     {maskSplit_maskSelect_hi_1[3415:3408]},
     {maskSplit_maskSelect_hi_1[3407:3400]},
     {maskSplit_maskSelect_hi_1[3399:3392]},
     {maskSplit_maskSelect_hi_1[3391:3384]},
     {maskSplit_maskSelect_hi_1[3383:3376]},
     {maskSplit_maskSelect_hi_1[3375:3368]},
     {maskSplit_maskSelect_hi_1[3367:3360]},
     {maskSplit_maskSelect_hi_1[3359:3352]},
     {maskSplit_maskSelect_hi_1[3351:3344]},
     {maskSplit_maskSelect_hi_1[3343:3336]},
     {maskSplit_maskSelect_hi_1[3335:3328]},
     {maskSplit_maskSelect_hi_1[3327:3320]},
     {maskSplit_maskSelect_hi_1[3319:3312]},
     {maskSplit_maskSelect_hi_1[3311:3304]},
     {maskSplit_maskSelect_hi_1[3303:3296]},
     {maskSplit_maskSelect_hi_1[3295:3288]},
     {maskSplit_maskSelect_hi_1[3287:3280]},
     {maskSplit_maskSelect_hi_1[3279:3272]},
     {maskSplit_maskSelect_hi_1[3271:3264]},
     {maskSplit_maskSelect_hi_1[3263:3256]},
     {maskSplit_maskSelect_hi_1[3255:3248]},
     {maskSplit_maskSelect_hi_1[3247:3240]},
     {maskSplit_maskSelect_hi_1[3239:3232]},
     {maskSplit_maskSelect_hi_1[3231:3224]},
     {maskSplit_maskSelect_hi_1[3223:3216]},
     {maskSplit_maskSelect_hi_1[3215:3208]},
     {maskSplit_maskSelect_hi_1[3207:3200]},
     {maskSplit_maskSelect_hi_1[3199:3192]},
     {maskSplit_maskSelect_hi_1[3191:3184]},
     {maskSplit_maskSelect_hi_1[3183:3176]},
     {maskSplit_maskSelect_hi_1[3175:3168]},
     {maskSplit_maskSelect_hi_1[3167:3160]},
     {maskSplit_maskSelect_hi_1[3159:3152]},
     {maskSplit_maskSelect_hi_1[3151:3144]},
     {maskSplit_maskSelect_hi_1[3143:3136]},
     {maskSplit_maskSelect_hi_1[3135:3128]},
     {maskSplit_maskSelect_hi_1[3127:3120]},
     {maskSplit_maskSelect_hi_1[3119:3112]},
     {maskSplit_maskSelect_hi_1[3111:3104]},
     {maskSplit_maskSelect_hi_1[3103:3096]},
     {maskSplit_maskSelect_hi_1[3095:3088]},
     {maskSplit_maskSelect_hi_1[3087:3080]},
     {maskSplit_maskSelect_hi_1[3079:3072]},
     {maskSplit_maskSelect_hi_1[3071:3064]},
     {maskSplit_maskSelect_hi_1[3063:3056]},
     {maskSplit_maskSelect_hi_1[3055:3048]},
     {maskSplit_maskSelect_hi_1[3047:3040]},
     {maskSplit_maskSelect_hi_1[3039:3032]},
     {maskSplit_maskSelect_hi_1[3031:3024]},
     {maskSplit_maskSelect_hi_1[3023:3016]},
     {maskSplit_maskSelect_hi_1[3015:3008]},
     {maskSplit_maskSelect_hi_1[3007:3000]},
     {maskSplit_maskSelect_hi_1[2999:2992]},
     {maskSplit_maskSelect_hi_1[2991:2984]},
     {maskSplit_maskSelect_hi_1[2983:2976]},
     {maskSplit_maskSelect_hi_1[2975:2968]},
     {maskSplit_maskSelect_hi_1[2967:2960]},
     {maskSplit_maskSelect_hi_1[2959:2952]},
     {maskSplit_maskSelect_hi_1[2951:2944]},
     {maskSplit_maskSelect_hi_1[2943:2936]},
     {maskSplit_maskSelect_hi_1[2935:2928]},
     {maskSplit_maskSelect_hi_1[2927:2920]},
     {maskSplit_maskSelect_hi_1[2919:2912]},
     {maskSplit_maskSelect_hi_1[2911:2904]},
     {maskSplit_maskSelect_hi_1[2903:2896]},
     {maskSplit_maskSelect_hi_1[2895:2888]},
     {maskSplit_maskSelect_hi_1[2887:2880]},
     {maskSplit_maskSelect_hi_1[2879:2872]},
     {maskSplit_maskSelect_hi_1[2871:2864]},
     {maskSplit_maskSelect_hi_1[2863:2856]},
     {maskSplit_maskSelect_hi_1[2855:2848]},
     {maskSplit_maskSelect_hi_1[2847:2840]},
     {maskSplit_maskSelect_hi_1[2839:2832]},
     {maskSplit_maskSelect_hi_1[2831:2824]},
     {maskSplit_maskSelect_hi_1[2823:2816]},
     {maskSplit_maskSelect_hi_1[2815:2808]},
     {maskSplit_maskSelect_hi_1[2807:2800]},
     {maskSplit_maskSelect_hi_1[2799:2792]},
     {maskSplit_maskSelect_hi_1[2791:2784]},
     {maskSplit_maskSelect_hi_1[2783:2776]},
     {maskSplit_maskSelect_hi_1[2775:2768]},
     {maskSplit_maskSelect_hi_1[2767:2760]},
     {maskSplit_maskSelect_hi_1[2759:2752]},
     {maskSplit_maskSelect_hi_1[2751:2744]},
     {maskSplit_maskSelect_hi_1[2743:2736]},
     {maskSplit_maskSelect_hi_1[2735:2728]},
     {maskSplit_maskSelect_hi_1[2727:2720]},
     {maskSplit_maskSelect_hi_1[2719:2712]},
     {maskSplit_maskSelect_hi_1[2711:2704]},
     {maskSplit_maskSelect_hi_1[2703:2696]},
     {maskSplit_maskSelect_hi_1[2695:2688]},
     {maskSplit_maskSelect_hi_1[2687:2680]},
     {maskSplit_maskSelect_hi_1[2679:2672]},
     {maskSplit_maskSelect_hi_1[2671:2664]},
     {maskSplit_maskSelect_hi_1[2663:2656]},
     {maskSplit_maskSelect_hi_1[2655:2648]},
     {maskSplit_maskSelect_hi_1[2647:2640]},
     {maskSplit_maskSelect_hi_1[2639:2632]},
     {maskSplit_maskSelect_hi_1[2631:2624]},
     {maskSplit_maskSelect_hi_1[2623:2616]},
     {maskSplit_maskSelect_hi_1[2615:2608]},
     {maskSplit_maskSelect_hi_1[2607:2600]},
     {maskSplit_maskSelect_hi_1[2599:2592]},
     {maskSplit_maskSelect_hi_1[2591:2584]},
     {maskSplit_maskSelect_hi_1[2583:2576]},
     {maskSplit_maskSelect_hi_1[2575:2568]},
     {maskSplit_maskSelect_hi_1[2567:2560]},
     {maskSplit_maskSelect_hi_1[2559:2552]},
     {maskSplit_maskSelect_hi_1[2551:2544]},
     {maskSplit_maskSelect_hi_1[2543:2536]},
     {maskSplit_maskSelect_hi_1[2535:2528]},
     {maskSplit_maskSelect_hi_1[2527:2520]},
     {maskSplit_maskSelect_hi_1[2519:2512]},
     {maskSplit_maskSelect_hi_1[2511:2504]},
     {maskSplit_maskSelect_hi_1[2503:2496]},
     {maskSplit_maskSelect_hi_1[2495:2488]},
     {maskSplit_maskSelect_hi_1[2487:2480]},
     {maskSplit_maskSelect_hi_1[2479:2472]},
     {maskSplit_maskSelect_hi_1[2471:2464]},
     {maskSplit_maskSelect_hi_1[2463:2456]},
     {maskSplit_maskSelect_hi_1[2455:2448]},
     {maskSplit_maskSelect_hi_1[2447:2440]},
     {maskSplit_maskSelect_hi_1[2439:2432]},
     {maskSplit_maskSelect_hi_1[2431:2424]},
     {maskSplit_maskSelect_hi_1[2423:2416]},
     {maskSplit_maskSelect_hi_1[2415:2408]},
     {maskSplit_maskSelect_hi_1[2407:2400]},
     {maskSplit_maskSelect_hi_1[2399:2392]},
     {maskSplit_maskSelect_hi_1[2391:2384]},
     {maskSplit_maskSelect_hi_1[2383:2376]},
     {maskSplit_maskSelect_hi_1[2375:2368]},
     {maskSplit_maskSelect_hi_1[2367:2360]},
     {maskSplit_maskSelect_hi_1[2359:2352]},
     {maskSplit_maskSelect_hi_1[2351:2344]},
     {maskSplit_maskSelect_hi_1[2343:2336]},
     {maskSplit_maskSelect_hi_1[2335:2328]},
     {maskSplit_maskSelect_hi_1[2327:2320]},
     {maskSplit_maskSelect_hi_1[2319:2312]},
     {maskSplit_maskSelect_hi_1[2311:2304]},
     {maskSplit_maskSelect_hi_1[2303:2296]},
     {maskSplit_maskSelect_hi_1[2295:2288]},
     {maskSplit_maskSelect_hi_1[2287:2280]},
     {maskSplit_maskSelect_hi_1[2279:2272]},
     {maskSplit_maskSelect_hi_1[2271:2264]},
     {maskSplit_maskSelect_hi_1[2263:2256]},
     {maskSplit_maskSelect_hi_1[2255:2248]},
     {maskSplit_maskSelect_hi_1[2247:2240]},
     {maskSplit_maskSelect_hi_1[2239:2232]},
     {maskSplit_maskSelect_hi_1[2231:2224]},
     {maskSplit_maskSelect_hi_1[2223:2216]},
     {maskSplit_maskSelect_hi_1[2215:2208]},
     {maskSplit_maskSelect_hi_1[2207:2200]},
     {maskSplit_maskSelect_hi_1[2199:2192]},
     {maskSplit_maskSelect_hi_1[2191:2184]},
     {maskSplit_maskSelect_hi_1[2183:2176]},
     {maskSplit_maskSelect_hi_1[2175:2168]},
     {maskSplit_maskSelect_hi_1[2167:2160]},
     {maskSplit_maskSelect_hi_1[2159:2152]},
     {maskSplit_maskSelect_hi_1[2151:2144]},
     {maskSplit_maskSelect_hi_1[2143:2136]},
     {maskSplit_maskSelect_hi_1[2135:2128]},
     {maskSplit_maskSelect_hi_1[2127:2120]},
     {maskSplit_maskSelect_hi_1[2119:2112]},
     {maskSplit_maskSelect_hi_1[2111:2104]},
     {maskSplit_maskSelect_hi_1[2103:2096]},
     {maskSplit_maskSelect_hi_1[2095:2088]},
     {maskSplit_maskSelect_hi_1[2087:2080]},
     {maskSplit_maskSelect_hi_1[2079:2072]},
     {maskSplit_maskSelect_hi_1[2071:2064]},
     {maskSplit_maskSelect_hi_1[2063:2056]},
     {maskSplit_maskSelect_hi_1[2055:2048]},
     {maskSplit_maskSelect_hi_1[2047:2040]},
     {maskSplit_maskSelect_hi_1[2039:2032]},
     {maskSplit_maskSelect_hi_1[2031:2024]},
     {maskSplit_maskSelect_hi_1[2023:2016]},
     {maskSplit_maskSelect_hi_1[2015:2008]},
     {maskSplit_maskSelect_hi_1[2007:2000]},
     {maskSplit_maskSelect_hi_1[1999:1992]},
     {maskSplit_maskSelect_hi_1[1991:1984]},
     {maskSplit_maskSelect_hi_1[1983:1976]},
     {maskSplit_maskSelect_hi_1[1975:1968]},
     {maskSplit_maskSelect_hi_1[1967:1960]},
     {maskSplit_maskSelect_hi_1[1959:1952]},
     {maskSplit_maskSelect_hi_1[1951:1944]},
     {maskSplit_maskSelect_hi_1[1943:1936]},
     {maskSplit_maskSelect_hi_1[1935:1928]},
     {maskSplit_maskSelect_hi_1[1927:1920]},
     {maskSplit_maskSelect_hi_1[1919:1912]},
     {maskSplit_maskSelect_hi_1[1911:1904]},
     {maskSplit_maskSelect_hi_1[1903:1896]},
     {maskSplit_maskSelect_hi_1[1895:1888]},
     {maskSplit_maskSelect_hi_1[1887:1880]},
     {maskSplit_maskSelect_hi_1[1879:1872]},
     {maskSplit_maskSelect_hi_1[1871:1864]},
     {maskSplit_maskSelect_hi_1[1863:1856]},
     {maskSplit_maskSelect_hi_1[1855:1848]},
     {maskSplit_maskSelect_hi_1[1847:1840]},
     {maskSplit_maskSelect_hi_1[1839:1832]},
     {maskSplit_maskSelect_hi_1[1831:1824]},
     {maskSplit_maskSelect_hi_1[1823:1816]},
     {maskSplit_maskSelect_hi_1[1815:1808]},
     {maskSplit_maskSelect_hi_1[1807:1800]},
     {maskSplit_maskSelect_hi_1[1799:1792]},
     {maskSplit_maskSelect_hi_1[1791:1784]},
     {maskSplit_maskSelect_hi_1[1783:1776]},
     {maskSplit_maskSelect_hi_1[1775:1768]},
     {maskSplit_maskSelect_hi_1[1767:1760]},
     {maskSplit_maskSelect_hi_1[1759:1752]},
     {maskSplit_maskSelect_hi_1[1751:1744]},
     {maskSplit_maskSelect_hi_1[1743:1736]},
     {maskSplit_maskSelect_hi_1[1735:1728]},
     {maskSplit_maskSelect_hi_1[1727:1720]},
     {maskSplit_maskSelect_hi_1[1719:1712]},
     {maskSplit_maskSelect_hi_1[1711:1704]},
     {maskSplit_maskSelect_hi_1[1703:1696]},
     {maskSplit_maskSelect_hi_1[1695:1688]},
     {maskSplit_maskSelect_hi_1[1687:1680]},
     {maskSplit_maskSelect_hi_1[1679:1672]},
     {maskSplit_maskSelect_hi_1[1671:1664]},
     {maskSplit_maskSelect_hi_1[1663:1656]},
     {maskSplit_maskSelect_hi_1[1655:1648]},
     {maskSplit_maskSelect_hi_1[1647:1640]},
     {maskSplit_maskSelect_hi_1[1639:1632]},
     {maskSplit_maskSelect_hi_1[1631:1624]},
     {maskSplit_maskSelect_hi_1[1623:1616]},
     {maskSplit_maskSelect_hi_1[1615:1608]},
     {maskSplit_maskSelect_hi_1[1607:1600]},
     {maskSplit_maskSelect_hi_1[1599:1592]},
     {maskSplit_maskSelect_hi_1[1591:1584]},
     {maskSplit_maskSelect_hi_1[1583:1576]},
     {maskSplit_maskSelect_hi_1[1575:1568]},
     {maskSplit_maskSelect_hi_1[1567:1560]},
     {maskSplit_maskSelect_hi_1[1559:1552]},
     {maskSplit_maskSelect_hi_1[1551:1544]},
     {maskSplit_maskSelect_hi_1[1543:1536]},
     {maskSplit_maskSelect_hi_1[1535:1528]},
     {maskSplit_maskSelect_hi_1[1527:1520]},
     {maskSplit_maskSelect_hi_1[1519:1512]},
     {maskSplit_maskSelect_hi_1[1511:1504]},
     {maskSplit_maskSelect_hi_1[1503:1496]},
     {maskSplit_maskSelect_hi_1[1495:1488]},
     {maskSplit_maskSelect_hi_1[1487:1480]},
     {maskSplit_maskSelect_hi_1[1479:1472]},
     {maskSplit_maskSelect_hi_1[1471:1464]},
     {maskSplit_maskSelect_hi_1[1463:1456]},
     {maskSplit_maskSelect_hi_1[1455:1448]},
     {maskSplit_maskSelect_hi_1[1447:1440]},
     {maskSplit_maskSelect_hi_1[1439:1432]},
     {maskSplit_maskSelect_hi_1[1431:1424]},
     {maskSplit_maskSelect_hi_1[1423:1416]},
     {maskSplit_maskSelect_hi_1[1415:1408]},
     {maskSplit_maskSelect_hi_1[1407:1400]},
     {maskSplit_maskSelect_hi_1[1399:1392]},
     {maskSplit_maskSelect_hi_1[1391:1384]},
     {maskSplit_maskSelect_hi_1[1383:1376]},
     {maskSplit_maskSelect_hi_1[1375:1368]},
     {maskSplit_maskSelect_hi_1[1367:1360]},
     {maskSplit_maskSelect_hi_1[1359:1352]},
     {maskSplit_maskSelect_hi_1[1351:1344]},
     {maskSplit_maskSelect_hi_1[1343:1336]},
     {maskSplit_maskSelect_hi_1[1335:1328]},
     {maskSplit_maskSelect_hi_1[1327:1320]},
     {maskSplit_maskSelect_hi_1[1319:1312]},
     {maskSplit_maskSelect_hi_1[1311:1304]},
     {maskSplit_maskSelect_hi_1[1303:1296]},
     {maskSplit_maskSelect_hi_1[1295:1288]},
     {maskSplit_maskSelect_hi_1[1287:1280]},
     {maskSplit_maskSelect_hi_1[1279:1272]},
     {maskSplit_maskSelect_hi_1[1271:1264]},
     {maskSplit_maskSelect_hi_1[1263:1256]},
     {maskSplit_maskSelect_hi_1[1255:1248]},
     {maskSplit_maskSelect_hi_1[1247:1240]},
     {maskSplit_maskSelect_hi_1[1239:1232]},
     {maskSplit_maskSelect_hi_1[1231:1224]},
     {maskSplit_maskSelect_hi_1[1223:1216]},
     {maskSplit_maskSelect_hi_1[1215:1208]},
     {maskSplit_maskSelect_hi_1[1207:1200]},
     {maskSplit_maskSelect_hi_1[1199:1192]},
     {maskSplit_maskSelect_hi_1[1191:1184]},
     {maskSplit_maskSelect_hi_1[1183:1176]},
     {maskSplit_maskSelect_hi_1[1175:1168]},
     {maskSplit_maskSelect_hi_1[1167:1160]},
     {maskSplit_maskSelect_hi_1[1159:1152]},
     {maskSplit_maskSelect_hi_1[1151:1144]},
     {maskSplit_maskSelect_hi_1[1143:1136]},
     {maskSplit_maskSelect_hi_1[1135:1128]},
     {maskSplit_maskSelect_hi_1[1127:1120]},
     {maskSplit_maskSelect_hi_1[1119:1112]},
     {maskSplit_maskSelect_hi_1[1111:1104]},
     {maskSplit_maskSelect_hi_1[1103:1096]},
     {maskSplit_maskSelect_hi_1[1095:1088]},
     {maskSplit_maskSelect_hi_1[1087:1080]},
     {maskSplit_maskSelect_hi_1[1079:1072]},
     {maskSplit_maskSelect_hi_1[1071:1064]},
     {maskSplit_maskSelect_hi_1[1063:1056]},
     {maskSplit_maskSelect_hi_1[1055:1048]},
     {maskSplit_maskSelect_hi_1[1047:1040]},
     {maskSplit_maskSelect_hi_1[1039:1032]},
     {maskSplit_maskSelect_hi_1[1031:1024]},
     {maskSplit_maskSelect_hi_1[1023:1016]},
     {maskSplit_maskSelect_hi_1[1015:1008]},
     {maskSplit_maskSelect_hi_1[1007:1000]},
     {maskSplit_maskSelect_hi_1[999:992]},
     {maskSplit_maskSelect_hi_1[991:984]},
     {maskSplit_maskSelect_hi_1[983:976]},
     {maskSplit_maskSelect_hi_1[975:968]},
     {maskSplit_maskSelect_hi_1[967:960]},
     {maskSplit_maskSelect_hi_1[959:952]},
     {maskSplit_maskSelect_hi_1[951:944]},
     {maskSplit_maskSelect_hi_1[943:936]},
     {maskSplit_maskSelect_hi_1[935:928]},
     {maskSplit_maskSelect_hi_1[927:920]},
     {maskSplit_maskSelect_hi_1[919:912]},
     {maskSplit_maskSelect_hi_1[911:904]},
     {maskSplit_maskSelect_hi_1[903:896]},
     {maskSplit_maskSelect_hi_1[895:888]},
     {maskSplit_maskSelect_hi_1[887:880]},
     {maskSplit_maskSelect_hi_1[879:872]},
     {maskSplit_maskSelect_hi_1[871:864]},
     {maskSplit_maskSelect_hi_1[863:856]},
     {maskSplit_maskSelect_hi_1[855:848]},
     {maskSplit_maskSelect_hi_1[847:840]},
     {maskSplit_maskSelect_hi_1[839:832]},
     {maskSplit_maskSelect_hi_1[831:824]},
     {maskSplit_maskSelect_hi_1[823:816]},
     {maskSplit_maskSelect_hi_1[815:808]},
     {maskSplit_maskSelect_hi_1[807:800]},
     {maskSplit_maskSelect_hi_1[799:792]},
     {maskSplit_maskSelect_hi_1[791:784]},
     {maskSplit_maskSelect_hi_1[783:776]},
     {maskSplit_maskSelect_hi_1[775:768]},
     {maskSplit_maskSelect_hi_1[767:760]},
     {maskSplit_maskSelect_hi_1[759:752]},
     {maskSplit_maskSelect_hi_1[751:744]},
     {maskSplit_maskSelect_hi_1[743:736]},
     {maskSplit_maskSelect_hi_1[735:728]},
     {maskSplit_maskSelect_hi_1[727:720]},
     {maskSplit_maskSelect_hi_1[719:712]},
     {maskSplit_maskSelect_hi_1[711:704]},
     {maskSplit_maskSelect_hi_1[703:696]},
     {maskSplit_maskSelect_hi_1[695:688]},
     {maskSplit_maskSelect_hi_1[687:680]},
     {maskSplit_maskSelect_hi_1[679:672]},
     {maskSplit_maskSelect_hi_1[671:664]},
     {maskSplit_maskSelect_hi_1[663:656]},
     {maskSplit_maskSelect_hi_1[655:648]},
     {maskSplit_maskSelect_hi_1[647:640]},
     {maskSplit_maskSelect_hi_1[639:632]},
     {maskSplit_maskSelect_hi_1[631:624]},
     {maskSplit_maskSelect_hi_1[623:616]},
     {maskSplit_maskSelect_hi_1[615:608]},
     {maskSplit_maskSelect_hi_1[607:600]},
     {maskSplit_maskSelect_hi_1[599:592]},
     {maskSplit_maskSelect_hi_1[591:584]},
     {maskSplit_maskSelect_hi_1[583:576]},
     {maskSplit_maskSelect_hi_1[575:568]},
     {maskSplit_maskSelect_hi_1[567:560]},
     {maskSplit_maskSelect_hi_1[559:552]},
     {maskSplit_maskSelect_hi_1[551:544]},
     {maskSplit_maskSelect_hi_1[543:536]},
     {maskSplit_maskSelect_hi_1[535:528]},
     {maskSplit_maskSelect_hi_1[527:520]},
     {maskSplit_maskSelect_hi_1[519:512]},
     {maskSplit_maskSelect_hi_1[511:504]},
     {maskSplit_maskSelect_hi_1[503:496]},
     {maskSplit_maskSelect_hi_1[495:488]},
     {maskSplit_maskSelect_hi_1[487:480]},
     {maskSplit_maskSelect_hi_1[479:472]},
     {maskSplit_maskSelect_hi_1[471:464]},
     {maskSplit_maskSelect_hi_1[463:456]},
     {maskSplit_maskSelect_hi_1[455:448]},
     {maskSplit_maskSelect_hi_1[447:440]},
     {maskSplit_maskSelect_hi_1[439:432]},
     {maskSplit_maskSelect_hi_1[431:424]},
     {maskSplit_maskSelect_hi_1[423:416]},
     {maskSplit_maskSelect_hi_1[415:408]},
     {maskSplit_maskSelect_hi_1[407:400]},
     {maskSplit_maskSelect_hi_1[399:392]},
     {maskSplit_maskSelect_hi_1[391:384]},
     {maskSplit_maskSelect_hi_1[383:376]},
     {maskSplit_maskSelect_hi_1[375:368]},
     {maskSplit_maskSelect_hi_1[367:360]},
     {maskSplit_maskSelect_hi_1[359:352]},
     {maskSplit_maskSelect_hi_1[351:344]},
     {maskSplit_maskSelect_hi_1[343:336]},
     {maskSplit_maskSelect_hi_1[335:328]},
     {maskSplit_maskSelect_hi_1[327:320]},
     {maskSplit_maskSelect_hi_1[319:312]},
     {maskSplit_maskSelect_hi_1[311:304]},
     {maskSplit_maskSelect_hi_1[303:296]},
     {maskSplit_maskSelect_hi_1[295:288]},
     {maskSplit_maskSelect_hi_1[287:280]},
     {maskSplit_maskSelect_hi_1[279:272]},
     {maskSplit_maskSelect_hi_1[271:264]},
     {maskSplit_maskSelect_hi_1[263:256]},
     {maskSplit_maskSelect_hi_1[255:248]},
     {maskSplit_maskSelect_hi_1[247:240]},
     {maskSplit_maskSelect_hi_1[239:232]},
     {maskSplit_maskSelect_hi_1[231:224]},
     {maskSplit_maskSelect_hi_1[223:216]},
     {maskSplit_maskSelect_hi_1[215:208]},
     {maskSplit_maskSelect_hi_1[207:200]},
     {maskSplit_maskSelect_hi_1[199:192]},
     {maskSplit_maskSelect_hi_1[191:184]},
     {maskSplit_maskSelect_hi_1[183:176]},
     {maskSplit_maskSelect_hi_1[175:168]},
     {maskSplit_maskSelect_hi_1[167:160]},
     {maskSplit_maskSelect_hi_1[159:152]},
     {maskSplit_maskSelect_hi_1[151:144]},
     {maskSplit_maskSelect_hi_1[143:136]},
     {maskSplit_maskSelect_hi_1[135:128]},
     {maskSplit_maskSelect_hi_1[127:120]},
     {maskSplit_maskSelect_hi_1[119:112]},
     {maskSplit_maskSelect_hi_1[111:104]},
     {maskSplit_maskSelect_hi_1[103:96]},
     {maskSplit_maskSelect_hi_1[95:88]},
     {maskSplit_maskSelect_hi_1[87:80]},
     {maskSplit_maskSelect_hi_1[79:72]},
     {maskSplit_maskSelect_hi_1[71:64]},
     {maskSplit_maskSelect_hi_1[63:56]},
     {maskSplit_maskSelect_hi_1[55:48]},
     {maskSplit_maskSelect_hi_1[47:40]},
     {maskSplit_maskSelect_hi_1[39:32]},
     {maskSplit_maskSelect_hi_1[31:24]},
     {maskSplit_maskSelect_hi_1[23:16]},
     {maskSplit_maskSelect_hi_1[15:8]},
     {maskSplit_maskSelect_hi_1[7:0]},
     {maskSplit_maskSelect_lo_1[4095:4088]},
     {maskSplit_maskSelect_lo_1[4087:4080]},
     {maskSplit_maskSelect_lo_1[4079:4072]},
     {maskSplit_maskSelect_lo_1[4071:4064]},
     {maskSplit_maskSelect_lo_1[4063:4056]},
     {maskSplit_maskSelect_lo_1[4055:4048]},
     {maskSplit_maskSelect_lo_1[4047:4040]},
     {maskSplit_maskSelect_lo_1[4039:4032]},
     {maskSplit_maskSelect_lo_1[4031:4024]},
     {maskSplit_maskSelect_lo_1[4023:4016]},
     {maskSplit_maskSelect_lo_1[4015:4008]},
     {maskSplit_maskSelect_lo_1[4007:4000]},
     {maskSplit_maskSelect_lo_1[3999:3992]},
     {maskSplit_maskSelect_lo_1[3991:3984]},
     {maskSplit_maskSelect_lo_1[3983:3976]},
     {maskSplit_maskSelect_lo_1[3975:3968]},
     {maskSplit_maskSelect_lo_1[3967:3960]},
     {maskSplit_maskSelect_lo_1[3959:3952]},
     {maskSplit_maskSelect_lo_1[3951:3944]},
     {maskSplit_maskSelect_lo_1[3943:3936]},
     {maskSplit_maskSelect_lo_1[3935:3928]},
     {maskSplit_maskSelect_lo_1[3927:3920]},
     {maskSplit_maskSelect_lo_1[3919:3912]},
     {maskSplit_maskSelect_lo_1[3911:3904]},
     {maskSplit_maskSelect_lo_1[3903:3896]},
     {maskSplit_maskSelect_lo_1[3895:3888]},
     {maskSplit_maskSelect_lo_1[3887:3880]},
     {maskSplit_maskSelect_lo_1[3879:3872]},
     {maskSplit_maskSelect_lo_1[3871:3864]},
     {maskSplit_maskSelect_lo_1[3863:3856]},
     {maskSplit_maskSelect_lo_1[3855:3848]},
     {maskSplit_maskSelect_lo_1[3847:3840]},
     {maskSplit_maskSelect_lo_1[3839:3832]},
     {maskSplit_maskSelect_lo_1[3831:3824]},
     {maskSplit_maskSelect_lo_1[3823:3816]},
     {maskSplit_maskSelect_lo_1[3815:3808]},
     {maskSplit_maskSelect_lo_1[3807:3800]},
     {maskSplit_maskSelect_lo_1[3799:3792]},
     {maskSplit_maskSelect_lo_1[3791:3784]},
     {maskSplit_maskSelect_lo_1[3783:3776]},
     {maskSplit_maskSelect_lo_1[3775:3768]},
     {maskSplit_maskSelect_lo_1[3767:3760]},
     {maskSplit_maskSelect_lo_1[3759:3752]},
     {maskSplit_maskSelect_lo_1[3751:3744]},
     {maskSplit_maskSelect_lo_1[3743:3736]},
     {maskSplit_maskSelect_lo_1[3735:3728]},
     {maskSplit_maskSelect_lo_1[3727:3720]},
     {maskSplit_maskSelect_lo_1[3719:3712]},
     {maskSplit_maskSelect_lo_1[3711:3704]},
     {maskSplit_maskSelect_lo_1[3703:3696]},
     {maskSplit_maskSelect_lo_1[3695:3688]},
     {maskSplit_maskSelect_lo_1[3687:3680]},
     {maskSplit_maskSelect_lo_1[3679:3672]},
     {maskSplit_maskSelect_lo_1[3671:3664]},
     {maskSplit_maskSelect_lo_1[3663:3656]},
     {maskSplit_maskSelect_lo_1[3655:3648]},
     {maskSplit_maskSelect_lo_1[3647:3640]},
     {maskSplit_maskSelect_lo_1[3639:3632]},
     {maskSplit_maskSelect_lo_1[3631:3624]},
     {maskSplit_maskSelect_lo_1[3623:3616]},
     {maskSplit_maskSelect_lo_1[3615:3608]},
     {maskSplit_maskSelect_lo_1[3607:3600]},
     {maskSplit_maskSelect_lo_1[3599:3592]},
     {maskSplit_maskSelect_lo_1[3591:3584]},
     {maskSplit_maskSelect_lo_1[3583:3576]},
     {maskSplit_maskSelect_lo_1[3575:3568]},
     {maskSplit_maskSelect_lo_1[3567:3560]},
     {maskSplit_maskSelect_lo_1[3559:3552]},
     {maskSplit_maskSelect_lo_1[3551:3544]},
     {maskSplit_maskSelect_lo_1[3543:3536]},
     {maskSplit_maskSelect_lo_1[3535:3528]},
     {maskSplit_maskSelect_lo_1[3527:3520]},
     {maskSplit_maskSelect_lo_1[3519:3512]},
     {maskSplit_maskSelect_lo_1[3511:3504]},
     {maskSplit_maskSelect_lo_1[3503:3496]},
     {maskSplit_maskSelect_lo_1[3495:3488]},
     {maskSplit_maskSelect_lo_1[3487:3480]},
     {maskSplit_maskSelect_lo_1[3479:3472]},
     {maskSplit_maskSelect_lo_1[3471:3464]},
     {maskSplit_maskSelect_lo_1[3463:3456]},
     {maskSplit_maskSelect_lo_1[3455:3448]},
     {maskSplit_maskSelect_lo_1[3447:3440]},
     {maskSplit_maskSelect_lo_1[3439:3432]},
     {maskSplit_maskSelect_lo_1[3431:3424]},
     {maskSplit_maskSelect_lo_1[3423:3416]},
     {maskSplit_maskSelect_lo_1[3415:3408]},
     {maskSplit_maskSelect_lo_1[3407:3400]},
     {maskSplit_maskSelect_lo_1[3399:3392]},
     {maskSplit_maskSelect_lo_1[3391:3384]},
     {maskSplit_maskSelect_lo_1[3383:3376]},
     {maskSplit_maskSelect_lo_1[3375:3368]},
     {maskSplit_maskSelect_lo_1[3367:3360]},
     {maskSplit_maskSelect_lo_1[3359:3352]},
     {maskSplit_maskSelect_lo_1[3351:3344]},
     {maskSplit_maskSelect_lo_1[3343:3336]},
     {maskSplit_maskSelect_lo_1[3335:3328]},
     {maskSplit_maskSelect_lo_1[3327:3320]},
     {maskSplit_maskSelect_lo_1[3319:3312]},
     {maskSplit_maskSelect_lo_1[3311:3304]},
     {maskSplit_maskSelect_lo_1[3303:3296]},
     {maskSplit_maskSelect_lo_1[3295:3288]},
     {maskSplit_maskSelect_lo_1[3287:3280]},
     {maskSplit_maskSelect_lo_1[3279:3272]},
     {maskSplit_maskSelect_lo_1[3271:3264]},
     {maskSplit_maskSelect_lo_1[3263:3256]},
     {maskSplit_maskSelect_lo_1[3255:3248]},
     {maskSplit_maskSelect_lo_1[3247:3240]},
     {maskSplit_maskSelect_lo_1[3239:3232]},
     {maskSplit_maskSelect_lo_1[3231:3224]},
     {maskSplit_maskSelect_lo_1[3223:3216]},
     {maskSplit_maskSelect_lo_1[3215:3208]},
     {maskSplit_maskSelect_lo_1[3207:3200]},
     {maskSplit_maskSelect_lo_1[3199:3192]},
     {maskSplit_maskSelect_lo_1[3191:3184]},
     {maskSplit_maskSelect_lo_1[3183:3176]},
     {maskSplit_maskSelect_lo_1[3175:3168]},
     {maskSplit_maskSelect_lo_1[3167:3160]},
     {maskSplit_maskSelect_lo_1[3159:3152]},
     {maskSplit_maskSelect_lo_1[3151:3144]},
     {maskSplit_maskSelect_lo_1[3143:3136]},
     {maskSplit_maskSelect_lo_1[3135:3128]},
     {maskSplit_maskSelect_lo_1[3127:3120]},
     {maskSplit_maskSelect_lo_1[3119:3112]},
     {maskSplit_maskSelect_lo_1[3111:3104]},
     {maskSplit_maskSelect_lo_1[3103:3096]},
     {maskSplit_maskSelect_lo_1[3095:3088]},
     {maskSplit_maskSelect_lo_1[3087:3080]},
     {maskSplit_maskSelect_lo_1[3079:3072]},
     {maskSplit_maskSelect_lo_1[3071:3064]},
     {maskSplit_maskSelect_lo_1[3063:3056]},
     {maskSplit_maskSelect_lo_1[3055:3048]},
     {maskSplit_maskSelect_lo_1[3047:3040]},
     {maskSplit_maskSelect_lo_1[3039:3032]},
     {maskSplit_maskSelect_lo_1[3031:3024]},
     {maskSplit_maskSelect_lo_1[3023:3016]},
     {maskSplit_maskSelect_lo_1[3015:3008]},
     {maskSplit_maskSelect_lo_1[3007:3000]},
     {maskSplit_maskSelect_lo_1[2999:2992]},
     {maskSplit_maskSelect_lo_1[2991:2984]},
     {maskSplit_maskSelect_lo_1[2983:2976]},
     {maskSplit_maskSelect_lo_1[2975:2968]},
     {maskSplit_maskSelect_lo_1[2967:2960]},
     {maskSplit_maskSelect_lo_1[2959:2952]},
     {maskSplit_maskSelect_lo_1[2951:2944]},
     {maskSplit_maskSelect_lo_1[2943:2936]},
     {maskSplit_maskSelect_lo_1[2935:2928]},
     {maskSplit_maskSelect_lo_1[2927:2920]},
     {maskSplit_maskSelect_lo_1[2919:2912]},
     {maskSplit_maskSelect_lo_1[2911:2904]},
     {maskSplit_maskSelect_lo_1[2903:2896]},
     {maskSplit_maskSelect_lo_1[2895:2888]},
     {maskSplit_maskSelect_lo_1[2887:2880]},
     {maskSplit_maskSelect_lo_1[2879:2872]},
     {maskSplit_maskSelect_lo_1[2871:2864]},
     {maskSplit_maskSelect_lo_1[2863:2856]},
     {maskSplit_maskSelect_lo_1[2855:2848]},
     {maskSplit_maskSelect_lo_1[2847:2840]},
     {maskSplit_maskSelect_lo_1[2839:2832]},
     {maskSplit_maskSelect_lo_1[2831:2824]},
     {maskSplit_maskSelect_lo_1[2823:2816]},
     {maskSplit_maskSelect_lo_1[2815:2808]},
     {maskSplit_maskSelect_lo_1[2807:2800]},
     {maskSplit_maskSelect_lo_1[2799:2792]},
     {maskSplit_maskSelect_lo_1[2791:2784]},
     {maskSplit_maskSelect_lo_1[2783:2776]},
     {maskSplit_maskSelect_lo_1[2775:2768]},
     {maskSplit_maskSelect_lo_1[2767:2760]},
     {maskSplit_maskSelect_lo_1[2759:2752]},
     {maskSplit_maskSelect_lo_1[2751:2744]},
     {maskSplit_maskSelect_lo_1[2743:2736]},
     {maskSplit_maskSelect_lo_1[2735:2728]},
     {maskSplit_maskSelect_lo_1[2727:2720]},
     {maskSplit_maskSelect_lo_1[2719:2712]},
     {maskSplit_maskSelect_lo_1[2711:2704]},
     {maskSplit_maskSelect_lo_1[2703:2696]},
     {maskSplit_maskSelect_lo_1[2695:2688]},
     {maskSplit_maskSelect_lo_1[2687:2680]},
     {maskSplit_maskSelect_lo_1[2679:2672]},
     {maskSplit_maskSelect_lo_1[2671:2664]},
     {maskSplit_maskSelect_lo_1[2663:2656]},
     {maskSplit_maskSelect_lo_1[2655:2648]},
     {maskSplit_maskSelect_lo_1[2647:2640]},
     {maskSplit_maskSelect_lo_1[2639:2632]},
     {maskSplit_maskSelect_lo_1[2631:2624]},
     {maskSplit_maskSelect_lo_1[2623:2616]},
     {maskSplit_maskSelect_lo_1[2615:2608]},
     {maskSplit_maskSelect_lo_1[2607:2600]},
     {maskSplit_maskSelect_lo_1[2599:2592]},
     {maskSplit_maskSelect_lo_1[2591:2584]},
     {maskSplit_maskSelect_lo_1[2583:2576]},
     {maskSplit_maskSelect_lo_1[2575:2568]},
     {maskSplit_maskSelect_lo_1[2567:2560]},
     {maskSplit_maskSelect_lo_1[2559:2552]},
     {maskSplit_maskSelect_lo_1[2551:2544]},
     {maskSplit_maskSelect_lo_1[2543:2536]},
     {maskSplit_maskSelect_lo_1[2535:2528]},
     {maskSplit_maskSelect_lo_1[2527:2520]},
     {maskSplit_maskSelect_lo_1[2519:2512]},
     {maskSplit_maskSelect_lo_1[2511:2504]},
     {maskSplit_maskSelect_lo_1[2503:2496]},
     {maskSplit_maskSelect_lo_1[2495:2488]},
     {maskSplit_maskSelect_lo_1[2487:2480]},
     {maskSplit_maskSelect_lo_1[2479:2472]},
     {maskSplit_maskSelect_lo_1[2471:2464]},
     {maskSplit_maskSelect_lo_1[2463:2456]},
     {maskSplit_maskSelect_lo_1[2455:2448]},
     {maskSplit_maskSelect_lo_1[2447:2440]},
     {maskSplit_maskSelect_lo_1[2439:2432]},
     {maskSplit_maskSelect_lo_1[2431:2424]},
     {maskSplit_maskSelect_lo_1[2423:2416]},
     {maskSplit_maskSelect_lo_1[2415:2408]},
     {maskSplit_maskSelect_lo_1[2407:2400]},
     {maskSplit_maskSelect_lo_1[2399:2392]},
     {maskSplit_maskSelect_lo_1[2391:2384]},
     {maskSplit_maskSelect_lo_1[2383:2376]},
     {maskSplit_maskSelect_lo_1[2375:2368]},
     {maskSplit_maskSelect_lo_1[2367:2360]},
     {maskSplit_maskSelect_lo_1[2359:2352]},
     {maskSplit_maskSelect_lo_1[2351:2344]},
     {maskSplit_maskSelect_lo_1[2343:2336]},
     {maskSplit_maskSelect_lo_1[2335:2328]},
     {maskSplit_maskSelect_lo_1[2327:2320]},
     {maskSplit_maskSelect_lo_1[2319:2312]},
     {maskSplit_maskSelect_lo_1[2311:2304]},
     {maskSplit_maskSelect_lo_1[2303:2296]},
     {maskSplit_maskSelect_lo_1[2295:2288]},
     {maskSplit_maskSelect_lo_1[2287:2280]},
     {maskSplit_maskSelect_lo_1[2279:2272]},
     {maskSplit_maskSelect_lo_1[2271:2264]},
     {maskSplit_maskSelect_lo_1[2263:2256]},
     {maskSplit_maskSelect_lo_1[2255:2248]},
     {maskSplit_maskSelect_lo_1[2247:2240]},
     {maskSplit_maskSelect_lo_1[2239:2232]},
     {maskSplit_maskSelect_lo_1[2231:2224]},
     {maskSplit_maskSelect_lo_1[2223:2216]},
     {maskSplit_maskSelect_lo_1[2215:2208]},
     {maskSplit_maskSelect_lo_1[2207:2200]},
     {maskSplit_maskSelect_lo_1[2199:2192]},
     {maskSplit_maskSelect_lo_1[2191:2184]},
     {maskSplit_maskSelect_lo_1[2183:2176]},
     {maskSplit_maskSelect_lo_1[2175:2168]},
     {maskSplit_maskSelect_lo_1[2167:2160]},
     {maskSplit_maskSelect_lo_1[2159:2152]},
     {maskSplit_maskSelect_lo_1[2151:2144]},
     {maskSplit_maskSelect_lo_1[2143:2136]},
     {maskSplit_maskSelect_lo_1[2135:2128]},
     {maskSplit_maskSelect_lo_1[2127:2120]},
     {maskSplit_maskSelect_lo_1[2119:2112]},
     {maskSplit_maskSelect_lo_1[2111:2104]},
     {maskSplit_maskSelect_lo_1[2103:2096]},
     {maskSplit_maskSelect_lo_1[2095:2088]},
     {maskSplit_maskSelect_lo_1[2087:2080]},
     {maskSplit_maskSelect_lo_1[2079:2072]},
     {maskSplit_maskSelect_lo_1[2071:2064]},
     {maskSplit_maskSelect_lo_1[2063:2056]},
     {maskSplit_maskSelect_lo_1[2055:2048]},
     {maskSplit_maskSelect_lo_1[2047:2040]},
     {maskSplit_maskSelect_lo_1[2039:2032]},
     {maskSplit_maskSelect_lo_1[2031:2024]},
     {maskSplit_maskSelect_lo_1[2023:2016]},
     {maskSplit_maskSelect_lo_1[2015:2008]},
     {maskSplit_maskSelect_lo_1[2007:2000]},
     {maskSplit_maskSelect_lo_1[1999:1992]},
     {maskSplit_maskSelect_lo_1[1991:1984]},
     {maskSplit_maskSelect_lo_1[1983:1976]},
     {maskSplit_maskSelect_lo_1[1975:1968]},
     {maskSplit_maskSelect_lo_1[1967:1960]},
     {maskSplit_maskSelect_lo_1[1959:1952]},
     {maskSplit_maskSelect_lo_1[1951:1944]},
     {maskSplit_maskSelect_lo_1[1943:1936]},
     {maskSplit_maskSelect_lo_1[1935:1928]},
     {maskSplit_maskSelect_lo_1[1927:1920]},
     {maskSplit_maskSelect_lo_1[1919:1912]},
     {maskSplit_maskSelect_lo_1[1911:1904]},
     {maskSplit_maskSelect_lo_1[1903:1896]},
     {maskSplit_maskSelect_lo_1[1895:1888]},
     {maskSplit_maskSelect_lo_1[1887:1880]},
     {maskSplit_maskSelect_lo_1[1879:1872]},
     {maskSplit_maskSelect_lo_1[1871:1864]},
     {maskSplit_maskSelect_lo_1[1863:1856]},
     {maskSplit_maskSelect_lo_1[1855:1848]},
     {maskSplit_maskSelect_lo_1[1847:1840]},
     {maskSplit_maskSelect_lo_1[1839:1832]},
     {maskSplit_maskSelect_lo_1[1831:1824]},
     {maskSplit_maskSelect_lo_1[1823:1816]},
     {maskSplit_maskSelect_lo_1[1815:1808]},
     {maskSplit_maskSelect_lo_1[1807:1800]},
     {maskSplit_maskSelect_lo_1[1799:1792]},
     {maskSplit_maskSelect_lo_1[1791:1784]},
     {maskSplit_maskSelect_lo_1[1783:1776]},
     {maskSplit_maskSelect_lo_1[1775:1768]},
     {maskSplit_maskSelect_lo_1[1767:1760]},
     {maskSplit_maskSelect_lo_1[1759:1752]},
     {maskSplit_maskSelect_lo_1[1751:1744]},
     {maskSplit_maskSelect_lo_1[1743:1736]},
     {maskSplit_maskSelect_lo_1[1735:1728]},
     {maskSplit_maskSelect_lo_1[1727:1720]},
     {maskSplit_maskSelect_lo_1[1719:1712]},
     {maskSplit_maskSelect_lo_1[1711:1704]},
     {maskSplit_maskSelect_lo_1[1703:1696]},
     {maskSplit_maskSelect_lo_1[1695:1688]},
     {maskSplit_maskSelect_lo_1[1687:1680]},
     {maskSplit_maskSelect_lo_1[1679:1672]},
     {maskSplit_maskSelect_lo_1[1671:1664]},
     {maskSplit_maskSelect_lo_1[1663:1656]},
     {maskSplit_maskSelect_lo_1[1655:1648]},
     {maskSplit_maskSelect_lo_1[1647:1640]},
     {maskSplit_maskSelect_lo_1[1639:1632]},
     {maskSplit_maskSelect_lo_1[1631:1624]},
     {maskSplit_maskSelect_lo_1[1623:1616]},
     {maskSplit_maskSelect_lo_1[1615:1608]},
     {maskSplit_maskSelect_lo_1[1607:1600]},
     {maskSplit_maskSelect_lo_1[1599:1592]},
     {maskSplit_maskSelect_lo_1[1591:1584]},
     {maskSplit_maskSelect_lo_1[1583:1576]},
     {maskSplit_maskSelect_lo_1[1575:1568]},
     {maskSplit_maskSelect_lo_1[1567:1560]},
     {maskSplit_maskSelect_lo_1[1559:1552]},
     {maskSplit_maskSelect_lo_1[1551:1544]},
     {maskSplit_maskSelect_lo_1[1543:1536]},
     {maskSplit_maskSelect_lo_1[1535:1528]},
     {maskSplit_maskSelect_lo_1[1527:1520]},
     {maskSplit_maskSelect_lo_1[1519:1512]},
     {maskSplit_maskSelect_lo_1[1511:1504]},
     {maskSplit_maskSelect_lo_1[1503:1496]},
     {maskSplit_maskSelect_lo_1[1495:1488]},
     {maskSplit_maskSelect_lo_1[1487:1480]},
     {maskSplit_maskSelect_lo_1[1479:1472]},
     {maskSplit_maskSelect_lo_1[1471:1464]},
     {maskSplit_maskSelect_lo_1[1463:1456]},
     {maskSplit_maskSelect_lo_1[1455:1448]},
     {maskSplit_maskSelect_lo_1[1447:1440]},
     {maskSplit_maskSelect_lo_1[1439:1432]},
     {maskSplit_maskSelect_lo_1[1431:1424]},
     {maskSplit_maskSelect_lo_1[1423:1416]},
     {maskSplit_maskSelect_lo_1[1415:1408]},
     {maskSplit_maskSelect_lo_1[1407:1400]},
     {maskSplit_maskSelect_lo_1[1399:1392]},
     {maskSplit_maskSelect_lo_1[1391:1384]},
     {maskSplit_maskSelect_lo_1[1383:1376]},
     {maskSplit_maskSelect_lo_1[1375:1368]},
     {maskSplit_maskSelect_lo_1[1367:1360]},
     {maskSplit_maskSelect_lo_1[1359:1352]},
     {maskSplit_maskSelect_lo_1[1351:1344]},
     {maskSplit_maskSelect_lo_1[1343:1336]},
     {maskSplit_maskSelect_lo_1[1335:1328]},
     {maskSplit_maskSelect_lo_1[1327:1320]},
     {maskSplit_maskSelect_lo_1[1319:1312]},
     {maskSplit_maskSelect_lo_1[1311:1304]},
     {maskSplit_maskSelect_lo_1[1303:1296]},
     {maskSplit_maskSelect_lo_1[1295:1288]},
     {maskSplit_maskSelect_lo_1[1287:1280]},
     {maskSplit_maskSelect_lo_1[1279:1272]},
     {maskSplit_maskSelect_lo_1[1271:1264]},
     {maskSplit_maskSelect_lo_1[1263:1256]},
     {maskSplit_maskSelect_lo_1[1255:1248]},
     {maskSplit_maskSelect_lo_1[1247:1240]},
     {maskSplit_maskSelect_lo_1[1239:1232]},
     {maskSplit_maskSelect_lo_1[1231:1224]},
     {maskSplit_maskSelect_lo_1[1223:1216]},
     {maskSplit_maskSelect_lo_1[1215:1208]},
     {maskSplit_maskSelect_lo_1[1207:1200]},
     {maskSplit_maskSelect_lo_1[1199:1192]},
     {maskSplit_maskSelect_lo_1[1191:1184]},
     {maskSplit_maskSelect_lo_1[1183:1176]},
     {maskSplit_maskSelect_lo_1[1175:1168]},
     {maskSplit_maskSelect_lo_1[1167:1160]},
     {maskSplit_maskSelect_lo_1[1159:1152]},
     {maskSplit_maskSelect_lo_1[1151:1144]},
     {maskSplit_maskSelect_lo_1[1143:1136]},
     {maskSplit_maskSelect_lo_1[1135:1128]},
     {maskSplit_maskSelect_lo_1[1127:1120]},
     {maskSplit_maskSelect_lo_1[1119:1112]},
     {maskSplit_maskSelect_lo_1[1111:1104]},
     {maskSplit_maskSelect_lo_1[1103:1096]},
     {maskSplit_maskSelect_lo_1[1095:1088]},
     {maskSplit_maskSelect_lo_1[1087:1080]},
     {maskSplit_maskSelect_lo_1[1079:1072]},
     {maskSplit_maskSelect_lo_1[1071:1064]},
     {maskSplit_maskSelect_lo_1[1063:1056]},
     {maskSplit_maskSelect_lo_1[1055:1048]},
     {maskSplit_maskSelect_lo_1[1047:1040]},
     {maskSplit_maskSelect_lo_1[1039:1032]},
     {maskSplit_maskSelect_lo_1[1031:1024]},
     {maskSplit_maskSelect_lo_1[1023:1016]},
     {maskSplit_maskSelect_lo_1[1015:1008]},
     {maskSplit_maskSelect_lo_1[1007:1000]},
     {maskSplit_maskSelect_lo_1[999:992]},
     {maskSplit_maskSelect_lo_1[991:984]},
     {maskSplit_maskSelect_lo_1[983:976]},
     {maskSplit_maskSelect_lo_1[975:968]},
     {maskSplit_maskSelect_lo_1[967:960]},
     {maskSplit_maskSelect_lo_1[959:952]},
     {maskSplit_maskSelect_lo_1[951:944]},
     {maskSplit_maskSelect_lo_1[943:936]},
     {maskSplit_maskSelect_lo_1[935:928]},
     {maskSplit_maskSelect_lo_1[927:920]},
     {maskSplit_maskSelect_lo_1[919:912]},
     {maskSplit_maskSelect_lo_1[911:904]},
     {maskSplit_maskSelect_lo_1[903:896]},
     {maskSplit_maskSelect_lo_1[895:888]},
     {maskSplit_maskSelect_lo_1[887:880]},
     {maskSplit_maskSelect_lo_1[879:872]},
     {maskSplit_maskSelect_lo_1[871:864]},
     {maskSplit_maskSelect_lo_1[863:856]},
     {maskSplit_maskSelect_lo_1[855:848]},
     {maskSplit_maskSelect_lo_1[847:840]},
     {maskSplit_maskSelect_lo_1[839:832]},
     {maskSplit_maskSelect_lo_1[831:824]},
     {maskSplit_maskSelect_lo_1[823:816]},
     {maskSplit_maskSelect_lo_1[815:808]},
     {maskSplit_maskSelect_lo_1[807:800]},
     {maskSplit_maskSelect_lo_1[799:792]},
     {maskSplit_maskSelect_lo_1[791:784]},
     {maskSplit_maskSelect_lo_1[783:776]},
     {maskSplit_maskSelect_lo_1[775:768]},
     {maskSplit_maskSelect_lo_1[767:760]},
     {maskSplit_maskSelect_lo_1[759:752]},
     {maskSplit_maskSelect_lo_1[751:744]},
     {maskSplit_maskSelect_lo_1[743:736]},
     {maskSplit_maskSelect_lo_1[735:728]},
     {maskSplit_maskSelect_lo_1[727:720]},
     {maskSplit_maskSelect_lo_1[719:712]},
     {maskSplit_maskSelect_lo_1[711:704]},
     {maskSplit_maskSelect_lo_1[703:696]},
     {maskSplit_maskSelect_lo_1[695:688]},
     {maskSplit_maskSelect_lo_1[687:680]},
     {maskSplit_maskSelect_lo_1[679:672]},
     {maskSplit_maskSelect_lo_1[671:664]},
     {maskSplit_maskSelect_lo_1[663:656]},
     {maskSplit_maskSelect_lo_1[655:648]},
     {maskSplit_maskSelect_lo_1[647:640]},
     {maskSplit_maskSelect_lo_1[639:632]},
     {maskSplit_maskSelect_lo_1[631:624]},
     {maskSplit_maskSelect_lo_1[623:616]},
     {maskSplit_maskSelect_lo_1[615:608]},
     {maskSplit_maskSelect_lo_1[607:600]},
     {maskSplit_maskSelect_lo_1[599:592]},
     {maskSplit_maskSelect_lo_1[591:584]},
     {maskSplit_maskSelect_lo_1[583:576]},
     {maskSplit_maskSelect_lo_1[575:568]},
     {maskSplit_maskSelect_lo_1[567:560]},
     {maskSplit_maskSelect_lo_1[559:552]},
     {maskSplit_maskSelect_lo_1[551:544]},
     {maskSplit_maskSelect_lo_1[543:536]},
     {maskSplit_maskSelect_lo_1[535:528]},
     {maskSplit_maskSelect_lo_1[527:520]},
     {maskSplit_maskSelect_lo_1[519:512]},
     {maskSplit_maskSelect_lo_1[511:504]},
     {maskSplit_maskSelect_lo_1[503:496]},
     {maskSplit_maskSelect_lo_1[495:488]},
     {maskSplit_maskSelect_lo_1[487:480]},
     {maskSplit_maskSelect_lo_1[479:472]},
     {maskSplit_maskSelect_lo_1[471:464]},
     {maskSplit_maskSelect_lo_1[463:456]},
     {maskSplit_maskSelect_lo_1[455:448]},
     {maskSplit_maskSelect_lo_1[447:440]},
     {maskSplit_maskSelect_lo_1[439:432]},
     {maskSplit_maskSelect_lo_1[431:424]},
     {maskSplit_maskSelect_lo_1[423:416]},
     {maskSplit_maskSelect_lo_1[415:408]},
     {maskSplit_maskSelect_lo_1[407:400]},
     {maskSplit_maskSelect_lo_1[399:392]},
     {maskSplit_maskSelect_lo_1[391:384]},
     {maskSplit_maskSelect_lo_1[383:376]},
     {maskSplit_maskSelect_lo_1[375:368]},
     {maskSplit_maskSelect_lo_1[367:360]},
     {maskSplit_maskSelect_lo_1[359:352]},
     {maskSplit_maskSelect_lo_1[351:344]},
     {maskSplit_maskSelect_lo_1[343:336]},
     {maskSplit_maskSelect_lo_1[335:328]},
     {maskSplit_maskSelect_lo_1[327:320]},
     {maskSplit_maskSelect_lo_1[319:312]},
     {maskSplit_maskSelect_lo_1[311:304]},
     {maskSplit_maskSelect_lo_1[303:296]},
     {maskSplit_maskSelect_lo_1[295:288]},
     {maskSplit_maskSelect_lo_1[287:280]},
     {maskSplit_maskSelect_lo_1[279:272]},
     {maskSplit_maskSelect_lo_1[271:264]},
     {maskSplit_maskSelect_lo_1[263:256]},
     {maskSplit_maskSelect_lo_1[255:248]},
     {maskSplit_maskSelect_lo_1[247:240]},
     {maskSplit_maskSelect_lo_1[239:232]},
     {maskSplit_maskSelect_lo_1[231:224]},
     {maskSplit_maskSelect_lo_1[223:216]},
     {maskSplit_maskSelect_lo_1[215:208]},
     {maskSplit_maskSelect_lo_1[207:200]},
     {maskSplit_maskSelect_lo_1[199:192]},
     {maskSplit_maskSelect_lo_1[191:184]},
     {maskSplit_maskSelect_lo_1[183:176]},
     {maskSplit_maskSelect_lo_1[175:168]},
     {maskSplit_maskSelect_lo_1[167:160]},
     {maskSplit_maskSelect_lo_1[159:152]},
     {maskSplit_maskSelect_lo_1[151:144]},
     {maskSplit_maskSelect_lo_1[143:136]},
     {maskSplit_maskSelect_lo_1[135:128]},
     {maskSplit_maskSelect_lo_1[127:120]},
     {maskSplit_maskSelect_lo_1[119:112]},
     {maskSplit_maskSelect_lo_1[111:104]},
     {maskSplit_maskSelect_lo_1[103:96]},
     {maskSplit_maskSelect_lo_1[95:88]},
     {maskSplit_maskSelect_lo_1[87:80]},
     {maskSplit_maskSelect_lo_1[79:72]},
     {maskSplit_maskSelect_lo_1[71:64]},
     {maskSplit_maskSelect_lo_1[63:56]},
     {maskSplit_maskSelect_lo_1[55:48]},
     {maskSplit_maskSelect_lo_1[47:40]},
     {maskSplit_maskSelect_lo_1[39:32]},
     {maskSplit_maskSelect_lo_1[31:24]},
     {maskSplit_maskSelect_lo_1[23:16]},
     {maskSplit_maskSelect_lo_1[15:8]},
     {maskSplit_maskSelect_lo_1[7:0]}};
  wire [7:0]         maskSplit_1_2 = (instReg_maskType ? _GEN_145[executeGroupCounter] : 8'hFF) & maskSplit_vlBoundaryCorrection_1;
  wire [3:0]         maskSplit_byteMask_lo_lo_1 = {{2{maskSplit_1_2[1]}}, {2{maskSplit_1_2[0]}}};
  wire [3:0]         maskSplit_byteMask_lo_hi_1 = {{2{maskSplit_1_2[3]}}, {2{maskSplit_1_2[2]}}};
  wire [7:0]         maskSplit_byteMask_lo_1 = {maskSplit_byteMask_lo_hi_1, maskSplit_byteMask_lo_lo_1};
  wire [3:0]         maskSplit_byteMask_hi_lo_1 = {{2{maskSplit_1_2[5]}}, {2{maskSplit_1_2[4]}}};
  wire [3:0]         maskSplit_byteMask_hi_hi_1 = {{2{maskSplit_1_2[7]}}, {2{maskSplit_1_2[6]}}};
  wire [7:0]         maskSplit_byteMask_hi_1 = {maskSplit_byteMask_hi_hi_1, maskSplit_byteMask_hi_lo_1};
  wire [15:0]        maskSplit_1_1 = {maskSplit_byteMask_hi_1, maskSplit_byteMask_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_lo_lo_lo_2 = {maskSplit_maskSelect_lo_lo_lo_lo_lo_lo_hi_2, maskSplit_maskSelect_lo_lo_lo_lo_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_lo_lo_hi_2 = {maskSplit_maskSelect_lo_lo_lo_lo_lo_hi_hi_2, maskSplit_maskSelect_lo_lo_lo_lo_lo_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_lo_lo_lo_lo_lo_2 = {maskSplit_maskSelect_lo_lo_lo_lo_lo_hi_2, maskSplit_maskSelect_lo_lo_lo_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_lo_hi_lo_2 = {maskSplit_maskSelect_lo_lo_lo_lo_hi_lo_hi_2, maskSplit_maskSelect_lo_lo_lo_lo_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_lo_hi_hi_2 = {maskSplit_maskSelect_lo_lo_lo_lo_hi_hi_hi_2, maskSplit_maskSelect_lo_lo_lo_lo_hi_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_lo_lo_lo_lo_hi_2 = {maskSplit_maskSelect_lo_lo_lo_lo_hi_hi_2, maskSplit_maskSelect_lo_lo_lo_lo_hi_lo_2};
  wire [511:0]       maskSplit_maskSelect_lo_lo_lo_lo_2 = {maskSplit_maskSelect_lo_lo_lo_lo_hi_2, maskSplit_maskSelect_lo_lo_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_hi_lo_lo_2 = {maskSplit_maskSelect_lo_lo_lo_hi_lo_lo_hi_2, maskSplit_maskSelect_lo_lo_lo_hi_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_hi_lo_hi_2 = {maskSplit_maskSelect_lo_lo_lo_hi_lo_hi_hi_2, maskSplit_maskSelect_lo_lo_lo_hi_lo_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_lo_lo_lo_hi_lo_2 = {maskSplit_maskSelect_lo_lo_lo_hi_lo_hi_2, maskSplit_maskSelect_lo_lo_lo_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_hi_hi_lo_2 = {maskSplit_maskSelect_lo_lo_lo_hi_hi_lo_hi_2, maskSplit_maskSelect_lo_lo_lo_hi_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_hi_hi_hi_2 = {maskSplit_maskSelect_lo_lo_lo_hi_hi_hi_hi_2, maskSplit_maskSelect_lo_lo_lo_hi_hi_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_lo_lo_lo_hi_hi_2 = {maskSplit_maskSelect_lo_lo_lo_hi_hi_hi_2, maskSplit_maskSelect_lo_lo_lo_hi_hi_lo_2};
  wire [511:0]       maskSplit_maskSelect_lo_lo_lo_hi_2 = {maskSplit_maskSelect_lo_lo_lo_hi_hi_2, maskSplit_maskSelect_lo_lo_lo_hi_lo_2};
  wire [1023:0]      maskSplit_maskSelect_lo_lo_lo_2 = {maskSplit_maskSelect_lo_lo_lo_hi_2, maskSplit_maskSelect_lo_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_lo_lo_lo_2 = {maskSplit_maskSelect_lo_lo_hi_lo_lo_lo_hi_2, maskSplit_maskSelect_lo_lo_hi_lo_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_lo_lo_hi_2 = {maskSplit_maskSelect_lo_lo_hi_lo_lo_hi_hi_2, maskSplit_maskSelect_lo_lo_hi_lo_lo_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_lo_lo_hi_lo_lo_2 = {maskSplit_maskSelect_lo_lo_hi_lo_lo_hi_2, maskSplit_maskSelect_lo_lo_hi_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_lo_hi_lo_2 = {maskSplit_maskSelect_lo_lo_hi_lo_hi_lo_hi_2, maskSplit_maskSelect_lo_lo_hi_lo_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_lo_hi_hi_2 = {maskSplit_maskSelect_lo_lo_hi_lo_hi_hi_hi_2, maskSplit_maskSelect_lo_lo_hi_lo_hi_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_lo_lo_hi_lo_hi_2 = {maskSplit_maskSelect_lo_lo_hi_lo_hi_hi_2, maskSplit_maskSelect_lo_lo_hi_lo_hi_lo_2};
  wire [511:0]       maskSplit_maskSelect_lo_lo_hi_lo_2 = {maskSplit_maskSelect_lo_lo_hi_lo_hi_2, maskSplit_maskSelect_lo_lo_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_hi_lo_lo_2 = {maskSplit_maskSelect_lo_lo_hi_hi_lo_lo_hi_2, maskSplit_maskSelect_lo_lo_hi_hi_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_hi_lo_hi_2 = {maskSplit_maskSelect_lo_lo_hi_hi_lo_hi_hi_2, maskSplit_maskSelect_lo_lo_hi_hi_lo_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_lo_lo_hi_hi_lo_2 = {maskSplit_maskSelect_lo_lo_hi_hi_lo_hi_2, maskSplit_maskSelect_lo_lo_hi_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_hi_hi_lo_2 = {maskSplit_maskSelect_lo_lo_hi_hi_hi_lo_hi_2, maskSplit_maskSelect_lo_lo_hi_hi_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_hi_hi_hi_2 = {maskSplit_maskSelect_lo_lo_hi_hi_hi_hi_hi_2, maskSplit_maskSelect_lo_lo_hi_hi_hi_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_lo_lo_hi_hi_hi_2 = {maskSplit_maskSelect_lo_lo_hi_hi_hi_hi_2, maskSplit_maskSelect_lo_lo_hi_hi_hi_lo_2};
  wire [511:0]       maskSplit_maskSelect_lo_lo_hi_hi_2 = {maskSplit_maskSelect_lo_lo_hi_hi_hi_2, maskSplit_maskSelect_lo_lo_hi_hi_lo_2};
  wire [1023:0]      maskSplit_maskSelect_lo_lo_hi_2 = {maskSplit_maskSelect_lo_lo_hi_hi_2, maskSplit_maskSelect_lo_lo_hi_lo_2};
  wire [2047:0]      maskSplit_maskSelect_lo_lo_2 = {maskSplit_maskSelect_lo_lo_hi_2, maskSplit_maskSelect_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_lo_lo_lo_2 = {maskSplit_maskSelect_lo_hi_lo_lo_lo_lo_hi_2, maskSplit_maskSelect_lo_hi_lo_lo_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_lo_lo_hi_2 = {maskSplit_maskSelect_lo_hi_lo_lo_lo_hi_hi_2, maskSplit_maskSelect_lo_hi_lo_lo_lo_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_lo_hi_lo_lo_lo_2 = {maskSplit_maskSelect_lo_hi_lo_lo_lo_hi_2, maskSplit_maskSelect_lo_hi_lo_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_lo_hi_lo_2 = {maskSplit_maskSelect_lo_hi_lo_lo_hi_lo_hi_2, maskSplit_maskSelect_lo_hi_lo_lo_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_lo_hi_hi_2 = {maskSplit_maskSelect_lo_hi_lo_lo_hi_hi_hi_2, maskSplit_maskSelect_lo_hi_lo_lo_hi_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_lo_hi_lo_lo_hi_2 = {maskSplit_maskSelect_lo_hi_lo_lo_hi_hi_2, maskSplit_maskSelect_lo_hi_lo_lo_hi_lo_2};
  wire [511:0]       maskSplit_maskSelect_lo_hi_lo_lo_2 = {maskSplit_maskSelect_lo_hi_lo_lo_hi_2, maskSplit_maskSelect_lo_hi_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_hi_lo_lo_2 = {maskSplit_maskSelect_lo_hi_lo_hi_lo_lo_hi_2, maskSplit_maskSelect_lo_hi_lo_hi_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_hi_lo_hi_2 = {maskSplit_maskSelect_lo_hi_lo_hi_lo_hi_hi_2, maskSplit_maskSelect_lo_hi_lo_hi_lo_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_lo_hi_lo_hi_lo_2 = {maskSplit_maskSelect_lo_hi_lo_hi_lo_hi_2, maskSplit_maskSelect_lo_hi_lo_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_hi_hi_lo_2 = {maskSplit_maskSelect_lo_hi_lo_hi_hi_lo_hi_2, maskSplit_maskSelect_lo_hi_lo_hi_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_hi_hi_hi_2 = {maskSplit_maskSelect_lo_hi_lo_hi_hi_hi_hi_2, maskSplit_maskSelect_lo_hi_lo_hi_hi_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_lo_hi_lo_hi_hi_2 = {maskSplit_maskSelect_lo_hi_lo_hi_hi_hi_2, maskSplit_maskSelect_lo_hi_lo_hi_hi_lo_2};
  wire [511:0]       maskSplit_maskSelect_lo_hi_lo_hi_2 = {maskSplit_maskSelect_lo_hi_lo_hi_hi_2, maskSplit_maskSelect_lo_hi_lo_hi_lo_2};
  wire [1023:0]      maskSplit_maskSelect_lo_hi_lo_2 = {maskSplit_maskSelect_lo_hi_lo_hi_2, maskSplit_maskSelect_lo_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_lo_lo_lo_2 = {maskSplit_maskSelect_lo_hi_hi_lo_lo_lo_hi_2, maskSplit_maskSelect_lo_hi_hi_lo_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_lo_lo_hi_2 = {maskSplit_maskSelect_lo_hi_hi_lo_lo_hi_hi_2, maskSplit_maskSelect_lo_hi_hi_lo_lo_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_lo_hi_hi_lo_lo_2 = {maskSplit_maskSelect_lo_hi_hi_lo_lo_hi_2, maskSplit_maskSelect_lo_hi_hi_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_lo_hi_lo_2 = {maskSplit_maskSelect_lo_hi_hi_lo_hi_lo_hi_2, maskSplit_maskSelect_lo_hi_hi_lo_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_lo_hi_hi_2 = {maskSplit_maskSelect_lo_hi_hi_lo_hi_hi_hi_2, maskSplit_maskSelect_lo_hi_hi_lo_hi_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_lo_hi_hi_lo_hi_2 = {maskSplit_maskSelect_lo_hi_hi_lo_hi_hi_2, maskSplit_maskSelect_lo_hi_hi_lo_hi_lo_2};
  wire [511:0]       maskSplit_maskSelect_lo_hi_hi_lo_2 = {maskSplit_maskSelect_lo_hi_hi_lo_hi_2, maskSplit_maskSelect_lo_hi_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_hi_lo_lo_2 = {maskSplit_maskSelect_lo_hi_hi_hi_lo_lo_hi_2, maskSplit_maskSelect_lo_hi_hi_hi_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_hi_lo_hi_2 = {maskSplit_maskSelect_lo_hi_hi_hi_lo_hi_hi_2, maskSplit_maskSelect_lo_hi_hi_hi_lo_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_lo_hi_hi_hi_lo_2 = {maskSplit_maskSelect_lo_hi_hi_hi_lo_hi_2, maskSplit_maskSelect_lo_hi_hi_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_hi_hi_lo_2 = {maskSplit_maskSelect_lo_hi_hi_hi_hi_lo_hi_2, maskSplit_maskSelect_lo_hi_hi_hi_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_hi_hi_hi_2 = {maskSplit_maskSelect_lo_hi_hi_hi_hi_hi_hi_2, maskSplit_maskSelect_lo_hi_hi_hi_hi_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_lo_hi_hi_hi_hi_2 = {maskSplit_maskSelect_lo_hi_hi_hi_hi_hi_2, maskSplit_maskSelect_lo_hi_hi_hi_hi_lo_2};
  wire [511:0]       maskSplit_maskSelect_lo_hi_hi_hi_2 = {maskSplit_maskSelect_lo_hi_hi_hi_hi_2, maskSplit_maskSelect_lo_hi_hi_hi_lo_2};
  wire [1023:0]      maskSplit_maskSelect_lo_hi_hi_2 = {maskSplit_maskSelect_lo_hi_hi_hi_2, maskSplit_maskSelect_lo_hi_hi_lo_2};
  wire [2047:0]      maskSplit_maskSelect_lo_hi_2 = {maskSplit_maskSelect_lo_hi_hi_2, maskSplit_maskSelect_lo_hi_lo_2};
  wire [4095:0]      maskSplit_maskSelect_lo_2 = {maskSplit_maskSelect_lo_hi_2, maskSplit_maskSelect_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_lo_lo_lo_2 = {maskSplit_maskSelect_hi_lo_lo_lo_lo_lo_hi_2, maskSplit_maskSelect_hi_lo_lo_lo_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_lo_lo_hi_2 = {maskSplit_maskSelect_hi_lo_lo_lo_lo_hi_hi_2, maskSplit_maskSelect_hi_lo_lo_lo_lo_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_hi_lo_lo_lo_lo_2 = {maskSplit_maskSelect_hi_lo_lo_lo_lo_hi_2, maskSplit_maskSelect_hi_lo_lo_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_lo_hi_lo_2 = {maskSplit_maskSelect_hi_lo_lo_lo_hi_lo_hi_2, maskSplit_maskSelect_hi_lo_lo_lo_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_lo_hi_hi_2 = {maskSplit_maskSelect_hi_lo_lo_lo_hi_hi_hi_2, maskSplit_maskSelect_hi_lo_lo_lo_hi_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_hi_lo_lo_lo_hi_2 = {maskSplit_maskSelect_hi_lo_lo_lo_hi_hi_2, maskSplit_maskSelect_hi_lo_lo_lo_hi_lo_2};
  wire [511:0]       maskSplit_maskSelect_hi_lo_lo_lo_2 = {maskSplit_maskSelect_hi_lo_lo_lo_hi_2, maskSplit_maskSelect_hi_lo_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_hi_lo_lo_2 = {maskSplit_maskSelect_hi_lo_lo_hi_lo_lo_hi_2, maskSplit_maskSelect_hi_lo_lo_hi_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_hi_lo_hi_2 = {maskSplit_maskSelect_hi_lo_lo_hi_lo_hi_hi_2, maskSplit_maskSelect_hi_lo_lo_hi_lo_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_hi_lo_lo_hi_lo_2 = {maskSplit_maskSelect_hi_lo_lo_hi_lo_hi_2, maskSplit_maskSelect_hi_lo_lo_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_hi_hi_lo_2 = {maskSplit_maskSelect_hi_lo_lo_hi_hi_lo_hi_2, maskSplit_maskSelect_hi_lo_lo_hi_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_hi_hi_hi_2 = {maskSplit_maskSelect_hi_lo_lo_hi_hi_hi_hi_2, maskSplit_maskSelect_hi_lo_lo_hi_hi_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_hi_lo_lo_hi_hi_2 = {maskSplit_maskSelect_hi_lo_lo_hi_hi_hi_2, maskSplit_maskSelect_hi_lo_lo_hi_hi_lo_2};
  wire [511:0]       maskSplit_maskSelect_hi_lo_lo_hi_2 = {maskSplit_maskSelect_hi_lo_lo_hi_hi_2, maskSplit_maskSelect_hi_lo_lo_hi_lo_2};
  wire [1023:0]      maskSplit_maskSelect_hi_lo_lo_2 = {maskSplit_maskSelect_hi_lo_lo_hi_2, maskSplit_maskSelect_hi_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_lo_lo_lo_2 = {maskSplit_maskSelect_hi_lo_hi_lo_lo_lo_hi_2, maskSplit_maskSelect_hi_lo_hi_lo_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_lo_lo_hi_2 = {maskSplit_maskSelect_hi_lo_hi_lo_lo_hi_hi_2, maskSplit_maskSelect_hi_lo_hi_lo_lo_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_hi_lo_hi_lo_lo_2 = {maskSplit_maskSelect_hi_lo_hi_lo_lo_hi_2, maskSplit_maskSelect_hi_lo_hi_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_lo_hi_lo_2 = {maskSplit_maskSelect_hi_lo_hi_lo_hi_lo_hi_2, maskSplit_maskSelect_hi_lo_hi_lo_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_lo_hi_hi_2 = {maskSplit_maskSelect_hi_lo_hi_lo_hi_hi_hi_2, maskSplit_maskSelect_hi_lo_hi_lo_hi_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_hi_lo_hi_lo_hi_2 = {maskSplit_maskSelect_hi_lo_hi_lo_hi_hi_2, maskSplit_maskSelect_hi_lo_hi_lo_hi_lo_2};
  wire [511:0]       maskSplit_maskSelect_hi_lo_hi_lo_2 = {maskSplit_maskSelect_hi_lo_hi_lo_hi_2, maskSplit_maskSelect_hi_lo_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_hi_lo_lo_2 = {maskSplit_maskSelect_hi_lo_hi_hi_lo_lo_hi_2, maskSplit_maskSelect_hi_lo_hi_hi_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_hi_lo_hi_2 = {maskSplit_maskSelect_hi_lo_hi_hi_lo_hi_hi_2, maskSplit_maskSelect_hi_lo_hi_hi_lo_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_hi_lo_hi_hi_lo_2 = {maskSplit_maskSelect_hi_lo_hi_hi_lo_hi_2, maskSplit_maskSelect_hi_lo_hi_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_hi_hi_lo_2 = {maskSplit_maskSelect_hi_lo_hi_hi_hi_lo_hi_2, maskSplit_maskSelect_hi_lo_hi_hi_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_hi_hi_hi_2 = {maskSplit_maskSelect_hi_lo_hi_hi_hi_hi_hi_2, maskSplit_maskSelect_hi_lo_hi_hi_hi_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_hi_lo_hi_hi_hi_2 = {maskSplit_maskSelect_hi_lo_hi_hi_hi_hi_2, maskSplit_maskSelect_hi_lo_hi_hi_hi_lo_2};
  wire [511:0]       maskSplit_maskSelect_hi_lo_hi_hi_2 = {maskSplit_maskSelect_hi_lo_hi_hi_hi_2, maskSplit_maskSelect_hi_lo_hi_hi_lo_2};
  wire [1023:0]      maskSplit_maskSelect_hi_lo_hi_2 = {maskSplit_maskSelect_hi_lo_hi_hi_2, maskSplit_maskSelect_hi_lo_hi_lo_2};
  wire [2047:0]      maskSplit_maskSelect_hi_lo_2 = {maskSplit_maskSelect_hi_lo_hi_2, maskSplit_maskSelect_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_lo_lo_lo_2 = {maskSplit_maskSelect_hi_hi_lo_lo_lo_lo_hi_2, maskSplit_maskSelect_hi_hi_lo_lo_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_lo_lo_hi_2 = {maskSplit_maskSelect_hi_hi_lo_lo_lo_hi_hi_2, maskSplit_maskSelect_hi_hi_lo_lo_lo_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_hi_hi_lo_lo_lo_2 = {maskSplit_maskSelect_hi_hi_lo_lo_lo_hi_2, maskSplit_maskSelect_hi_hi_lo_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_lo_hi_lo_2 = {maskSplit_maskSelect_hi_hi_lo_lo_hi_lo_hi_2, maskSplit_maskSelect_hi_hi_lo_lo_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_lo_hi_hi_2 = {maskSplit_maskSelect_hi_hi_lo_lo_hi_hi_hi_2, maskSplit_maskSelect_hi_hi_lo_lo_hi_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_hi_hi_lo_lo_hi_2 = {maskSplit_maskSelect_hi_hi_lo_lo_hi_hi_2, maskSplit_maskSelect_hi_hi_lo_lo_hi_lo_2};
  wire [511:0]       maskSplit_maskSelect_hi_hi_lo_lo_2 = {maskSplit_maskSelect_hi_hi_lo_lo_hi_2, maskSplit_maskSelect_hi_hi_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_hi_lo_lo_2 = {maskSplit_maskSelect_hi_hi_lo_hi_lo_lo_hi_2, maskSplit_maskSelect_hi_hi_lo_hi_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_hi_lo_hi_2 = {maskSplit_maskSelect_hi_hi_lo_hi_lo_hi_hi_2, maskSplit_maskSelect_hi_hi_lo_hi_lo_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_hi_hi_lo_hi_lo_2 = {maskSplit_maskSelect_hi_hi_lo_hi_lo_hi_2, maskSplit_maskSelect_hi_hi_lo_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_hi_hi_lo_2 = {maskSplit_maskSelect_hi_hi_lo_hi_hi_lo_hi_2, maskSplit_maskSelect_hi_hi_lo_hi_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_hi_hi_hi_2 = {maskSplit_maskSelect_hi_hi_lo_hi_hi_hi_hi_2, maskSplit_maskSelect_hi_hi_lo_hi_hi_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_hi_hi_lo_hi_hi_2 = {maskSplit_maskSelect_hi_hi_lo_hi_hi_hi_2, maskSplit_maskSelect_hi_hi_lo_hi_hi_lo_2};
  wire [511:0]       maskSplit_maskSelect_hi_hi_lo_hi_2 = {maskSplit_maskSelect_hi_hi_lo_hi_hi_2, maskSplit_maskSelect_hi_hi_lo_hi_lo_2};
  wire [1023:0]      maskSplit_maskSelect_hi_hi_lo_2 = {maskSplit_maskSelect_hi_hi_lo_hi_2, maskSplit_maskSelect_hi_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_lo_lo_lo_2 = {maskSplit_maskSelect_hi_hi_hi_lo_lo_lo_hi_2, maskSplit_maskSelect_hi_hi_hi_lo_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_lo_lo_hi_2 = {maskSplit_maskSelect_hi_hi_hi_lo_lo_hi_hi_2, maskSplit_maskSelect_hi_hi_hi_lo_lo_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_hi_hi_hi_lo_lo_2 = {maskSplit_maskSelect_hi_hi_hi_lo_lo_hi_2, maskSplit_maskSelect_hi_hi_hi_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_lo_hi_lo_2 = {maskSplit_maskSelect_hi_hi_hi_lo_hi_lo_hi_2, maskSplit_maskSelect_hi_hi_hi_lo_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_lo_hi_hi_2 = {maskSplit_maskSelect_hi_hi_hi_lo_hi_hi_hi_2, maskSplit_maskSelect_hi_hi_hi_lo_hi_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_hi_hi_hi_lo_hi_2 = {maskSplit_maskSelect_hi_hi_hi_lo_hi_hi_2, maskSplit_maskSelect_hi_hi_hi_lo_hi_lo_2};
  wire [511:0]       maskSplit_maskSelect_hi_hi_hi_lo_2 = {maskSplit_maskSelect_hi_hi_hi_lo_hi_2, maskSplit_maskSelect_hi_hi_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_hi_lo_lo_2 = {maskSplit_maskSelect_hi_hi_hi_hi_lo_lo_hi_2, maskSplit_maskSelect_hi_hi_hi_hi_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_hi_lo_hi_2 = {maskSplit_maskSelect_hi_hi_hi_hi_lo_hi_hi_2, maskSplit_maskSelect_hi_hi_hi_hi_lo_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_hi_hi_hi_hi_lo_2 = {maskSplit_maskSelect_hi_hi_hi_hi_lo_hi_2, maskSplit_maskSelect_hi_hi_hi_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_hi_hi_lo_2 = {maskSplit_maskSelect_hi_hi_hi_hi_hi_lo_hi_2, maskSplit_maskSelect_hi_hi_hi_hi_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_hi_hi_hi_2 = {maskSplit_maskSelect_hi_hi_hi_hi_hi_hi_hi_2, maskSplit_maskSelect_hi_hi_hi_hi_hi_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_hi_hi_hi_hi_hi_2 = {maskSplit_maskSelect_hi_hi_hi_hi_hi_hi_2, maskSplit_maskSelect_hi_hi_hi_hi_hi_lo_2};
  wire [511:0]       maskSplit_maskSelect_hi_hi_hi_hi_2 = {maskSplit_maskSelect_hi_hi_hi_hi_hi_2, maskSplit_maskSelect_hi_hi_hi_hi_lo_2};
  wire [1023:0]      maskSplit_maskSelect_hi_hi_hi_2 = {maskSplit_maskSelect_hi_hi_hi_hi_2, maskSplit_maskSelect_hi_hi_hi_lo_2};
  wire [2047:0]      maskSplit_maskSelect_hi_hi_2 = {maskSplit_maskSelect_hi_hi_hi_2, maskSplit_maskSelect_hi_hi_lo_2};
  wire [4095:0]      maskSplit_maskSelect_hi_2 = {maskSplit_maskSelect_hi_hi_2, maskSplit_maskSelect_hi_lo_2};
  wire               maskSplit_vlMisAlign_2;
  assign maskSplit_vlMisAlign_2 = |(instReg_vl[1:0]);
  wire [11:0]        maskSplit_lastexecuteGroup_2 = instReg_vl[13:2] - {11'h0, ~maskSplit_vlMisAlign_2};
  wire [11:0]        _GEN_146 = {2'h0, executeGroupCounter};
  wire               maskSplit_isVlBoundary_2 = _GEN_146 == maskSplit_lastexecuteGroup_2;
  wire               maskSplit_validExecuteGroup_2 = _GEN_146 <= maskSplit_lastexecuteGroup_2;
  wire [3:0]         _maskSplit_vlBoundaryCorrection_T_40 = _maskSplit_vlBoundaryCorrection_T_37 | {_maskSplit_vlBoundaryCorrection_T_37[2:0], 1'h0};
  wire [3:0]         maskSplit_vlBoundaryCorrection_2 =
    ~({4{maskSplit_vlMisAlign_2 & maskSplit_isVlBoundary_2}} & (_maskSplit_vlBoundaryCorrection_T_40 | {_maskSplit_vlBoundaryCorrection_T_40[1:0], 2'h0})) & {4{maskSplit_validExecuteGroup_2}};
  wire [1023:0][3:0] _GEN_147 =
    {{maskSplit_maskSelect_lo_2[4095:4092]},
     {maskSplit_maskSelect_lo_2[4091:4088]},
     {maskSplit_maskSelect_lo_2[4087:4084]},
     {maskSplit_maskSelect_lo_2[4083:4080]},
     {maskSplit_maskSelect_lo_2[4079:4076]},
     {maskSplit_maskSelect_lo_2[4075:4072]},
     {maskSplit_maskSelect_lo_2[4071:4068]},
     {maskSplit_maskSelect_lo_2[4067:4064]},
     {maskSplit_maskSelect_lo_2[4063:4060]},
     {maskSplit_maskSelect_lo_2[4059:4056]},
     {maskSplit_maskSelect_lo_2[4055:4052]},
     {maskSplit_maskSelect_lo_2[4051:4048]},
     {maskSplit_maskSelect_lo_2[4047:4044]},
     {maskSplit_maskSelect_lo_2[4043:4040]},
     {maskSplit_maskSelect_lo_2[4039:4036]},
     {maskSplit_maskSelect_lo_2[4035:4032]},
     {maskSplit_maskSelect_lo_2[4031:4028]},
     {maskSplit_maskSelect_lo_2[4027:4024]},
     {maskSplit_maskSelect_lo_2[4023:4020]},
     {maskSplit_maskSelect_lo_2[4019:4016]},
     {maskSplit_maskSelect_lo_2[4015:4012]},
     {maskSplit_maskSelect_lo_2[4011:4008]},
     {maskSplit_maskSelect_lo_2[4007:4004]},
     {maskSplit_maskSelect_lo_2[4003:4000]},
     {maskSplit_maskSelect_lo_2[3999:3996]},
     {maskSplit_maskSelect_lo_2[3995:3992]},
     {maskSplit_maskSelect_lo_2[3991:3988]},
     {maskSplit_maskSelect_lo_2[3987:3984]},
     {maskSplit_maskSelect_lo_2[3983:3980]},
     {maskSplit_maskSelect_lo_2[3979:3976]},
     {maskSplit_maskSelect_lo_2[3975:3972]},
     {maskSplit_maskSelect_lo_2[3971:3968]},
     {maskSplit_maskSelect_lo_2[3967:3964]},
     {maskSplit_maskSelect_lo_2[3963:3960]},
     {maskSplit_maskSelect_lo_2[3959:3956]},
     {maskSplit_maskSelect_lo_2[3955:3952]},
     {maskSplit_maskSelect_lo_2[3951:3948]},
     {maskSplit_maskSelect_lo_2[3947:3944]},
     {maskSplit_maskSelect_lo_2[3943:3940]},
     {maskSplit_maskSelect_lo_2[3939:3936]},
     {maskSplit_maskSelect_lo_2[3935:3932]},
     {maskSplit_maskSelect_lo_2[3931:3928]},
     {maskSplit_maskSelect_lo_2[3927:3924]},
     {maskSplit_maskSelect_lo_2[3923:3920]},
     {maskSplit_maskSelect_lo_2[3919:3916]},
     {maskSplit_maskSelect_lo_2[3915:3912]},
     {maskSplit_maskSelect_lo_2[3911:3908]},
     {maskSplit_maskSelect_lo_2[3907:3904]},
     {maskSplit_maskSelect_lo_2[3903:3900]},
     {maskSplit_maskSelect_lo_2[3899:3896]},
     {maskSplit_maskSelect_lo_2[3895:3892]},
     {maskSplit_maskSelect_lo_2[3891:3888]},
     {maskSplit_maskSelect_lo_2[3887:3884]},
     {maskSplit_maskSelect_lo_2[3883:3880]},
     {maskSplit_maskSelect_lo_2[3879:3876]},
     {maskSplit_maskSelect_lo_2[3875:3872]},
     {maskSplit_maskSelect_lo_2[3871:3868]},
     {maskSplit_maskSelect_lo_2[3867:3864]},
     {maskSplit_maskSelect_lo_2[3863:3860]},
     {maskSplit_maskSelect_lo_2[3859:3856]},
     {maskSplit_maskSelect_lo_2[3855:3852]},
     {maskSplit_maskSelect_lo_2[3851:3848]},
     {maskSplit_maskSelect_lo_2[3847:3844]},
     {maskSplit_maskSelect_lo_2[3843:3840]},
     {maskSplit_maskSelect_lo_2[3839:3836]},
     {maskSplit_maskSelect_lo_2[3835:3832]},
     {maskSplit_maskSelect_lo_2[3831:3828]},
     {maskSplit_maskSelect_lo_2[3827:3824]},
     {maskSplit_maskSelect_lo_2[3823:3820]},
     {maskSplit_maskSelect_lo_2[3819:3816]},
     {maskSplit_maskSelect_lo_2[3815:3812]},
     {maskSplit_maskSelect_lo_2[3811:3808]},
     {maskSplit_maskSelect_lo_2[3807:3804]},
     {maskSplit_maskSelect_lo_2[3803:3800]},
     {maskSplit_maskSelect_lo_2[3799:3796]},
     {maskSplit_maskSelect_lo_2[3795:3792]},
     {maskSplit_maskSelect_lo_2[3791:3788]},
     {maskSplit_maskSelect_lo_2[3787:3784]},
     {maskSplit_maskSelect_lo_2[3783:3780]},
     {maskSplit_maskSelect_lo_2[3779:3776]},
     {maskSplit_maskSelect_lo_2[3775:3772]},
     {maskSplit_maskSelect_lo_2[3771:3768]},
     {maskSplit_maskSelect_lo_2[3767:3764]},
     {maskSplit_maskSelect_lo_2[3763:3760]},
     {maskSplit_maskSelect_lo_2[3759:3756]},
     {maskSplit_maskSelect_lo_2[3755:3752]},
     {maskSplit_maskSelect_lo_2[3751:3748]},
     {maskSplit_maskSelect_lo_2[3747:3744]},
     {maskSplit_maskSelect_lo_2[3743:3740]},
     {maskSplit_maskSelect_lo_2[3739:3736]},
     {maskSplit_maskSelect_lo_2[3735:3732]},
     {maskSplit_maskSelect_lo_2[3731:3728]},
     {maskSplit_maskSelect_lo_2[3727:3724]},
     {maskSplit_maskSelect_lo_2[3723:3720]},
     {maskSplit_maskSelect_lo_2[3719:3716]},
     {maskSplit_maskSelect_lo_2[3715:3712]},
     {maskSplit_maskSelect_lo_2[3711:3708]},
     {maskSplit_maskSelect_lo_2[3707:3704]},
     {maskSplit_maskSelect_lo_2[3703:3700]},
     {maskSplit_maskSelect_lo_2[3699:3696]},
     {maskSplit_maskSelect_lo_2[3695:3692]},
     {maskSplit_maskSelect_lo_2[3691:3688]},
     {maskSplit_maskSelect_lo_2[3687:3684]},
     {maskSplit_maskSelect_lo_2[3683:3680]},
     {maskSplit_maskSelect_lo_2[3679:3676]},
     {maskSplit_maskSelect_lo_2[3675:3672]},
     {maskSplit_maskSelect_lo_2[3671:3668]},
     {maskSplit_maskSelect_lo_2[3667:3664]},
     {maskSplit_maskSelect_lo_2[3663:3660]},
     {maskSplit_maskSelect_lo_2[3659:3656]},
     {maskSplit_maskSelect_lo_2[3655:3652]},
     {maskSplit_maskSelect_lo_2[3651:3648]},
     {maskSplit_maskSelect_lo_2[3647:3644]},
     {maskSplit_maskSelect_lo_2[3643:3640]},
     {maskSplit_maskSelect_lo_2[3639:3636]},
     {maskSplit_maskSelect_lo_2[3635:3632]},
     {maskSplit_maskSelect_lo_2[3631:3628]},
     {maskSplit_maskSelect_lo_2[3627:3624]},
     {maskSplit_maskSelect_lo_2[3623:3620]},
     {maskSplit_maskSelect_lo_2[3619:3616]},
     {maskSplit_maskSelect_lo_2[3615:3612]},
     {maskSplit_maskSelect_lo_2[3611:3608]},
     {maskSplit_maskSelect_lo_2[3607:3604]},
     {maskSplit_maskSelect_lo_2[3603:3600]},
     {maskSplit_maskSelect_lo_2[3599:3596]},
     {maskSplit_maskSelect_lo_2[3595:3592]},
     {maskSplit_maskSelect_lo_2[3591:3588]},
     {maskSplit_maskSelect_lo_2[3587:3584]},
     {maskSplit_maskSelect_lo_2[3583:3580]},
     {maskSplit_maskSelect_lo_2[3579:3576]},
     {maskSplit_maskSelect_lo_2[3575:3572]},
     {maskSplit_maskSelect_lo_2[3571:3568]},
     {maskSplit_maskSelect_lo_2[3567:3564]},
     {maskSplit_maskSelect_lo_2[3563:3560]},
     {maskSplit_maskSelect_lo_2[3559:3556]},
     {maskSplit_maskSelect_lo_2[3555:3552]},
     {maskSplit_maskSelect_lo_2[3551:3548]},
     {maskSplit_maskSelect_lo_2[3547:3544]},
     {maskSplit_maskSelect_lo_2[3543:3540]},
     {maskSplit_maskSelect_lo_2[3539:3536]},
     {maskSplit_maskSelect_lo_2[3535:3532]},
     {maskSplit_maskSelect_lo_2[3531:3528]},
     {maskSplit_maskSelect_lo_2[3527:3524]},
     {maskSplit_maskSelect_lo_2[3523:3520]},
     {maskSplit_maskSelect_lo_2[3519:3516]},
     {maskSplit_maskSelect_lo_2[3515:3512]},
     {maskSplit_maskSelect_lo_2[3511:3508]},
     {maskSplit_maskSelect_lo_2[3507:3504]},
     {maskSplit_maskSelect_lo_2[3503:3500]},
     {maskSplit_maskSelect_lo_2[3499:3496]},
     {maskSplit_maskSelect_lo_2[3495:3492]},
     {maskSplit_maskSelect_lo_2[3491:3488]},
     {maskSplit_maskSelect_lo_2[3487:3484]},
     {maskSplit_maskSelect_lo_2[3483:3480]},
     {maskSplit_maskSelect_lo_2[3479:3476]},
     {maskSplit_maskSelect_lo_2[3475:3472]},
     {maskSplit_maskSelect_lo_2[3471:3468]},
     {maskSplit_maskSelect_lo_2[3467:3464]},
     {maskSplit_maskSelect_lo_2[3463:3460]},
     {maskSplit_maskSelect_lo_2[3459:3456]},
     {maskSplit_maskSelect_lo_2[3455:3452]},
     {maskSplit_maskSelect_lo_2[3451:3448]},
     {maskSplit_maskSelect_lo_2[3447:3444]},
     {maskSplit_maskSelect_lo_2[3443:3440]},
     {maskSplit_maskSelect_lo_2[3439:3436]},
     {maskSplit_maskSelect_lo_2[3435:3432]},
     {maskSplit_maskSelect_lo_2[3431:3428]},
     {maskSplit_maskSelect_lo_2[3427:3424]},
     {maskSplit_maskSelect_lo_2[3423:3420]},
     {maskSplit_maskSelect_lo_2[3419:3416]},
     {maskSplit_maskSelect_lo_2[3415:3412]},
     {maskSplit_maskSelect_lo_2[3411:3408]},
     {maskSplit_maskSelect_lo_2[3407:3404]},
     {maskSplit_maskSelect_lo_2[3403:3400]},
     {maskSplit_maskSelect_lo_2[3399:3396]},
     {maskSplit_maskSelect_lo_2[3395:3392]},
     {maskSplit_maskSelect_lo_2[3391:3388]},
     {maskSplit_maskSelect_lo_2[3387:3384]},
     {maskSplit_maskSelect_lo_2[3383:3380]},
     {maskSplit_maskSelect_lo_2[3379:3376]},
     {maskSplit_maskSelect_lo_2[3375:3372]},
     {maskSplit_maskSelect_lo_2[3371:3368]},
     {maskSplit_maskSelect_lo_2[3367:3364]},
     {maskSplit_maskSelect_lo_2[3363:3360]},
     {maskSplit_maskSelect_lo_2[3359:3356]},
     {maskSplit_maskSelect_lo_2[3355:3352]},
     {maskSplit_maskSelect_lo_2[3351:3348]},
     {maskSplit_maskSelect_lo_2[3347:3344]},
     {maskSplit_maskSelect_lo_2[3343:3340]},
     {maskSplit_maskSelect_lo_2[3339:3336]},
     {maskSplit_maskSelect_lo_2[3335:3332]},
     {maskSplit_maskSelect_lo_2[3331:3328]},
     {maskSplit_maskSelect_lo_2[3327:3324]},
     {maskSplit_maskSelect_lo_2[3323:3320]},
     {maskSplit_maskSelect_lo_2[3319:3316]},
     {maskSplit_maskSelect_lo_2[3315:3312]},
     {maskSplit_maskSelect_lo_2[3311:3308]},
     {maskSplit_maskSelect_lo_2[3307:3304]},
     {maskSplit_maskSelect_lo_2[3303:3300]},
     {maskSplit_maskSelect_lo_2[3299:3296]},
     {maskSplit_maskSelect_lo_2[3295:3292]},
     {maskSplit_maskSelect_lo_2[3291:3288]},
     {maskSplit_maskSelect_lo_2[3287:3284]},
     {maskSplit_maskSelect_lo_2[3283:3280]},
     {maskSplit_maskSelect_lo_2[3279:3276]},
     {maskSplit_maskSelect_lo_2[3275:3272]},
     {maskSplit_maskSelect_lo_2[3271:3268]},
     {maskSplit_maskSelect_lo_2[3267:3264]},
     {maskSplit_maskSelect_lo_2[3263:3260]},
     {maskSplit_maskSelect_lo_2[3259:3256]},
     {maskSplit_maskSelect_lo_2[3255:3252]},
     {maskSplit_maskSelect_lo_2[3251:3248]},
     {maskSplit_maskSelect_lo_2[3247:3244]},
     {maskSplit_maskSelect_lo_2[3243:3240]},
     {maskSplit_maskSelect_lo_2[3239:3236]},
     {maskSplit_maskSelect_lo_2[3235:3232]},
     {maskSplit_maskSelect_lo_2[3231:3228]},
     {maskSplit_maskSelect_lo_2[3227:3224]},
     {maskSplit_maskSelect_lo_2[3223:3220]},
     {maskSplit_maskSelect_lo_2[3219:3216]},
     {maskSplit_maskSelect_lo_2[3215:3212]},
     {maskSplit_maskSelect_lo_2[3211:3208]},
     {maskSplit_maskSelect_lo_2[3207:3204]},
     {maskSplit_maskSelect_lo_2[3203:3200]},
     {maskSplit_maskSelect_lo_2[3199:3196]},
     {maskSplit_maskSelect_lo_2[3195:3192]},
     {maskSplit_maskSelect_lo_2[3191:3188]},
     {maskSplit_maskSelect_lo_2[3187:3184]},
     {maskSplit_maskSelect_lo_2[3183:3180]},
     {maskSplit_maskSelect_lo_2[3179:3176]},
     {maskSplit_maskSelect_lo_2[3175:3172]},
     {maskSplit_maskSelect_lo_2[3171:3168]},
     {maskSplit_maskSelect_lo_2[3167:3164]},
     {maskSplit_maskSelect_lo_2[3163:3160]},
     {maskSplit_maskSelect_lo_2[3159:3156]},
     {maskSplit_maskSelect_lo_2[3155:3152]},
     {maskSplit_maskSelect_lo_2[3151:3148]},
     {maskSplit_maskSelect_lo_2[3147:3144]},
     {maskSplit_maskSelect_lo_2[3143:3140]},
     {maskSplit_maskSelect_lo_2[3139:3136]},
     {maskSplit_maskSelect_lo_2[3135:3132]},
     {maskSplit_maskSelect_lo_2[3131:3128]},
     {maskSplit_maskSelect_lo_2[3127:3124]},
     {maskSplit_maskSelect_lo_2[3123:3120]},
     {maskSplit_maskSelect_lo_2[3119:3116]},
     {maskSplit_maskSelect_lo_2[3115:3112]},
     {maskSplit_maskSelect_lo_2[3111:3108]},
     {maskSplit_maskSelect_lo_2[3107:3104]},
     {maskSplit_maskSelect_lo_2[3103:3100]},
     {maskSplit_maskSelect_lo_2[3099:3096]},
     {maskSplit_maskSelect_lo_2[3095:3092]},
     {maskSplit_maskSelect_lo_2[3091:3088]},
     {maskSplit_maskSelect_lo_2[3087:3084]},
     {maskSplit_maskSelect_lo_2[3083:3080]},
     {maskSplit_maskSelect_lo_2[3079:3076]},
     {maskSplit_maskSelect_lo_2[3075:3072]},
     {maskSplit_maskSelect_lo_2[3071:3068]},
     {maskSplit_maskSelect_lo_2[3067:3064]},
     {maskSplit_maskSelect_lo_2[3063:3060]},
     {maskSplit_maskSelect_lo_2[3059:3056]},
     {maskSplit_maskSelect_lo_2[3055:3052]},
     {maskSplit_maskSelect_lo_2[3051:3048]},
     {maskSplit_maskSelect_lo_2[3047:3044]},
     {maskSplit_maskSelect_lo_2[3043:3040]},
     {maskSplit_maskSelect_lo_2[3039:3036]},
     {maskSplit_maskSelect_lo_2[3035:3032]},
     {maskSplit_maskSelect_lo_2[3031:3028]},
     {maskSplit_maskSelect_lo_2[3027:3024]},
     {maskSplit_maskSelect_lo_2[3023:3020]},
     {maskSplit_maskSelect_lo_2[3019:3016]},
     {maskSplit_maskSelect_lo_2[3015:3012]},
     {maskSplit_maskSelect_lo_2[3011:3008]},
     {maskSplit_maskSelect_lo_2[3007:3004]},
     {maskSplit_maskSelect_lo_2[3003:3000]},
     {maskSplit_maskSelect_lo_2[2999:2996]},
     {maskSplit_maskSelect_lo_2[2995:2992]},
     {maskSplit_maskSelect_lo_2[2991:2988]},
     {maskSplit_maskSelect_lo_2[2987:2984]},
     {maskSplit_maskSelect_lo_2[2983:2980]},
     {maskSplit_maskSelect_lo_2[2979:2976]},
     {maskSplit_maskSelect_lo_2[2975:2972]},
     {maskSplit_maskSelect_lo_2[2971:2968]},
     {maskSplit_maskSelect_lo_2[2967:2964]},
     {maskSplit_maskSelect_lo_2[2963:2960]},
     {maskSplit_maskSelect_lo_2[2959:2956]},
     {maskSplit_maskSelect_lo_2[2955:2952]},
     {maskSplit_maskSelect_lo_2[2951:2948]},
     {maskSplit_maskSelect_lo_2[2947:2944]},
     {maskSplit_maskSelect_lo_2[2943:2940]},
     {maskSplit_maskSelect_lo_2[2939:2936]},
     {maskSplit_maskSelect_lo_2[2935:2932]},
     {maskSplit_maskSelect_lo_2[2931:2928]},
     {maskSplit_maskSelect_lo_2[2927:2924]},
     {maskSplit_maskSelect_lo_2[2923:2920]},
     {maskSplit_maskSelect_lo_2[2919:2916]},
     {maskSplit_maskSelect_lo_2[2915:2912]},
     {maskSplit_maskSelect_lo_2[2911:2908]},
     {maskSplit_maskSelect_lo_2[2907:2904]},
     {maskSplit_maskSelect_lo_2[2903:2900]},
     {maskSplit_maskSelect_lo_2[2899:2896]},
     {maskSplit_maskSelect_lo_2[2895:2892]},
     {maskSplit_maskSelect_lo_2[2891:2888]},
     {maskSplit_maskSelect_lo_2[2887:2884]},
     {maskSplit_maskSelect_lo_2[2883:2880]},
     {maskSplit_maskSelect_lo_2[2879:2876]},
     {maskSplit_maskSelect_lo_2[2875:2872]},
     {maskSplit_maskSelect_lo_2[2871:2868]},
     {maskSplit_maskSelect_lo_2[2867:2864]},
     {maskSplit_maskSelect_lo_2[2863:2860]},
     {maskSplit_maskSelect_lo_2[2859:2856]},
     {maskSplit_maskSelect_lo_2[2855:2852]},
     {maskSplit_maskSelect_lo_2[2851:2848]},
     {maskSplit_maskSelect_lo_2[2847:2844]},
     {maskSplit_maskSelect_lo_2[2843:2840]},
     {maskSplit_maskSelect_lo_2[2839:2836]},
     {maskSplit_maskSelect_lo_2[2835:2832]},
     {maskSplit_maskSelect_lo_2[2831:2828]},
     {maskSplit_maskSelect_lo_2[2827:2824]},
     {maskSplit_maskSelect_lo_2[2823:2820]},
     {maskSplit_maskSelect_lo_2[2819:2816]},
     {maskSplit_maskSelect_lo_2[2815:2812]},
     {maskSplit_maskSelect_lo_2[2811:2808]},
     {maskSplit_maskSelect_lo_2[2807:2804]},
     {maskSplit_maskSelect_lo_2[2803:2800]},
     {maskSplit_maskSelect_lo_2[2799:2796]},
     {maskSplit_maskSelect_lo_2[2795:2792]},
     {maskSplit_maskSelect_lo_2[2791:2788]},
     {maskSplit_maskSelect_lo_2[2787:2784]},
     {maskSplit_maskSelect_lo_2[2783:2780]},
     {maskSplit_maskSelect_lo_2[2779:2776]},
     {maskSplit_maskSelect_lo_2[2775:2772]},
     {maskSplit_maskSelect_lo_2[2771:2768]},
     {maskSplit_maskSelect_lo_2[2767:2764]},
     {maskSplit_maskSelect_lo_2[2763:2760]},
     {maskSplit_maskSelect_lo_2[2759:2756]},
     {maskSplit_maskSelect_lo_2[2755:2752]},
     {maskSplit_maskSelect_lo_2[2751:2748]},
     {maskSplit_maskSelect_lo_2[2747:2744]},
     {maskSplit_maskSelect_lo_2[2743:2740]},
     {maskSplit_maskSelect_lo_2[2739:2736]},
     {maskSplit_maskSelect_lo_2[2735:2732]},
     {maskSplit_maskSelect_lo_2[2731:2728]},
     {maskSplit_maskSelect_lo_2[2727:2724]},
     {maskSplit_maskSelect_lo_2[2723:2720]},
     {maskSplit_maskSelect_lo_2[2719:2716]},
     {maskSplit_maskSelect_lo_2[2715:2712]},
     {maskSplit_maskSelect_lo_2[2711:2708]},
     {maskSplit_maskSelect_lo_2[2707:2704]},
     {maskSplit_maskSelect_lo_2[2703:2700]},
     {maskSplit_maskSelect_lo_2[2699:2696]},
     {maskSplit_maskSelect_lo_2[2695:2692]},
     {maskSplit_maskSelect_lo_2[2691:2688]},
     {maskSplit_maskSelect_lo_2[2687:2684]},
     {maskSplit_maskSelect_lo_2[2683:2680]},
     {maskSplit_maskSelect_lo_2[2679:2676]},
     {maskSplit_maskSelect_lo_2[2675:2672]},
     {maskSplit_maskSelect_lo_2[2671:2668]},
     {maskSplit_maskSelect_lo_2[2667:2664]},
     {maskSplit_maskSelect_lo_2[2663:2660]},
     {maskSplit_maskSelect_lo_2[2659:2656]},
     {maskSplit_maskSelect_lo_2[2655:2652]},
     {maskSplit_maskSelect_lo_2[2651:2648]},
     {maskSplit_maskSelect_lo_2[2647:2644]},
     {maskSplit_maskSelect_lo_2[2643:2640]},
     {maskSplit_maskSelect_lo_2[2639:2636]},
     {maskSplit_maskSelect_lo_2[2635:2632]},
     {maskSplit_maskSelect_lo_2[2631:2628]},
     {maskSplit_maskSelect_lo_2[2627:2624]},
     {maskSplit_maskSelect_lo_2[2623:2620]},
     {maskSplit_maskSelect_lo_2[2619:2616]},
     {maskSplit_maskSelect_lo_2[2615:2612]},
     {maskSplit_maskSelect_lo_2[2611:2608]},
     {maskSplit_maskSelect_lo_2[2607:2604]},
     {maskSplit_maskSelect_lo_2[2603:2600]},
     {maskSplit_maskSelect_lo_2[2599:2596]},
     {maskSplit_maskSelect_lo_2[2595:2592]},
     {maskSplit_maskSelect_lo_2[2591:2588]},
     {maskSplit_maskSelect_lo_2[2587:2584]},
     {maskSplit_maskSelect_lo_2[2583:2580]},
     {maskSplit_maskSelect_lo_2[2579:2576]},
     {maskSplit_maskSelect_lo_2[2575:2572]},
     {maskSplit_maskSelect_lo_2[2571:2568]},
     {maskSplit_maskSelect_lo_2[2567:2564]},
     {maskSplit_maskSelect_lo_2[2563:2560]},
     {maskSplit_maskSelect_lo_2[2559:2556]},
     {maskSplit_maskSelect_lo_2[2555:2552]},
     {maskSplit_maskSelect_lo_2[2551:2548]},
     {maskSplit_maskSelect_lo_2[2547:2544]},
     {maskSplit_maskSelect_lo_2[2543:2540]},
     {maskSplit_maskSelect_lo_2[2539:2536]},
     {maskSplit_maskSelect_lo_2[2535:2532]},
     {maskSplit_maskSelect_lo_2[2531:2528]},
     {maskSplit_maskSelect_lo_2[2527:2524]},
     {maskSplit_maskSelect_lo_2[2523:2520]},
     {maskSplit_maskSelect_lo_2[2519:2516]},
     {maskSplit_maskSelect_lo_2[2515:2512]},
     {maskSplit_maskSelect_lo_2[2511:2508]},
     {maskSplit_maskSelect_lo_2[2507:2504]},
     {maskSplit_maskSelect_lo_2[2503:2500]},
     {maskSplit_maskSelect_lo_2[2499:2496]},
     {maskSplit_maskSelect_lo_2[2495:2492]},
     {maskSplit_maskSelect_lo_2[2491:2488]},
     {maskSplit_maskSelect_lo_2[2487:2484]},
     {maskSplit_maskSelect_lo_2[2483:2480]},
     {maskSplit_maskSelect_lo_2[2479:2476]},
     {maskSplit_maskSelect_lo_2[2475:2472]},
     {maskSplit_maskSelect_lo_2[2471:2468]},
     {maskSplit_maskSelect_lo_2[2467:2464]},
     {maskSplit_maskSelect_lo_2[2463:2460]},
     {maskSplit_maskSelect_lo_2[2459:2456]},
     {maskSplit_maskSelect_lo_2[2455:2452]},
     {maskSplit_maskSelect_lo_2[2451:2448]},
     {maskSplit_maskSelect_lo_2[2447:2444]},
     {maskSplit_maskSelect_lo_2[2443:2440]},
     {maskSplit_maskSelect_lo_2[2439:2436]},
     {maskSplit_maskSelect_lo_2[2435:2432]},
     {maskSplit_maskSelect_lo_2[2431:2428]},
     {maskSplit_maskSelect_lo_2[2427:2424]},
     {maskSplit_maskSelect_lo_2[2423:2420]},
     {maskSplit_maskSelect_lo_2[2419:2416]},
     {maskSplit_maskSelect_lo_2[2415:2412]},
     {maskSplit_maskSelect_lo_2[2411:2408]},
     {maskSplit_maskSelect_lo_2[2407:2404]},
     {maskSplit_maskSelect_lo_2[2403:2400]},
     {maskSplit_maskSelect_lo_2[2399:2396]},
     {maskSplit_maskSelect_lo_2[2395:2392]},
     {maskSplit_maskSelect_lo_2[2391:2388]},
     {maskSplit_maskSelect_lo_2[2387:2384]},
     {maskSplit_maskSelect_lo_2[2383:2380]},
     {maskSplit_maskSelect_lo_2[2379:2376]},
     {maskSplit_maskSelect_lo_2[2375:2372]},
     {maskSplit_maskSelect_lo_2[2371:2368]},
     {maskSplit_maskSelect_lo_2[2367:2364]},
     {maskSplit_maskSelect_lo_2[2363:2360]},
     {maskSplit_maskSelect_lo_2[2359:2356]},
     {maskSplit_maskSelect_lo_2[2355:2352]},
     {maskSplit_maskSelect_lo_2[2351:2348]},
     {maskSplit_maskSelect_lo_2[2347:2344]},
     {maskSplit_maskSelect_lo_2[2343:2340]},
     {maskSplit_maskSelect_lo_2[2339:2336]},
     {maskSplit_maskSelect_lo_2[2335:2332]},
     {maskSplit_maskSelect_lo_2[2331:2328]},
     {maskSplit_maskSelect_lo_2[2327:2324]},
     {maskSplit_maskSelect_lo_2[2323:2320]},
     {maskSplit_maskSelect_lo_2[2319:2316]},
     {maskSplit_maskSelect_lo_2[2315:2312]},
     {maskSplit_maskSelect_lo_2[2311:2308]},
     {maskSplit_maskSelect_lo_2[2307:2304]},
     {maskSplit_maskSelect_lo_2[2303:2300]},
     {maskSplit_maskSelect_lo_2[2299:2296]},
     {maskSplit_maskSelect_lo_2[2295:2292]},
     {maskSplit_maskSelect_lo_2[2291:2288]},
     {maskSplit_maskSelect_lo_2[2287:2284]},
     {maskSplit_maskSelect_lo_2[2283:2280]},
     {maskSplit_maskSelect_lo_2[2279:2276]},
     {maskSplit_maskSelect_lo_2[2275:2272]},
     {maskSplit_maskSelect_lo_2[2271:2268]},
     {maskSplit_maskSelect_lo_2[2267:2264]},
     {maskSplit_maskSelect_lo_2[2263:2260]},
     {maskSplit_maskSelect_lo_2[2259:2256]},
     {maskSplit_maskSelect_lo_2[2255:2252]},
     {maskSplit_maskSelect_lo_2[2251:2248]},
     {maskSplit_maskSelect_lo_2[2247:2244]},
     {maskSplit_maskSelect_lo_2[2243:2240]},
     {maskSplit_maskSelect_lo_2[2239:2236]},
     {maskSplit_maskSelect_lo_2[2235:2232]},
     {maskSplit_maskSelect_lo_2[2231:2228]},
     {maskSplit_maskSelect_lo_2[2227:2224]},
     {maskSplit_maskSelect_lo_2[2223:2220]},
     {maskSplit_maskSelect_lo_2[2219:2216]},
     {maskSplit_maskSelect_lo_2[2215:2212]},
     {maskSplit_maskSelect_lo_2[2211:2208]},
     {maskSplit_maskSelect_lo_2[2207:2204]},
     {maskSplit_maskSelect_lo_2[2203:2200]},
     {maskSplit_maskSelect_lo_2[2199:2196]},
     {maskSplit_maskSelect_lo_2[2195:2192]},
     {maskSplit_maskSelect_lo_2[2191:2188]},
     {maskSplit_maskSelect_lo_2[2187:2184]},
     {maskSplit_maskSelect_lo_2[2183:2180]},
     {maskSplit_maskSelect_lo_2[2179:2176]},
     {maskSplit_maskSelect_lo_2[2175:2172]},
     {maskSplit_maskSelect_lo_2[2171:2168]},
     {maskSplit_maskSelect_lo_2[2167:2164]},
     {maskSplit_maskSelect_lo_2[2163:2160]},
     {maskSplit_maskSelect_lo_2[2159:2156]},
     {maskSplit_maskSelect_lo_2[2155:2152]},
     {maskSplit_maskSelect_lo_2[2151:2148]},
     {maskSplit_maskSelect_lo_2[2147:2144]},
     {maskSplit_maskSelect_lo_2[2143:2140]},
     {maskSplit_maskSelect_lo_2[2139:2136]},
     {maskSplit_maskSelect_lo_2[2135:2132]},
     {maskSplit_maskSelect_lo_2[2131:2128]},
     {maskSplit_maskSelect_lo_2[2127:2124]},
     {maskSplit_maskSelect_lo_2[2123:2120]},
     {maskSplit_maskSelect_lo_2[2119:2116]},
     {maskSplit_maskSelect_lo_2[2115:2112]},
     {maskSplit_maskSelect_lo_2[2111:2108]},
     {maskSplit_maskSelect_lo_2[2107:2104]},
     {maskSplit_maskSelect_lo_2[2103:2100]},
     {maskSplit_maskSelect_lo_2[2099:2096]},
     {maskSplit_maskSelect_lo_2[2095:2092]},
     {maskSplit_maskSelect_lo_2[2091:2088]},
     {maskSplit_maskSelect_lo_2[2087:2084]},
     {maskSplit_maskSelect_lo_2[2083:2080]},
     {maskSplit_maskSelect_lo_2[2079:2076]},
     {maskSplit_maskSelect_lo_2[2075:2072]},
     {maskSplit_maskSelect_lo_2[2071:2068]},
     {maskSplit_maskSelect_lo_2[2067:2064]},
     {maskSplit_maskSelect_lo_2[2063:2060]},
     {maskSplit_maskSelect_lo_2[2059:2056]},
     {maskSplit_maskSelect_lo_2[2055:2052]},
     {maskSplit_maskSelect_lo_2[2051:2048]},
     {maskSplit_maskSelect_lo_2[2047:2044]},
     {maskSplit_maskSelect_lo_2[2043:2040]},
     {maskSplit_maskSelect_lo_2[2039:2036]},
     {maskSplit_maskSelect_lo_2[2035:2032]},
     {maskSplit_maskSelect_lo_2[2031:2028]},
     {maskSplit_maskSelect_lo_2[2027:2024]},
     {maskSplit_maskSelect_lo_2[2023:2020]},
     {maskSplit_maskSelect_lo_2[2019:2016]},
     {maskSplit_maskSelect_lo_2[2015:2012]},
     {maskSplit_maskSelect_lo_2[2011:2008]},
     {maskSplit_maskSelect_lo_2[2007:2004]},
     {maskSplit_maskSelect_lo_2[2003:2000]},
     {maskSplit_maskSelect_lo_2[1999:1996]},
     {maskSplit_maskSelect_lo_2[1995:1992]},
     {maskSplit_maskSelect_lo_2[1991:1988]},
     {maskSplit_maskSelect_lo_2[1987:1984]},
     {maskSplit_maskSelect_lo_2[1983:1980]},
     {maskSplit_maskSelect_lo_2[1979:1976]},
     {maskSplit_maskSelect_lo_2[1975:1972]},
     {maskSplit_maskSelect_lo_2[1971:1968]},
     {maskSplit_maskSelect_lo_2[1967:1964]},
     {maskSplit_maskSelect_lo_2[1963:1960]},
     {maskSplit_maskSelect_lo_2[1959:1956]},
     {maskSplit_maskSelect_lo_2[1955:1952]},
     {maskSplit_maskSelect_lo_2[1951:1948]},
     {maskSplit_maskSelect_lo_2[1947:1944]},
     {maskSplit_maskSelect_lo_2[1943:1940]},
     {maskSplit_maskSelect_lo_2[1939:1936]},
     {maskSplit_maskSelect_lo_2[1935:1932]},
     {maskSplit_maskSelect_lo_2[1931:1928]},
     {maskSplit_maskSelect_lo_2[1927:1924]},
     {maskSplit_maskSelect_lo_2[1923:1920]},
     {maskSplit_maskSelect_lo_2[1919:1916]},
     {maskSplit_maskSelect_lo_2[1915:1912]},
     {maskSplit_maskSelect_lo_2[1911:1908]},
     {maskSplit_maskSelect_lo_2[1907:1904]},
     {maskSplit_maskSelect_lo_2[1903:1900]},
     {maskSplit_maskSelect_lo_2[1899:1896]},
     {maskSplit_maskSelect_lo_2[1895:1892]},
     {maskSplit_maskSelect_lo_2[1891:1888]},
     {maskSplit_maskSelect_lo_2[1887:1884]},
     {maskSplit_maskSelect_lo_2[1883:1880]},
     {maskSplit_maskSelect_lo_2[1879:1876]},
     {maskSplit_maskSelect_lo_2[1875:1872]},
     {maskSplit_maskSelect_lo_2[1871:1868]},
     {maskSplit_maskSelect_lo_2[1867:1864]},
     {maskSplit_maskSelect_lo_2[1863:1860]},
     {maskSplit_maskSelect_lo_2[1859:1856]},
     {maskSplit_maskSelect_lo_2[1855:1852]},
     {maskSplit_maskSelect_lo_2[1851:1848]},
     {maskSplit_maskSelect_lo_2[1847:1844]},
     {maskSplit_maskSelect_lo_2[1843:1840]},
     {maskSplit_maskSelect_lo_2[1839:1836]},
     {maskSplit_maskSelect_lo_2[1835:1832]},
     {maskSplit_maskSelect_lo_2[1831:1828]},
     {maskSplit_maskSelect_lo_2[1827:1824]},
     {maskSplit_maskSelect_lo_2[1823:1820]},
     {maskSplit_maskSelect_lo_2[1819:1816]},
     {maskSplit_maskSelect_lo_2[1815:1812]},
     {maskSplit_maskSelect_lo_2[1811:1808]},
     {maskSplit_maskSelect_lo_2[1807:1804]},
     {maskSplit_maskSelect_lo_2[1803:1800]},
     {maskSplit_maskSelect_lo_2[1799:1796]},
     {maskSplit_maskSelect_lo_2[1795:1792]},
     {maskSplit_maskSelect_lo_2[1791:1788]},
     {maskSplit_maskSelect_lo_2[1787:1784]},
     {maskSplit_maskSelect_lo_2[1783:1780]},
     {maskSplit_maskSelect_lo_2[1779:1776]},
     {maskSplit_maskSelect_lo_2[1775:1772]},
     {maskSplit_maskSelect_lo_2[1771:1768]},
     {maskSplit_maskSelect_lo_2[1767:1764]},
     {maskSplit_maskSelect_lo_2[1763:1760]},
     {maskSplit_maskSelect_lo_2[1759:1756]},
     {maskSplit_maskSelect_lo_2[1755:1752]},
     {maskSplit_maskSelect_lo_2[1751:1748]},
     {maskSplit_maskSelect_lo_2[1747:1744]},
     {maskSplit_maskSelect_lo_2[1743:1740]},
     {maskSplit_maskSelect_lo_2[1739:1736]},
     {maskSplit_maskSelect_lo_2[1735:1732]},
     {maskSplit_maskSelect_lo_2[1731:1728]},
     {maskSplit_maskSelect_lo_2[1727:1724]},
     {maskSplit_maskSelect_lo_2[1723:1720]},
     {maskSplit_maskSelect_lo_2[1719:1716]},
     {maskSplit_maskSelect_lo_2[1715:1712]},
     {maskSplit_maskSelect_lo_2[1711:1708]},
     {maskSplit_maskSelect_lo_2[1707:1704]},
     {maskSplit_maskSelect_lo_2[1703:1700]},
     {maskSplit_maskSelect_lo_2[1699:1696]},
     {maskSplit_maskSelect_lo_2[1695:1692]},
     {maskSplit_maskSelect_lo_2[1691:1688]},
     {maskSplit_maskSelect_lo_2[1687:1684]},
     {maskSplit_maskSelect_lo_2[1683:1680]},
     {maskSplit_maskSelect_lo_2[1679:1676]},
     {maskSplit_maskSelect_lo_2[1675:1672]},
     {maskSplit_maskSelect_lo_2[1671:1668]},
     {maskSplit_maskSelect_lo_2[1667:1664]},
     {maskSplit_maskSelect_lo_2[1663:1660]},
     {maskSplit_maskSelect_lo_2[1659:1656]},
     {maskSplit_maskSelect_lo_2[1655:1652]},
     {maskSplit_maskSelect_lo_2[1651:1648]},
     {maskSplit_maskSelect_lo_2[1647:1644]},
     {maskSplit_maskSelect_lo_2[1643:1640]},
     {maskSplit_maskSelect_lo_2[1639:1636]},
     {maskSplit_maskSelect_lo_2[1635:1632]},
     {maskSplit_maskSelect_lo_2[1631:1628]},
     {maskSplit_maskSelect_lo_2[1627:1624]},
     {maskSplit_maskSelect_lo_2[1623:1620]},
     {maskSplit_maskSelect_lo_2[1619:1616]},
     {maskSplit_maskSelect_lo_2[1615:1612]},
     {maskSplit_maskSelect_lo_2[1611:1608]},
     {maskSplit_maskSelect_lo_2[1607:1604]},
     {maskSplit_maskSelect_lo_2[1603:1600]},
     {maskSplit_maskSelect_lo_2[1599:1596]},
     {maskSplit_maskSelect_lo_2[1595:1592]},
     {maskSplit_maskSelect_lo_2[1591:1588]},
     {maskSplit_maskSelect_lo_2[1587:1584]},
     {maskSplit_maskSelect_lo_2[1583:1580]},
     {maskSplit_maskSelect_lo_2[1579:1576]},
     {maskSplit_maskSelect_lo_2[1575:1572]},
     {maskSplit_maskSelect_lo_2[1571:1568]},
     {maskSplit_maskSelect_lo_2[1567:1564]},
     {maskSplit_maskSelect_lo_2[1563:1560]},
     {maskSplit_maskSelect_lo_2[1559:1556]},
     {maskSplit_maskSelect_lo_2[1555:1552]},
     {maskSplit_maskSelect_lo_2[1551:1548]},
     {maskSplit_maskSelect_lo_2[1547:1544]},
     {maskSplit_maskSelect_lo_2[1543:1540]},
     {maskSplit_maskSelect_lo_2[1539:1536]},
     {maskSplit_maskSelect_lo_2[1535:1532]},
     {maskSplit_maskSelect_lo_2[1531:1528]},
     {maskSplit_maskSelect_lo_2[1527:1524]},
     {maskSplit_maskSelect_lo_2[1523:1520]},
     {maskSplit_maskSelect_lo_2[1519:1516]},
     {maskSplit_maskSelect_lo_2[1515:1512]},
     {maskSplit_maskSelect_lo_2[1511:1508]},
     {maskSplit_maskSelect_lo_2[1507:1504]},
     {maskSplit_maskSelect_lo_2[1503:1500]},
     {maskSplit_maskSelect_lo_2[1499:1496]},
     {maskSplit_maskSelect_lo_2[1495:1492]},
     {maskSplit_maskSelect_lo_2[1491:1488]},
     {maskSplit_maskSelect_lo_2[1487:1484]},
     {maskSplit_maskSelect_lo_2[1483:1480]},
     {maskSplit_maskSelect_lo_2[1479:1476]},
     {maskSplit_maskSelect_lo_2[1475:1472]},
     {maskSplit_maskSelect_lo_2[1471:1468]},
     {maskSplit_maskSelect_lo_2[1467:1464]},
     {maskSplit_maskSelect_lo_2[1463:1460]},
     {maskSplit_maskSelect_lo_2[1459:1456]},
     {maskSplit_maskSelect_lo_2[1455:1452]},
     {maskSplit_maskSelect_lo_2[1451:1448]},
     {maskSplit_maskSelect_lo_2[1447:1444]},
     {maskSplit_maskSelect_lo_2[1443:1440]},
     {maskSplit_maskSelect_lo_2[1439:1436]},
     {maskSplit_maskSelect_lo_2[1435:1432]},
     {maskSplit_maskSelect_lo_2[1431:1428]},
     {maskSplit_maskSelect_lo_2[1427:1424]},
     {maskSplit_maskSelect_lo_2[1423:1420]},
     {maskSplit_maskSelect_lo_2[1419:1416]},
     {maskSplit_maskSelect_lo_2[1415:1412]},
     {maskSplit_maskSelect_lo_2[1411:1408]},
     {maskSplit_maskSelect_lo_2[1407:1404]},
     {maskSplit_maskSelect_lo_2[1403:1400]},
     {maskSplit_maskSelect_lo_2[1399:1396]},
     {maskSplit_maskSelect_lo_2[1395:1392]},
     {maskSplit_maskSelect_lo_2[1391:1388]},
     {maskSplit_maskSelect_lo_2[1387:1384]},
     {maskSplit_maskSelect_lo_2[1383:1380]},
     {maskSplit_maskSelect_lo_2[1379:1376]},
     {maskSplit_maskSelect_lo_2[1375:1372]},
     {maskSplit_maskSelect_lo_2[1371:1368]},
     {maskSplit_maskSelect_lo_2[1367:1364]},
     {maskSplit_maskSelect_lo_2[1363:1360]},
     {maskSplit_maskSelect_lo_2[1359:1356]},
     {maskSplit_maskSelect_lo_2[1355:1352]},
     {maskSplit_maskSelect_lo_2[1351:1348]},
     {maskSplit_maskSelect_lo_2[1347:1344]},
     {maskSplit_maskSelect_lo_2[1343:1340]},
     {maskSplit_maskSelect_lo_2[1339:1336]},
     {maskSplit_maskSelect_lo_2[1335:1332]},
     {maskSplit_maskSelect_lo_2[1331:1328]},
     {maskSplit_maskSelect_lo_2[1327:1324]},
     {maskSplit_maskSelect_lo_2[1323:1320]},
     {maskSplit_maskSelect_lo_2[1319:1316]},
     {maskSplit_maskSelect_lo_2[1315:1312]},
     {maskSplit_maskSelect_lo_2[1311:1308]},
     {maskSplit_maskSelect_lo_2[1307:1304]},
     {maskSplit_maskSelect_lo_2[1303:1300]},
     {maskSplit_maskSelect_lo_2[1299:1296]},
     {maskSplit_maskSelect_lo_2[1295:1292]},
     {maskSplit_maskSelect_lo_2[1291:1288]},
     {maskSplit_maskSelect_lo_2[1287:1284]},
     {maskSplit_maskSelect_lo_2[1283:1280]},
     {maskSplit_maskSelect_lo_2[1279:1276]},
     {maskSplit_maskSelect_lo_2[1275:1272]},
     {maskSplit_maskSelect_lo_2[1271:1268]},
     {maskSplit_maskSelect_lo_2[1267:1264]},
     {maskSplit_maskSelect_lo_2[1263:1260]},
     {maskSplit_maskSelect_lo_2[1259:1256]},
     {maskSplit_maskSelect_lo_2[1255:1252]},
     {maskSplit_maskSelect_lo_2[1251:1248]},
     {maskSplit_maskSelect_lo_2[1247:1244]},
     {maskSplit_maskSelect_lo_2[1243:1240]},
     {maskSplit_maskSelect_lo_2[1239:1236]},
     {maskSplit_maskSelect_lo_2[1235:1232]},
     {maskSplit_maskSelect_lo_2[1231:1228]},
     {maskSplit_maskSelect_lo_2[1227:1224]},
     {maskSplit_maskSelect_lo_2[1223:1220]},
     {maskSplit_maskSelect_lo_2[1219:1216]},
     {maskSplit_maskSelect_lo_2[1215:1212]},
     {maskSplit_maskSelect_lo_2[1211:1208]},
     {maskSplit_maskSelect_lo_2[1207:1204]},
     {maskSplit_maskSelect_lo_2[1203:1200]},
     {maskSplit_maskSelect_lo_2[1199:1196]},
     {maskSplit_maskSelect_lo_2[1195:1192]},
     {maskSplit_maskSelect_lo_2[1191:1188]},
     {maskSplit_maskSelect_lo_2[1187:1184]},
     {maskSplit_maskSelect_lo_2[1183:1180]},
     {maskSplit_maskSelect_lo_2[1179:1176]},
     {maskSplit_maskSelect_lo_2[1175:1172]},
     {maskSplit_maskSelect_lo_2[1171:1168]},
     {maskSplit_maskSelect_lo_2[1167:1164]},
     {maskSplit_maskSelect_lo_2[1163:1160]},
     {maskSplit_maskSelect_lo_2[1159:1156]},
     {maskSplit_maskSelect_lo_2[1155:1152]},
     {maskSplit_maskSelect_lo_2[1151:1148]},
     {maskSplit_maskSelect_lo_2[1147:1144]},
     {maskSplit_maskSelect_lo_2[1143:1140]},
     {maskSplit_maskSelect_lo_2[1139:1136]},
     {maskSplit_maskSelect_lo_2[1135:1132]},
     {maskSplit_maskSelect_lo_2[1131:1128]},
     {maskSplit_maskSelect_lo_2[1127:1124]},
     {maskSplit_maskSelect_lo_2[1123:1120]},
     {maskSplit_maskSelect_lo_2[1119:1116]},
     {maskSplit_maskSelect_lo_2[1115:1112]},
     {maskSplit_maskSelect_lo_2[1111:1108]},
     {maskSplit_maskSelect_lo_2[1107:1104]},
     {maskSplit_maskSelect_lo_2[1103:1100]},
     {maskSplit_maskSelect_lo_2[1099:1096]},
     {maskSplit_maskSelect_lo_2[1095:1092]},
     {maskSplit_maskSelect_lo_2[1091:1088]},
     {maskSplit_maskSelect_lo_2[1087:1084]},
     {maskSplit_maskSelect_lo_2[1083:1080]},
     {maskSplit_maskSelect_lo_2[1079:1076]},
     {maskSplit_maskSelect_lo_2[1075:1072]},
     {maskSplit_maskSelect_lo_2[1071:1068]},
     {maskSplit_maskSelect_lo_2[1067:1064]},
     {maskSplit_maskSelect_lo_2[1063:1060]},
     {maskSplit_maskSelect_lo_2[1059:1056]},
     {maskSplit_maskSelect_lo_2[1055:1052]},
     {maskSplit_maskSelect_lo_2[1051:1048]},
     {maskSplit_maskSelect_lo_2[1047:1044]},
     {maskSplit_maskSelect_lo_2[1043:1040]},
     {maskSplit_maskSelect_lo_2[1039:1036]},
     {maskSplit_maskSelect_lo_2[1035:1032]},
     {maskSplit_maskSelect_lo_2[1031:1028]},
     {maskSplit_maskSelect_lo_2[1027:1024]},
     {maskSplit_maskSelect_lo_2[1023:1020]},
     {maskSplit_maskSelect_lo_2[1019:1016]},
     {maskSplit_maskSelect_lo_2[1015:1012]},
     {maskSplit_maskSelect_lo_2[1011:1008]},
     {maskSplit_maskSelect_lo_2[1007:1004]},
     {maskSplit_maskSelect_lo_2[1003:1000]},
     {maskSplit_maskSelect_lo_2[999:996]},
     {maskSplit_maskSelect_lo_2[995:992]},
     {maskSplit_maskSelect_lo_2[991:988]},
     {maskSplit_maskSelect_lo_2[987:984]},
     {maskSplit_maskSelect_lo_2[983:980]},
     {maskSplit_maskSelect_lo_2[979:976]},
     {maskSplit_maskSelect_lo_2[975:972]},
     {maskSplit_maskSelect_lo_2[971:968]},
     {maskSplit_maskSelect_lo_2[967:964]},
     {maskSplit_maskSelect_lo_2[963:960]},
     {maskSplit_maskSelect_lo_2[959:956]},
     {maskSplit_maskSelect_lo_2[955:952]},
     {maskSplit_maskSelect_lo_2[951:948]},
     {maskSplit_maskSelect_lo_2[947:944]},
     {maskSplit_maskSelect_lo_2[943:940]},
     {maskSplit_maskSelect_lo_2[939:936]},
     {maskSplit_maskSelect_lo_2[935:932]},
     {maskSplit_maskSelect_lo_2[931:928]},
     {maskSplit_maskSelect_lo_2[927:924]},
     {maskSplit_maskSelect_lo_2[923:920]},
     {maskSplit_maskSelect_lo_2[919:916]},
     {maskSplit_maskSelect_lo_2[915:912]},
     {maskSplit_maskSelect_lo_2[911:908]},
     {maskSplit_maskSelect_lo_2[907:904]},
     {maskSplit_maskSelect_lo_2[903:900]},
     {maskSplit_maskSelect_lo_2[899:896]},
     {maskSplit_maskSelect_lo_2[895:892]},
     {maskSplit_maskSelect_lo_2[891:888]},
     {maskSplit_maskSelect_lo_2[887:884]},
     {maskSplit_maskSelect_lo_2[883:880]},
     {maskSplit_maskSelect_lo_2[879:876]},
     {maskSplit_maskSelect_lo_2[875:872]},
     {maskSplit_maskSelect_lo_2[871:868]},
     {maskSplit_maskSelect_lo_2[867:864]},
     {maskSplit_maskSelect_lo_2[863:860]},
     {maskSplit_maskSelect_lo_2[859:856]},
     {maskSplit_maskSelect_lo_2[855:852]},
     {maskSplit_maskSelect_lo_2[851:848]},
     {maskSplit_maskSelect_lo_2[847:844]},
     {maskSplit_maskSelect_lo_2[843:840]},
     {maskSplit_maskSelect_lo_2[839:836]},
     {maskSplit_maskSelect_lo_2[835:832]},
     {maskSplit_maskSelect_lo_2[831:828]},
     {maskSplit_maskSelect_lo_2[827:824]},
     {maskSplit_maskSelect_lo_2[823:820]},
     {maskSplit_maskSelect_lo_2[819:816]},
     {maskSplit_maskSelect_lo_2[815:812]},
     {maskSplit_maskSelect_lo_2[811:808]},
     {maskSplit_maskSelect_lo_2[807:804]},
     {maskSplit_maskSelect_lo_2[803:800]},
     {maskSplit_maskSelect_lo_2[799:796]},
     {maskSplit_maskSelect_lo_2[795:792]},
     {maskSplit_maskSelect_lo_2[791:788]},
     {maskSplit_maskSelect_lo_2[787:784]},
     {maskSplit_maskSelect_lo_2[783:780]},
     {maskSplit_maskSelect_lo_2[779:776]},
     {maskSplit_maskSelect_lo_2[775:772]},
     {maskSplit_maskSelect_lo_2[771:768]},
     {maskSplit_maskSelect_lo_2[767:764]},
     {maskSplit_maskSelect_lo_2[763:760]},
     {maskSplit_maskSelect_lo_2[759:756]},
     {maskSplit_maskSelect_lo_2[755:752]},
     {maskSplit_maskSelect_lo_2[751:748]},
     {maskSplit_maskSelect_lo_2[747:744]},
     {maskSplit_maskSelect_lo_2[743:740]},
     {maskSplit_maskSelect_lo_2[739:736]},
     {maskSplit_maskSelect_lo_2[735:732]},
     {maskSplit_maskSelect_lo_2[731:728]},
     {maskSplit_maskSelect_lo_2[727:724]},
     {maskSplit_maskSelect_lo_2[723:720]},
     {maskSplit_maskSelect_lo_2[719:716]},
     {maskSplit_maskSelect_lo_2[715:712]},
     {maskSplit_maskSelect_lo_2[711:708]},
     {maskSplit_maskSelect_lo_2[707:704]},
     {maskSplit_maskSelect_lo_2[703:700]},
     {maskSplit_maskSelect_lo_2[699:696]},
     {maskSplit_maskSelect_lo_2[695:692]},
     {maskSplit_maskSelect_lo_2[691:688]},
     {maskSplit_maskSelect_lo_2[687:684]},
     {maskSplit_maskSelect_lo_2[683:680]},
     {maskSplit_maskSelect_lo_2[679:676]},
     {maskSplit_maskSelect_lo_2[675:672]},
     {maskSplit_maskSelect_lo_2[671:668]},
     {maskSplit_maskSelect_lo_2[667:664]},
     {maskSplit_maskSelect_lo_2[663:660]},
     {maskSplit_maskSelect_lo_2[659:656]},
     {maskSplit_maskSelect_lo_2[655:652]},
     {maskSplit_maskSelect_lo_2[651:648]},
     {maskSplit_maskSelect_lo_2[647:644]},
     {maskSplit_maskSelect_lo_2[643:640]},
     {maskSplit_maskSelect_lo_2[639:636]},
     {maskSplit_maskSelect_lo_2[635:632]},
     {maskSplit_maskSelect_lo_2[631:628]},
     {maskSplit_maskSelect_lo_2[627:624]},
     {maskSplit_maskSelect_lo_2[623:620]},
     {maskSplit_maskSelect_lo_2[619:616]},
     {maskSplit_maskSelect_lo_2[615:612]},
     {maskSplit_maskSelect_lo_2[611:608]},
     {maskSplit_maskSelect_lo_2[607:604]},
     {maskSplit_maskSelect_lo_2[603:600]},
     {maskSplit_maskSelect_lo_2[599:596]},
     {maskSplit_maskSelect_lo_2[595:592]},
     {maskSplit_maskSelect_lo_2[591:588]},
     {maskSplit_maskSelect_lo_2[587:584]},
     {maskSplit_maskSelect_lo_2[583:580]},
     {maskSplit_maskSelect_lo_2[579:576]},
     {maskSplit_maskSelect_lo_2[575:572]},
     {maskSplit_maskSelect_lo_2[571:568]},
     {maskSplit_maskSelect_lo_2[567:564]},
     {maskSplit_maskSelect_lo_2[563:560]},
     {maskSplit_maskSelect_lo_2[559:556]},
     {maskSplit_maskSelect_lo_2[555:552]},
     {maskSplit_maskSelect_lo_2[551:548]},
     {maskSplit_maskSelect_lo_2[547:544]},
     {maskSplit_maskSelect_lo_2[543:540]},
     {maskSplit_maskSelect_lo_2[539:536]},
     {maskSplit_maskSelect_lo_2[535:532]},
     {maskSplit_maskSelect_lo_2[531:528]},
     {maskSplit_maskSelect_lo_2[527:524]},
     {maskSplit_maskSelect_lo_2[523:520]},
     {maskSplit_maskSelect_lo_2[519:516]},
     {maskSplit_maskSelect_lo_2[515:512]},
     {maskSplit_maskSelect_lo_2[511:508]},
     {maskSplit_maskSelect_lo_2[507:504]},
     {maskSplit_maskSelect_lo_2[503:500]},
     {maskSplit_maskSelect_lo_2[499:496]},
     {maskSplit_maskSelect_lo_2[495:492]},
     {maskSplit_maskSelect_lo_2[491:488]},
     {maskSplit_maskSelect_lo_2[487:484]},
     {maskSplit_maskSelect_lo_2[483:480]},
     {maskSplit_maskSelect_lo_2[479:476]},
     {maskSplit_maskSelect_lo_2[475:472]},
     {maskSplit_maskSelect_lo_2[471:468]},
     {maskSplit_maskSelect_lo_2[467:464]},
     {maskSplit_maskSelect_lo_2[463:460]},
     {maskSplit_maskSelect_lo_2[459:456]},
     {maskSplit_maskSelect_lo_2[455:452]},
     {maskSplit_maskSelect_lo_2[451:448]},
     {maskSplit_maskSelect_lo_2[447:444]},
     {maskSplit_maskSelect_lo_2[443:440]},
     {maskSplit_maskSelect_lo_2[439:436]},
     {maskSplit_maskSelect_lo_2[435:432]},
     {maskSplit_maskSelect_lo_2[431:428]},
     {maskSplit_maskSelect_lo_2[427:424]},
     {maskSplit_maskSelect_lo_2[423:420]},
     {maskSplit_maskSelect_lo_2[419:416]},
     {maskSplit_maskSelect_lo_2[415:412]},
     {maskSplit_maskSelect_lo_2[411:408]},
     {maskSplit_maskSelect_lo_2[407:404]},
     {maskSplit_maskSelect_lo_2[403:400]},
     {maskSplit_maskSelect_lo_2[399:396]},
     {maskSplit_maskSelect_lo_2[395:392]},
     {maskSplit_maskSelect_lo_2[391:388]},
     {maskSplit_maskSelect_lo_2[387:384]},
     {maskSplit_maskSelect_lo_2[383:380]},
     {maskSplit_maskSelect_lo_2[379:376]},
     {maskSplit_maskSelect_lo_2[375:372]},
     {maskSplit_maskSelect_lo_2[371:368]},
     {maskSplit_maskSelect_lo_2[367:364]},
     {maskSplit_maskSelect_lo_2[363:360]},
     {maskSplit_maskSelect_lo_2[359:356]},
     {maskSplit_maskSelect_lo_2[355:352]},
     {maskSplit_maskSelect_lo_2[351:348]},
     {maskSplit_maskSelect_lo_2[347:344]},
     {maskSplit_maskSelect_lo_2[343:340]},
     {maskSplit_maskSelect_lo_2[339:336]},
     {maskSplit_maskSelect_lo_2[335:332]},
     {maskSplit_maskSelect_lo_2[331:328]},
     {maskSplit_maskSelect_lo_2[327:324]},
     {maskSplit_maskSelect_lo_2[323:320]},
     {maskSplit_maskSelect_lo_2[319:316]},
     {maskSplit_maskSelect_lo_2[315:312]},
     {maskSplit_maskSelect_lo_2[311:308]},
     {maskSplit_maskSelect_lo_2[307:304]},
     {maskSplit_maskSelect_lo_2[303:300]},
     {maskSplit_maskSelect_lo_2[299:296]},
     {maskSplit_maskSelect_lo_2[295:292]},
     {maskSplit_maskSelect_lo_2[291:288]},
     {maskSplit_maskSelect_lo_2[287:284]},
     {maskSplit_maskSelect_lo_2[283:280]},
     {maskSplit_maskSelect_lo_2[279:276]},
     {maskSplit_maskSelect_lo_2[275:272]},
     {maskSplit_maskSelect_lo_2[271:268]},
     {maskSplit_maskSelect_lo_2[267:264]},
     {maskSplit_maskSelect_lo_2[263:260]},
     {maskSplit_maskSelect_lo_2[259:256]},
     {maskSplit_maskSelect_lo_2[255:252]},
     {maskSplit_maskSelect_lo_2[251:248]},
     {maskSplit_maskSelect_lo_2[247:244]},
     {maskSplit_maskSelect_lo_2[243:240]},
     {maskSplit_maskSelect_lo_2[239:236]},
     {maskSplit_maskSelect_lo_2[235:232]},
     {maskSplit_maskSelect_lo_2[231:228]},
     {maskSplit_maskSelect_lo_2[227:224]},
     {maskSplit_maskSelect_lo_2[223:220]},
     {maskSplit_maskSelect_lo_2[219:216]},
     {maskSplit_maskSelect_lo_2[215:212]},
     {maskSplit_maskSelect_lo_2[211:208]},
     {maskSplit_maskSelect_lo_2[207:204]},
     {maskSplit_maskSelect_lo_2[203:200]},
     {maskSplit_maskSelect_lo_2[199:196]},
     {maskSplit_maskSelect_lo_2[195:192]},
     {maskSplit_maskSelect_lo_2[191:188]},
     {maskSplit_maskSelect_lo_2[187:184]},
     {maskSplit_maskSelect_lo_2[183:180]},
     {maskSplit_maskSelect_lo_2[179:176]},
     {maskSplit_maskSelect_lo_2[175:172]},
     {maskSplit_maskSelect_lo_2[171:168]},
     {maskSplit_maskSelect_lo_2[167:164]},
     {maskSplit_maskSelect_lo_2[163:160]},
     {maskSplit_maskSelect_lo_2[159:156]},
     {maskSplit_maskSelect_lo_2[155:152]},
     {maskSplit_maskSelect_lo_2[151:148]},
     {maskSplit_maskSelect_lo_2[147:144]},
     {maskSplit_maskSelect_lo_2[143:140]},
     {maskSplit_maskSelect_lo_2[139:136]},
     {maskSplit_maskSelect_lo_2[135:132]},
     {maskSplit_maskSelect_lo_2[131:128]},
     {maskSplit_maskSelect_lo_2[127:124]},
     {maskSplit_maskSelect_lo_2[123:120]},
     {maskSplit_maskSelect_lo_2[119:116]},
     {maskSplit_maskSelect_lo_2[115:112]},
     {maskSplit_maskSelect_lo_2[111:108]},
     {maskSplit_maskSelect_lo_2[107:104]},
     {maskSplit_maskSelect_lo_2[103:100]},
     {maskSplit_maskSelect_lo_2[99:96]},
     {maskSplit_maskSelect_lo_2[95:92]},
     {maskSplit_maskSelect_lo_2[91:88]},
     {maskSplit_maskSelect_lo_2[87:84]},
     {maskSplit_maskSelect_lo_2[83:80]},
     {maskSplit_maskSelect_lo_2[79:76]},
     {maskSplit_maskSelect_lo_2[75:72]},
     {maskSplit_maskSelect_lo_2[71:68]},
     {maskSplit_maskSelect_lo_2[67:64]},
     {maskSplit_maskSelect_lo_2[63:60]},
     {maskSplit_maskSelect_lo_2[59:56]},
     {maskSplit_maskSelect_lo_2[55:52]},
     {maskSplit_maskSelect_lo_2[51:48]},
     {maskSplit_maskSelect_lo_2[47:44]},
     {maskSplit_maskSelect_lo_2[43:40]},
     {maskSplit_maskSelect_lo_2[39:36]},
     {maskSplit_maskSelect_lo_2[35:32]},
     {maskSplit_maskSelect_lo_2[31:28]},
     {maskSplit_maskSelect_lo_2[27:24]},
     {maskSplit_maskSelect_lo_2[23:20]},
     {maskSplit_maskSelect_lo_2[19:16]},
     {maskSplit_maskSelect_lo_2[15:12]},
     {maskSplit_maskSelect_lo_2[11:8]},
     {maskSplit_maskSelect_lo_2[7:4]},
     {maskSplit_maskSelect_lo_2[3:0]}};
  wire [3:0]         maskSplit_2_2 = (instReg_maskType ? _GEN_147[executeGroupCounter] : 4'hF) & maskSplit_vlBoundaryCorrection_2;
  wire [7:0]         maskSplit_byteMask_lo_2 = {{4{maskSplit_2_2[1]}}, {4{maskSplit_2_2[0]}}};
  wire [7:0]         maskSplit_byteMask_hi_2 = {{4{maskSplit_2_2[3]}}, {4{maskSplit_2_2[2]}}};
  wire [15:0]        maskSplit_2_1 = {maskSplit_byteMask_hi_2, maskSplit_byteMask_lo_2};
  wire [15:0]        executeByteMask = (sew1H[0] ? maskSplit_0_1 : 16'h0) | (sew1H[1] ? maskSplit_1_1 : 16'h0) | (sew1H[2] ? maskSplit_2_1 : 16'h0);
  wire [15:0]        _executeElementMask_T_3 = sew1H[0] ? maskSplit_0_2 : 16'h0;
  wire [7:0]         _GEN_148 = _executeElementMask_T_3[7:0] | (sew1H[1] ? maskSplit_1_2 : 8'h0);
  wire [15:0]        executeElementMask = {_executeElementMask_T_3[15:8], _GEN_148[7:4], _GEN_148[3:0] | (sew1H[2] ? maskSplit_2_2 : 4'h0)};
  wire [127:0]       maskForDestination_lo_lo_lo_lo_lo_lo = {maskForDestination_lo_lo_lo_lo_lo_lo_hi, maskForDestination_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]       maskForDestination_lo_lo_lo_lo_lo_hi = {maskForDestination_lo_lo_lo_lo_lo_hi_hi, maskForDestination_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]       maskForDestination_lo_lo_lo_lo_lo = {maskForDestination_lo_lo_lo_lo_lo_hi, maskForDestination_lo_lo_lo_lo_lo_lo};
  wire [127:0]       maskForDestination_lo_lo_lo_lo_hi_lo = {maskForDestination_lo_lo_lo_lo_hi_lo_hi, maskForDestination_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]       maskForDestination_lo_lo_lo_lo_hi_hi = {maskForDestination_lo_lo_lo_lo_hi_hi_hi, maskForDestination_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]       maskForDestination_lo_lo_lo_lo_hi = {maskForDestination_lo_lo_lo_lo_hi_hi, maskForDestination_lo_lo_lo_lo_hi_lo};
  wire [511:0]       maskForDestination_lo_lo_lo_lo = {maskForDestination_lo_lo_lo_lo_hi, maskForDestination_lo_lo_lo_lo_lo};
  wire [127:0]       maskForDestination_lo_lo_lo_hi_lo_lo = {maskForDestination_lo_lo_lo_hi_lo_lo_hi, maskForDestination_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]       maskForDestination_lo_lo_lo_hi_lo_hi = {maskForDestination_lo_lo_lo_hi_lo_hi_hi, maskForDestination_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]       maskForDestination_lo_lo_lo_hi_lo = {maskForDestination_lo_lo_lo_hi_lo_hi, maskForDestination_lo_lo_lo_hi_lo_lo};
  wire [127:0]       maskForDestination_lo_lo_lo_hi_hi_lo = {maskForDestination_lo_lo_lo_hi_hi_lo_hi, maskForDestination_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]       maskForDestination_lo_lo_lo_hi_hi_hi = {maskForDestination_lo_lo_lo_hi_hi_hi_hi, maskForDestination_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]       maskForDestination_lo_lo_lo_hi_hi = {maskForDestination_lo_lo_lo_hi_hi_hi, maskForDestination_lo_lo_lo_hi_hi_lo};
  wire [511:0]       maskForDestination_lo_lo_lo_hi = {maskForDestination_lo_lo_lo_hi_hi, maskForDestination_lo_lo_lo_hi_lo};
  wire [1023:0]      maskForDestination_lo_lo_lo = {maskForDestination_lo_lo_lo_hi, maskForDestination_lo_lo_lo_lo};
  wire [127:0]       maskForDestination_lo_lo_hi_lo_lo_lo = {maskForDestination_lo_lo_hi_lo_lo_lo_hi, maskForDestination_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]       maskForDestination_lo_lo_hi_lo_lo_hi = {maskForDestination_lo_lo_hi_lo_lo_hi_hi, maskForDestination_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]       maskForDestination_lo_lo_hi_lo_lo = {maskForDestination_lo_lo_hi_lo_lo_hi, maskForDestination_lo_lo_hi_lo_lo_lo};
  wire [127:0]       maskForDestination_lo_lo_hi_lo_hi_lo = {maskForDestination_lo_lo_hi_lo_hi_lo_hi, maskForDestination_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]       maskForDestination_lo_lo_hi_lo_hi_hi = {maskForDestination_lo_lo_hi_lo_hi_hi_hi, maskForDestination_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]       maskForDestination_lo_lo_hi_lo_hi = {maskForDestination_lo_lo_hi_lo_hi_hi, maskForDestination_lo_lo_hi_lo_hi_lo};
  wire [511:0]       maskForDestination_lo_lo_hi_lo = {maskForDestination_lo_lo_hi_lo_hi, maskForDestination_lo_lo_hi_lo_lo};
  wire [127:0]       maskForDestination_lo_lo_hi_hi_lo_lo = {maskForDestination_lo_lo_hi_hi_lo_lo_hi, maskForDestination_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]       maskForDestination_lo_lo_hi_hi_lo_hi = {maskForDestination_lo_lo_hi_hi_lo_hi_hi, maskForDestination_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]       maskForDestination_lo_lo_hi_hi_lo = {maskForDestination_lo_lo_hi_hi_lo_hi, maskForDestination_lo_lo_hi_hi_lo_lo};
  wire [127:0]       maskForDestination_lo_lo_hi_hi_hi_lo = {maskForDestination_lo_lo_hi_hi_hi_lo_hi, maskForDestination_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]       maskForDestination_lo_lo_hi_hi_hi_hi = {maskForDestination_lo_lo_hi_hi_hi_hi_hi, maskForDestination_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]       maskForDestination_lo_lo_hi_hi_hi = {maskForDestination_lo_lo_hi_hi_hi_hi, maskForDestination_lo_lo_hi_hi_hi_lo};
  wire [511:0]       maskForDestination_lo_lo_hi_hi = {maskForDestination_lo_lo_hi_hi_hi, maskForDestination_lo_lo_hi_hi_lo};
  wire [1023:0]      maskForDestination_lo_lo_hi = {maskForDestination_lo_lo_hi_hi, maskForDestination_lo_lo_hi_lo};
  wire [2047:0]      maskForDestination_lo_lo = {maskForDestination_lo_lo_hi, maskForDestination_lo_lo_lo};
  wire [127:0]       maskForDestination_lo_hi_lo_lo_lo_lo = {maskForDestination_lo_hi_lo_lo_lo_lo_hi, maskForDestination_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]       maskForDestination_lo_hi_lo_lo_lo_hi = {maskForDestination_lo_hi_lo_lo_lo_hi_hi, maskForDestination_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]       maskForDestination_lo_hi_lo_lo_lo = {maskForDestination_lo_hi_lo_lo_lo_hi, maskForDestination_lo_hi_lo_lo_lo_lo};
  wire [127:0]       maskForDestination_lo_hi_lo_lo_hi_lo = {maskForDestination_lo_hi_lo_lo_hi_lo_hi, maskForDestination_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]       maskForDestination_lo_hi_lo_lo_hi_hi = {maskForDestination_lo_hi_lo_lo_hi_hi_hi, maskForDestination_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]       maskForDestination_lo_hi_lo_lo_hi = {maskForDestination_lo_hi_lo_lo_hi_hi, maskForDestination_lo_hi_lo_lo_hi_lo};
  wire [511:0]       maskForDestination_lo_hi_lo_lo = {maskForDestination_lo_hi_lo_lo_hi, maskForDestination_lo_hi_lo_lo_lo};
  wire [127:0]       maskForDestination_lo_hi_lo_hi_lo_lo = {maskForDestination_lo_hi_lo_hi_lo_lo_hi, maskForDestination_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]       maskForDestination_lo_hi_lo_hi_lo_hi = {maskForDestination_lo_hi_lo_hi_lo_hi_hi, maskForDestination_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]       maskForDestination_lo_hi_lo_hi_lo = {maskForDestination_lo_hi_lo_hi_lo_hi, maskForDestination_lo_hi_lo_hi_lo_lo};
  wire [127:0]       maskForDestination_lo_hi_lo_hi_hi_lo = {maskForDestination_lo_hi_lo_hi_hi_lo_hi, maskForDestination_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]       maskForDestination_lo_hi_lo_hi_hi_hi = {maskForDestination_lo_hi_lo_hi_hi_hi_hi, maskForDestination_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]       maskForDestination_lo_hi_lo_hi_hi = {maskForDestination_lo_hi_lo_hi_hi_hi, maskForDestination_lo_hi_lo_hi_hi_lo};
  wire [511:0]       maskForDestination_lo_hi_lo_hi = {maskForDestination_lo_hi_lo_hi_hi, maskForDestination_lo_hi_lo_hi_lo};
  wire [1023:0]      maskForDestination_lo_hi_lo = {maskForDestination_lo_hi_lo_hi, maskForDestination_lo_hi_lo_lo};
  wire [127:0]       maskForDestination_lo_hi_hi_lo_lo_lo = {maskForDestination_lo_hi_hi_lo_lo_lo_hi, maskForDestination_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]       maskForDestination_lo_hi_hi_lo_lo_hi = {maskForDestination_lo_hi_hi_lo_lo_hi_hi, maskForDestination_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]       maskForDestination_lo_hi_hi_lo_lo = {maskForDestination_lo_hi_hi_lo_lo_hi, maskForDestination_lo_hi_hi_lo_lo_lo};
  wire [127:0]       maskForDestination_lo_hi_hi_lo_hi_lo = {maskForDestination_lo_hi_hi_lo_hi_lo_hi, maskForDestination_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]       maskForDestination_lo_hi_hi_lo_hi_hi = {maskForDestination_lo_hi_hi_lo_hi_hi_hi, maskForDestination_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]       maskForDestination_lo_hi_hi_lo_hi = {maskForDestination_lo_hi_hi_lo_hi_hi, maskForDestination_lo_hi_hi_lo_hi_lo};
  wire [511:0]       maskForDestination_lo_hi_hi_lo = {maskForDestination_lo_hi_hi_lo_hi, maskForDestination_lo_hi_hi_lo_lo};
  wire [127:0]       maskForDestination_lo_hi_hi_hi_lo_lo = {maskForDestination_lo_hi_hi_hi_lo_lo_hi, maskForDestination_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]       maskForDestination_lo_hi_hi_hi_lo_hi = {maskForDestination_lo_hi_hi_hi_lo_hi_hi, maskForDestination_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]       maskForDestination_lo_hi_hi_hi_lo = {maskForDestination_lo_hi_hi_hi_lo_hi, maskForDestination_lo_hi_hi_hi_lo_lo};
  wire [127:0]       maskForDestination_lo_hi_hi_hi_hi_lo = {maskForDestination_lo_hi_hi_hi_hi_lo_hi, maskForDestination_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]       maskForDestination_lo_hi_hi_hi_hi_hi = {maskForDestination_lo_hi_hi_hi_hi_hi_hi, maskForDestination_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]       maskForDestination_lo_hi_hi_hi_hi = {maskForDestination_lo_hi_hi_hi_hi_hi, maskForDestination_lo_hi_hi_hi_hi_lo};
  wire [511:0]       maskForDestination_lo_hi_hi_hi = {maskForDestination_lo_hi_hi_hi_hi, maskForDestination_lo_hi_hi_hi_lo};
  wire [1023:0]      maskForDestination_lo_hi_hi = {maskForDestination_lo_hi_hi_hi, maskForDestination_lo_hi_hi_lo};
  wire [2047:0]      maskForDestination_lo_hi = {maskForDestination_lo_hi_hi, maskForDestination_lo_hi_lo};
  wire [4095:0]      maskForDestination_lo = {maskForDestination_lo_hi, maskForDestination_lo_lo};
  wire [127:0]       maskForDestination_hi_lo_lo_lo_lo_lo = {maskForDestination_hi_lo_lo_lo_lo_lo_hi, maskForDestination_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]       maskForDestination_hi_lo_lo_lo_lo_hi = {maskForDestination_hi_lo_lo_lo_lo_hi_hi, maskForDestination_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]       maskForDestination_hi_lo_lo_lo_lo = {maskForDestination_hi_lo_lo_lo_lo_hi, maskForDestination_hi_lo_lo_lo_lo_lo};
  wire [127:0]       maskForDestination_hi_lo_lo_lo_hi_lo = {maskForDestination_hi_lo_lo_lo_hi_lo_hi, maskForDestination_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]       maskForDestination_hi_lo_lo_lo_hi_hi = {maskForDestination_hi_lo_lo_lo_hi_hi_hi, maskForDestination_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]       maskForDestination_hi_lo_lo_lo_hi = {maskForDestination_hi_lo_lo_lo_hi_hi, maskForDestination_hi_lo_lo_lo_hi_lo};
  wire [511:0]       maskForDestination_hi_lo_lo_lo = {maskForDestination_hi_lo_lo_lo_hi, maskForDestination_hi_lo_lo_lo_lo};
  wire [127:0]       maskForDestination_hi_lo_lo_hi_lo_lo = {maskForDestination_hi_lo_lo_hi_lo_lo_hi, maskForDestination_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]       maskForDestination_hi_lo_lo_hi_lo_hi = {maskForDestination_hi_lo_lo_hi_lo_hi_hi, maskForDestination_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]       maskForDestination_hi_lo_lo_hi_lo = {maskForDestination_hi_lo_lo_hi_lo_hi, maskForDestination_hi_lo_lo_hi_lo_lo};
  wire [127:0]       maskForDestination_hi_lo_lo_hi_hi_lo = {maskForDestination_hi_lo_lo_hi_hi_lo_hi, maskForDestination_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]       maskForDestination_hi_lo_lo_hi_hi_hi = {maskForDestination_hi_lo_lo_hi_hi_hi_hi, maskForDestination_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]       maskForDestination_hi_lo_lo_hi_hi = {maskForDestination_hi_lo_lo_hi_hi_hi, maskForDestination_hi_lo_lo_hi_hi_lo};
  wire [511:0]       maskForDestination_hi_lo_lo_hi = {maskForDestination_hi_lo_lo_hi_hi, maskForDestination_hi_lo_lo_hi_lo};
  wire [1023:0]      maskForDestination_hi_lo_lo = {maskForDestination_hi_lo_lo_hi, maskForDestination_hi_lo_lo_lo};
  wire [127:0]       maskForDestination_hi_lo_hi_lo_lo_lo = {maskForDestination_hi_lo_hi_lo_lo_lo_hi, maskForDestination_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]       maskForDestination_hi_lo_hi_lo_lo_hi = {maskForDestination_hi_lo_hi_lo_lo_hi_hi, maskForDestination_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]       maskForDestination_hi_lo_hi_lo_lo = {maskForDestination_hi_lo_hi_lo_lo_hi, maskForDestination_hi_lo_hi_lo_lo_lo};
  wire [127:0]       maskForDestination_hi_lo_hi_lo_hi_lo = {maskForDestination_hi_lo_hi_lo_hi_lo_hi, maskForDestination_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]       maskForDestination_hi_lo_hi_lo_hi_hi = {maskForDestination_hi_lo_hi_lo_hi_hi_hi, maskForDestination_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]       maskForDestination_hi_lo_hi_lo_hi = {maskForDestination_hi_lo_hi_lo_hi_hi, maskForDestination_hi_lo_hi_lo_hi_lo};
  wire [511:0]       maskForDestination_hi_lo_hi_lo = {maskForDestination_hi_lo_hi_lo_hi, maskForDestination_hi_lo_hi_lo_lo};
  wire [127:0]       maskForDestination_hi_lo_hi_hi_lo_lo = {maskForDestination_hi_lo_hi_hi_lo_lo_hi, maskForDestination_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]       maskForDestination_hi_lo_hi_hi_lo_hi = {maskForDestination_hi_lo_hi_hi_lo_hi_hi, maskForDestination_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]       maskForDestination_hi_lo_hi_hi_lo = {maskForDestination_hi_lo_hi_hi_lo_hi, maskForDestination_hi_lo_hi_hi_lo_lo};
  wire [127:0]       maskForDestination_hi_lo_hi_hi_hi_lo = {maskForDestination_hi_lo_hi_hi_hi_lo_hi, maskForDestination_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]       maskForDestination_hi_lo_hi_hi_hi_hi = {maskForDestination_hi_lo_hi_hi_hi_hi_hi, maskForDestination_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]       maskForDestination_hi_lo_hi_hi_hi = {maskForDestination_hi_lo_hi_hi_hi_hi, maskForDestination_hi_lo_hi_hi_hi_lo};
  wire [511:0]       maskForDestination_hi_lo_hi_hi = {maskForDestination_hi_lo_hi_hi_hi, maskForDestination_hi_lo_hi_hi_lo};
  wire [1023:0]      maskForDestination_hi_lo_hi = {maskForDestination_hi_lo_hi_hi, maskForDestination_hi_lo_hi_lo};
  wire [2047:0]      maskForDestination_hi_lo = {maskForDestination_hi_lo_hi, maskForDestination_hi_lo_lo};
  wire [127:0]       maskForDestination_hi_hi_lo_lo_lo_lo = {maskForDestination_hi_hi_lo_lo_lo_lo_hi, maskForDestination_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]       maskForDestination_hi_hi_lo_lo_lo_hi = {maskForDestination_hi_hi_lo_lo_lo_hi_hi, maskForDestination_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]       maskForDestination_hi_hi_lo_lo_lo = {maskForDestination_hi_hi_lo_lo_lo_hi, maskForDestination_hi_hi_lo_lo_lo_lo};
  wire [127:0]       maskForDestination_hi_hi_lo_lo_hi_lo = {maskForDestination_hi_hi_lo_lo_hi_lo_hi, maskForDestination_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]       maskForDestination_hi_hi_lo_lo_hi_hi = {maskForDestination_hi_hi_lo_lo_hi_hi_hi, maskForDestination_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]       maskForDestination_hi_hi_lo_lo_hi = {maskForDestination_hi_hi_lo_lo_hi_hi, maskForDestination_hi_hi_lo_lo_hi_lo};
  wire [511:0]       maskForDestination_hi_hi_lo_lo = {maskForDestination_hi_hi_lo_lo_hi, maskForDestination_hi_hi_lo_lo_lo};
  wire [127:0]       maskForDestination_hi_hi_lo_hi_lo_lo = {maskForDestination_hi_hi_lo_hi_lo_lo_hi, maskForDestination_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]       maskForDestination_hi_hi_lo_hi_lo_hi = {maskForDestination_hi_hi_lo_hi_lo_hi_hi, maskForDestination_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]       maskForDestination_hi_hi_lo_hi_lo = {maskForDestination_hi_hi_lo_hi_lo_hi, maskForDestination_hi_hi_lo_hi_lo_lo};
  wire [127:0]       maskForDestination_hi_hi_lo_hi_hi_lo = {maskForDestination_hi_hi_lo_hi_hi_lo_hi, maskForDestination_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]       maskForDestination_hi_hi_lo_hi_hi_hi = {maskForDestination_hi_hi_lo_hi_hi_hi_hi, maskForDestination_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]       maskForDestination_hi_hi_lo_hi_hi = {maskForDestination_hi_hi_lo_hi_hi_hi, maskForDestination_hi_hi_lo_hi_hi_lo};
  wire [511:0]       maskForDestination_hi_hi_lo_hi = {maskForDestination_hi_hi_lo_hi_hi, maskForDestination_hi_hi_lo_hi_lo};
  wire [1023:0]      maskForDestination_hi_hi_lo = {maskForDestination_hi_hi_lo_hi, maskForDestination_hi_hi_lo_lo};
  wire [127:0]       maskForDestination_hi_hi_hi_lo_lo_lo = {maskForDestination_hi_hi_hi_lo_lo_lo_hi, maskForDestination_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]       maskForDestination_hi_hi_hi_lo_lo_hi = {maskForDestination_hi_hi_hi_lo_lo_hi_hi, maskForDestination_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]       maskForDestination_hi_hi_hi_lo_lo = {maskForDestination_hi_hi_hi_lo_lo_hi, maskForDestination_hi_hi_hi_lo_lo_lo};
  wire [127:0]       maskForDestination_hi_hi_hi_lo_hi_lo = {maskForDestination_hi_hi_hi_lo_hi_lo_hi, maskForDestination_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]       maskForDestination_hi_hi_hi_lo_hi_hi = {maskForDestination_hi_hi_hi_lo_hi_hi_hi, maskForDestination_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]       maskForDestination_hi_hi_hi_lo_hi = {maskForDestination_hi_hi_hi_lo_hi_hi, maskForDestination_hi_hi_hi_lo_hi_lo};
  wire [511:0]       maskForDestination_hi_hi_hi_lo = {maskForDestination_hi_hi_hi_lo_hi, maskForDestination_hi_hi_hi_lo_lo};
  wire [127:0]       maskForDestination_hi_hi_hi_hi_lo_lo = {maskForDestination_hi_hi_hi_hi_lo_lo_hi, maskForDestination_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]       maskForDestination_hi_hi_hi_hi_lo_hi = {maskForDestination_hi_hi_hi_hi_lo_hi_hi, maskForDestination_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]       maskForDestination_hi_hi_hi_hi_lo = {maskForDestination_hi_hi_hi_hi_lo_hi, maskForDestination_hi_hi_hi_hi_lo_lo};
  wire [127:0]       maskForDestination_hi_hi_hi_hi_hi_lo = {maskForDestination_hi_hi_hi_hi_hi_lo_hi, maskForDestination_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]       maskForDestination_hi_hi_hi_hi_hi_hi = {maskForDestination_hi_hi_hi_hi_hi_hi_hi, maskForDestination_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]       maskForDestination_hi_hi_hi_hi_hi = {maskForDestination_hi_hi_hi_hi_hi_hi, maskForDestination_hi_hi_hi_hi_hi_lo};
  wire [511:0]       maskForDestination_hi_hi_hi_hi = {maskForDestination_hi_hi_hi_hi_hi, maskForDestination_hi_hi_hi_hi_lo};
  wire [1023:0]      maskForDestination_hi_hi_hi = {maskForDestination_hi_hi_hi_hi, maskForDestination_hi_hi_hi_lo};
  wire [2047:0]      maskForDestination_hi_hi = {maskForDestination_hi_hi_hi, maskForDestination_hi_hi_lo};
  wire [4095:0]      maskForDestination_hi = {maskForDestination_hi_hi, maskForDestination_hi_lo};
  wire [127:0]       _lastGroupMask_T = 128'h1 << elementTailForMaskDestination;
  wire [126:0]       _GEN_149 = _lastGroupMask_T[126:0] | _lastGroupMask_T[127:1];
  wire [125:0]       _GEN_150 = _GEN_149[125:0] | {_lastGroupMask_T[127], _GEN_149[126:2]};
  wire [123:0]       _GEN_151 = _GEN_150[123:0] | {_lastGroupMask_T[127], _GEN_149[126], _GEN_150[125:4]};
  wire [119:0]       _GEN_152 = _GEN_151[119:0] | {_lastGroupMask_T[127], _GEN_149[126], _GEN_150[125:124], _GEN_151[123:8]};
  wire [111:0]       _GEN_153 = _GEN_152[111:0] | {_lastGroupMask_T[127], _GEN_149[126], _GEN_150[125:124], _GEN_151[123:120], _GEN_152[119:16]};
  wire [95:0]        _GEN_154 = _GEN_153[95:0] | {_lastGroupMask_T[127], _GEN_149[126], _GEN_150[125:124], _GEN_151[123:120], _GEN_152[119:112], _GEN_153[111:32]};
  wire [127:0]       lastGroupMask =
    {_lastGroupMask_T[127],
     _GEN_149[126],
     _GEN_150[125:124],
     _GEN_151[123:120],
     _GEN_152[119:112],
     _GEN_153[111:96],
     _GEN_154[95:64],
     _GEN_154[63:0] | {_lastGroupMask_T[127], _GEN_149[126], _GEN_150[125:124], _GEN_151[123:120], _GEN_152[119:112], _GEN_153[111:96], _GEN_154[95:64]}};
  wire [63:0][127:0] _GEN_155 =
    {{maskForDestination_hi[4095:3968]},
     {maskForDestination_hi[3967:3840]},
     {maskForDestination_hi[3839:3712]},
     {maskForDestination_hi[3711:3584]},
     {maskForDestination_hi[3583:3456]},
     {maskForDestination_hi[3455:3328]},
     {maskForDestination_hi[3327:3200]},
     {maskForDestination_hi[3199:3072]},
     {maskForDestination_hi[3071:2944]},
     {maskForDestination_hi[2943:2816]},
     {maskForDestination_hi[2815:2688]},
     {maskForDestination_hi[2687:2560]},
     {maskForDestination_hi[2559:2432]},
     {maskForDestination_hi[2431:2304]},
     {maskForDestination_hi[2303:2176]},
     {maskForDestination_hi[2175:2048]},
     {maskForDestination_hi[2047:1920]},
     {maskForDestination_hi[1919:1792]},
     {maskForDestination_hi[1791:1664]},
     {maskForDestination_hi[1663:1536]},
     {maskForDestination_hi[1535:1408]},
     {maskForDestination_hi[1407:1280]},
     {maskForDestination_hi[1279:1152]},
     {maskForDestination_hi[1151:1024]},
     {maskForDestination_hi[1023:896]},
     {maskForDestination_hi[895:768]},
     {maskForDestination_hi[767:640]},
     {maskForDestination_hi[639:512]},
     {maskForDestination_hi[511:384]},
     {maskForDestination_hi[383:256]},
     {maskForDestination_hi[255:128]},
     {maskForDestination_hi[127:0]},
     {maskForDestination_lo[4095:3968]},
     {maskForDestination_lo[3967:3840]},
     {maskForDestination_lo[3839:3712]},
     {maskForDestination_lo[3711:3584]},
     {maskForDestination_lo[3583:3456]},
     {maskForDestination_lo[3455:3328]},
     {maskForDestination_lo[3327:3200]},
     {maskForDestination_lo[3199:3072]},
     {maskForDestination_lo[3071:2944]},
     {maskForDestination_lo[2943:2816]},
     {maskForDestination_lo[2815:2688]},
     {maskForDestination_lo[2687:2560]},
     {maskForDestination_lo[2559:2432]},
     {maskForDestination_lo[2431:2304]},
     {maskForDestination_lo[2303:2176]},
     {maskForDestination_lo[2175:2048]},
     {maskForDestination_lo[2047:1920]},
     {maskForDestination_lo[1919:1792]},
     {maskForDestination_lo[1791:1664]},
     {maskForDestination_lo[1663:1536]},
     {maskForDestination_lo[1535:1408]},
     {maskForDestination_lo[1407:1280]},
     {maskForDestination_lo[1279:1152]},
     {maskForDestination_lo[1151:1024]},
     {maskForDestination_lo[1023:896]},
     {maskForDestination_lo[895:768]},
     {maskForDestination_lo[767:640]},
     {maskForDestination_lo[639:512]},
     {maskForDestination_lo[511:384]},
     {maskForDestination_lo[383:256]},
     {maskForDestination_lo[255:128]},
     {maskForDestination_lo[127:0]}};
  wire [127:0]       currentMaskGroupForDestination =
    (lastGroup ? lastGroupMask : 128'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF) & (instReg_maskType & ~instReg_decodeResult_maskSource ? _GEN_155[requestCounter[5:0]] : 128'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF);
  wire [63:0]        _GEN_156 = {exeReqReg_1_bits_source1, exeReqReg_0_bits_source1};
  wire [63:0]        groupSourceData_lo;
  assign groupSourceData_lo = _GEN_156;
  wire [63:0]        source1_lo;
  assign source1_lo = _GEN_156;
  wire [63:0]        _GEN_157 = {exeReqReg_3_bits_source1, exeReqReg_2_bits_source1};
  wire [63:0]        groupSourceData_hi;
  assign groupSourceData_hi = _GEN_157;
  wire [63:0]        source1_hi;
  assign source1_hi = _GEN_157;
  wire [127:0]       groupSourceData = {groupSourceData_hi, groupSourceData_lo};
  wire [1:0]         _GEN_158 = {exeReqReg_1_valid, exeReqReg_0_valid};
  wire [1:0]         groupSourceValid_lo;
  assign groupSourceValid_lo = _GEN_158;
  wire [1:0]         view__in_bits_validInput_lo;
  assign view__in_bits_validInput_lo = _GEN_158;
  wire [1:0]         view__in_bits_sourceValid_lo;
  assign view__in_bits_sourceValid_lo = _GEN_158;
  wire [1:0]         _GEN_159 = {exeReqReg_3_valid, exeReqReg_2_valid};
  wire [1:0]         groupSourceValid_hi;
  assign groupSourceValid_hi = _GEN_159;
  wire [1:0]         view__in_bits_validInput_hi;
  assign view__in_bits_validInput_hi = _GEN_159;
  wire [1:0]         view__in_bits_sourceValid_hi;
  assign view__in_bits_sourceValid_hi = _GEN_159;
  wire [3:0]         groupSourceValid = {groupSourceValid_hi, groupSourceValid_lo};
  wire [1:0]         shifterSize = (sourceDataEEW1H[0] ? executeIndex : 2'h0) | (sourceDataEEW1H[1] ? {executeIndex[1], 1'h0} : 2'h0);
  wire [3:0]         _shifterSource_T = 4'h1 << shifterSize;
  wire [127:0]       _shifterSource_T_8 = _shifterSource_T[0] ? groupSourceData : 128'h0;
  wire [95:0]        _GEN_160 = _shifterSource_T_8[95:0] | (_shifterSource_T[1] ? groupSourceData[127:32] : 96'h0);
  wire [63:0]        _GEN_161 = _GEN_160[63:0] | (_shifterSource_T[2] ? groupSourceData[127:64] : 64'h0);
  wire [127:0]       shifterSource = {_shifterSource_T_8[127:96], _GEN_160[95:64], _GEN_161[63:32], _GEN_161[31:0] | (_shifterSource_T[3] ? groupSourceData[127:96] : 32'h0)};
  wire [7:0]         selectValid_lo = {{4{groupSourceValid[1]}}, {4{groupSourceValid[0]}}};
  wire [7:0]         selectValid_hi = {{4{groupSourceValid[3]}}, {4{groupSourceValid[2]}}};
  wire [3:0]         selectValid_lo_1 = {{2{groupSourceValid[1]}}, {2{groupSourceValid[0]}}};
  wire [3:0]         selectValid_hi_1 = {{2{groupSourceValid[3]}}, {2{groupSourceValid[2]}}};
  wire [3:0][3:0]    _GEN_162 = {{selectValid_hi[7:4]}, {selectValid_hi[3:0]}, {selectValid_lo[7:4]}, {selectValid_lo[3:0]}};
  wire [3:0]         selectValid = (sourceDataEEW1H[0] ? _GEN_162[executeIndex] : 4'h0) | (sourceDataEEW1H[1] ? (executeIndex[1] ? selectValid_hi_1 : selectValid_lo_1) : 4'h0) | (sourceDataEEW1H[2] ? groupSourceValid : 4'h0);
  wire [31:0]        source_0 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[7:0] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[15:0] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[31:0] : 32'h0);
  wire [31:0]        source_1 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[15:8] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[31:16] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[63:32] : 32'h0);
  wire [31:0]        source_2 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[23:16] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[47:32] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[95:64] : 32'h0);
  wire [31:0]        source_3 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[31:24] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[63:48] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[127:96] : 32'h0);
  wire [3:0]         _GEN_163 = selectValid & readMaskCorrection;
  wire [3:0]         checkVec_validVec;
  assign checkVec_validVec = _GEN_163;
  wire [3:0]         checkVec_validVec_1;
  assign checkVec_validVec_1 = _GEN_163;
  wire [3:0]         checkVec_validVec_2;
  assign checkVec_validVec_2 = _GEN_163;
  wire               checkVec_checkResultVec_0_6 = checkVec_validVec[0];
  wire [3:0]         _GEN_164 = 4'h1 << instReg_vlmul[1:0];
  wire [3:0]         checkVec_checkResultVec_intLMULInput;
  assign checkVec_checkResultVec_intLMULInput = _GEN_164;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_1;
  assign checkVec_checkResultVec_intLMULInput_1 = _GEN_164;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_2;
  assign checkVec_checkResultVec_intLMULInput_2 = _GEN_164;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_3;
  assign checkVec_checkResultVec_intLMULInput_3 = _GEN_164;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_4;
  assign checkVec_checkResultVec_intLMULInput_4 = _GEN_164;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_5;
  assign checkVec_checkResultVec_intLMULInput_5 = _GEN_164;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_6;
  assign checkVec_checkResultVec_intLMULInput_6 = _GEN_164;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_7;
  assign checkVec_checkResultVec_intLMULInput_7 = _GEN_164;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_8;
  assign checkVec_checkResultVec_intLMULInput_8 = _GEN_164;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_9;
  assign checkVec_checkResultVec_intLMULInput_9 = _GEN_164;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_10;
  assign checkVec_checkResultVec_intLMULInput_10 = _GEN_164;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_11;
  assign checkVec_checkResultVec_intLMULInput_11 = _GEN_164;
  wire [12:0]        checkVec_checkResultVec_dataPosition = source_0[12:0];
  wire [3:0]         checkVec_checkResultVec_0_0 = 4'h1 << checkVec_checkResultVec_dataPosition[1:0];
  wire [1:0]         checkVec_checkResultVec_0_1 = checkVec_checkResultVec_dataPosition[1:0];
  wire [1:0]         checkVec_checkResultVec_0_2 = checkVec_checkResultVec_dataPosition[3:2];
  wire [8:0]         checkVec_checkResultVec_dataGroup = checkVec_checkResultVec_dataPosition[12:4];
  wire [5:0]         checkVec_checkResultVec_0_3 = checkVec_checkResultVec_dataGroup[5:0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth = checkVec_checkResultVec_dataGroup[8:6];
  wire [2:0]         checkVec_checkResultVec_0_4 = checkVec_checkResultVec_accessRegGrowth;
  wire [7:0]         checkVec_checkResultVec_decimalProportion = {checkVec_checkResultVec_0_3, checkVec_checkResultVec_0_2};
  wire [2:0]         checkVec_checkResultVec_decimal = checkVec_checkResultVec_decimalProportion[7:5];
  wire               checkVec_checkResultVec_overlap =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal >= checkVec_checkResultVec_intLMULInput[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth} >= checkVec_checkResultVec_intLMULInput, source_0[31:13]};
  wire               checkVec_checkResultVec_0_5 = checkVec_checkResultVec_overlap | ~checkVec_checkResultVec_0_6;
  wire               checkVec_checkResultVec_1_6 = checkVec_validVec[1];
  wire [12:0]        checkVec_checkResultVec_dataPosition_1 = source_1[12:0];
  wire [3:0]         checkVec_checkResultVec_1_0 = 4'h1 << checkVec_checkResultVec_dataPosition_1[1:0];
  wire [1:0]         checkVec_checkResultVec_1_1 = checkVec_checkResultVec_dataPosition_1[1:0];
  wire [1:0]         checkVec_checkResultVec_1_2 = checkVec_checkResultVec_dataPosition_1[3:2];
  wire [8:0]         checkVec_checkResultVec_dataGroup_1 = checkVec_checkResultVec_dataPosition_1[12:4];
  wire [5:0]         checkVec_checkResultVec_1_3 = checkVec_checkResultVec_dataGroup_1[5:0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_1 = checkVec_checkResultVec_dataGroup_1[8:6];
  wire [2:0]         checkVec_checkResultVec_1_4 = checkVec_checkResultVec_accessRegGrowth_1;
  wire [7:0]         checkVec_checkResultVec_decimalProportion_1 = {checkVec_checkResultVec_1_3, checkVec_checkResultVec_1_2};
  wire [2:0]         checkVec_checkResultVec_decimal_1 = checkVec_checkResultVec_decimalProportion_1[7:5];
  wire               checkVec_checkResultVec_overlap_1 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_1 >= checkVec_checkResultVec_intLMULInput_1[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_1} >= checkVec_checkResultVec_intLMULInput_1, source_1[31:13]};
  wire               checkVec_checkResultVec_1_5 = checkVec_checkResultVec_overlap_1 | ~checkVec_checkResultVec_1_6;
  wire               checkVec_checkResultVec_2_6 = checkVec_validVec[2];
  wire [12:0]        checkVec_checkResultVec_dataPosition_2 = source_2[12:0];
  wire [3:0]         checkVec_checkResultVec_2_0 = 4'h1 << checkVec_checkResultVec_dataPosition_2[1:0];
  wire [1:0]         checkVec_checkResultVec_2_1 = checkVec_checkResultVec_dataPosition_2[1:0];
  wire [1:0]         checkVec_checkResultVec_2_2 = checkVec_checkResultVec_dataPosition_2[3:2];
  wire [8:0]         checkVec_checkResultVec_dataGroup_2 = checkVec_checkResultVec_dataPosition_2[12:4];
  wire [5:0]         checkVec_checkResultVec_2_3 = checkVec_checkResultVec_dataGroup_2[5:0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_2 = checkVec_checkResultVec_dataGroup_2[8:6];
  wire [2:0]         checkVec_checkResultVec_2_4 = checkVec_checkResultVec_accessRegGrowth_2;
  wire [7:0]         checkVec_checkResultVec_decimalProportion_2 = {checkVec_checkResultVec_2_3, checkVec_checkResultVec_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_2 = checkVec_checkResultVec_decimalProportion_2[7:5];
  wire               checkVec_checkResultVec_overlap_2 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_2 >= checkVec_checkResultVec_intLMULInput_2[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_2} >= checkVec_checkResultVec_intLMULInput_2, source_2[31:13]};
  wire               checkVec_checkResultVec_2_5 = checkVec_checkResultVec_overlap_2 | ~checkVec_checkResultVec_2_6;
  wire               checkVec_checkResultVec_3_6 = checkVec_validVec[3];
  wire [12:0]        checkVec_checkResultVec_dataPosition_3 = source_3[12:0];
  wire [3:0]         checkVec_checkResultVec_3_0 = 4'h1 << checkVec_checkResultVec_dataPosition_3[1:0];
  wire [1:0]         checkVec_checkResultVec_3_1 = checkVec_checkResultVec_dataPosition_3[1:0];
  wire [1:0]         checkVec_checkResultVec_3_2 = checkVec_checkResultVec_dataPosition_3[3:2];
  wire [8:0]         checkVec_checkResultVec_dataGroup_3 = checkVec_checkResultVec_dataPosition_3[12:4];
  wire [5:0]         checkVec_checkResultVec_3_3 = checkVec_checkResultVec_dataGroup_3[5:0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_3 = checkVec_checkResultVec_dataGroup_3[8:6];
  wire [2:0]         checkVec_checkResultVec_3_4 = checkVec_checkResultVec_accessRegGrowth_3;
  wire [7:0]         checkVec_checkResultVec_decimalProportion_3 = {checkVec_checkResultVec_3_3, checkVec_checkResultVec_3_2};
  wire [2:0]         checkVec_checkResultVec_decimal_3 = checkVec_checkResultVec_decimalProportion_3[7:5];
  wire               checkVec_checkResultVec_overlap_3 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_3 >= checkVec_checkResultVec_intLMULInput_3[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_3} >= checkVec_checkResultVec_intLMULInput_3, source_3[31:13]};
  wire               checkVec_checkResultVec_3_5 = checkVec_checkResultVec_overlap_3 | ~checkVec_checkResultVec_3_6;
  wire [7:0]         checkVec_checkResult_lo = {checkVec_checkResultVec_1_0, checkVec_checkResultVec_0_0};
  wire [7:0]         checkVec_checkResult_hi = {checkVec_checkResultVec_3_0, checkVec_checkResultVec_2_0};
  wire [15:0]        checkVec_0_0 = {checkVec_checkResult_hi, checkVec_checkResult_lo};
  wire [3:0]         checkVec_checkResult_lo_1 = {checkVec_checkResultVec_1_1, checkVec_checkResultVec_0_1};
  wire [3:0]         checkVec_checkResult_hi_1 = {checkVec_checkResultVec_3_1, checkVec_checkResultVec_2_1};
  wire [7:0]         checkVec_0_1 = {checkVec_checkResult_hi_1, checkVec_checkResult_lo_1};
  wire [3:0]         checkVec_checkResult_lo_2 = {checkVec_checkResultVec_1_2, checkVec_checkResultVec_0_2};
  wire [3:0]         checkVec_checkResult_hi_2 = {checkVec_checkResultVec_3_2, checkVec_checkResultVec_2_2};
  wire [7:0]         checkVec_0_2 = {checkVec_checkResult_hi_2, checkVec_checkResult_lo_2};
  wire [11:0]        checkVec_checkResult_lo_3 = {checkVec_checkResultVec_1_3, checkVec_checkResultVec_0_3};
  wire [11:0]        checkVec_checkResult_hi_3 = {checkVec_checkResultVec_3_3, checkVec_checkResultVec_2_3};
  wire [23:0]        checkVec_0_3 = {checkVec_checkResult_hi_3, checkVec_checkResult_lo_3};
  wire [5:0]         checkVec_checkResult_lo_4 = {checkVec_checkResultVec_1_4, checkVec_checkResultVec_0_4};
  wire [5:0]         checkVec_checkResult_hi_4 = {checkVec_checkResultVec_3_4, checkVec_checkResultVec_2_4};
  wire [11:0]        checkVec_0_4 = {checkVec_checkResult_hi_4, checkVec_checkResult_lo_4};
  wire [1:0]         checkVec_checkResult_lo_5 = {checkVec_checkResultVec_1_5, checkVec_checkResultVec_0_5};
  wire [1:0]         checkVec_checkResult_hi_5 = {checkVec_checkResultVec_3_5, checkVec_checkResultVec_2_5};
  wire [3:0]         checkVec_0_5 = {checkVec_checkResult_hi_5, checkVec_checkResult_lo_5};
  wire [1:0]         checkVec_checkResult_lo_6 = {checkVec_checkResultVec_1_6, checkVec_checkResultVec_0_6};
  wire [1:0]         checkVec_checkResult_hi_6 = {checkVec_checkResultVec_3_6, checkVec_checkResultVec_2_6};
  wire [3:0]         checkVec_0_6 = {checkVec_checkResult_hi_6, checkVec_checkResult_lo_6};
  wire               checkVec_checkResultVec_0_6_1 = checkVec_validVec_1[0];
  wire [12:0]        checkVec_checkResultVec_dataPosition_4 = {source_0[11:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_35 = 2'h1 << checkVec_checkResultVec_dataPosition_4[1];
  wire [3:0]         checkVec_checkResultVec_0_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_35[1]}}, {2{_checkVec_checkResultVec_accessMask_T_35[0]}}};
  wire [1:0]         checkVec_checkResultVec_0_1_1 = {checkVec_checkResultVec_dataPosition_4[1], 1'h0};
  wire [1:0]         checkVec_checkResultVec_0_2_1 = checkVec_checkResultVec_dataPosition_4[3:2];
  wire [8:0]         checkVec_checkResultVec_dataGroup_4 = checkVec_checkResultVec_dataPosition_4[12:4];
  wire [5:0]         checkVec_checkResultVec_0_3_1 = checkVec_checkResultVec_dataGroup_4[5:0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_4 = checkVec_checkResultVec_dataGroup_4[8:6];
  wire [2:0]         checkVec_checkResultVec_0_4_1 = checkVec_checkResultVec_accessRegGrowth_4;
  wire [7:0]         checkVec_checkResultVec_decimalProportion_4 = {checkVec_checkResultVec_0_3_1, checkVec_checkResultVec_0_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_4 = checkVec_checkResultVec_decimalProportion_4[7:5];
  wire               checkVec_checkResultVec_overlap_4 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_4 >= checkVec_checkResultVec_intLMULInput_4[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_4} >= checkVec_checkResultVec_intLMULInput_4, source_0[31:13]};
  wire               checkVec_checkResultVec_0_5_1 = checkVec_checkResultVec_overlap_4 | ~checkVec_checkResultVec_0_6_1;
  wire               checkVec_checkResultVec_1_6_1 = checkVec_validVec_1[1];
  wire [12:0]        checkVec_checkResultVec_dataPosition_5 = {source_1[11:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_43 = 2'h1 << checkVec_checkResultVec_dataPosition_5[1];
  wire [3:0]         checkVec_checkResultVec_1_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_43[1]}}, {2{_checkVec_checkResultVec_accessMask_T_43[0]}}};
  wire [1:0]         checkVec_checkResultVec_1_1_1 = {checkVec_checkResultVec_dataPosition_5[1], 1'h0};
  wire [1:0]         checkVec_checkResultVec_1_2_1 = checkVec_checkResultVec_dataPosition_5[3:2];
  wire [8:0]         checkVec_checkResultVec_dataGroup_5 = checkVec_checkResultVec_dataPosition_5[12:4];
  wire [5:0]         checkVec_checkResultVec_1_3_1 = checkVec_checkResultVec_dataGroup_5[5:0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_5 = checkVec_checkResultVec_dataGroup_5[8:6];
  wire [2:0]         checkVec_checkResultVec_1_4_1 = checkVec_checkResultVec_accessRegGrowth_5;
  wire [7:0]         checkVec_checkResultVec_decimalProportion_5 = {checkVec_checkResultVec_1_3_1, checkVec_checkResultVec_1_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_5 = checkVec_checkResultVec_decimalProportion_5[7:5];
  wire               checkVec_checkResultVec_overlap_5 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_5 >= checkVec_checkResultVec_intLMULInput_5[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_5} >= checkVec_checkResultVec_intLMULInput_5, source_1[31:13]};
  wire               checkVec_checkResultVec_1_5_1 = checkVec_checkResultVec_overlap_5 | ~checkVec_checkResultVec_1_6_1;
  wire               checkVec_checkResultVec_2_6_1 = checkVec_validVec_1[2];
  wire [12:0]        checkVec_checkResultVec_dataPosition_6 = {source_2[11:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_51 = 2'h1 << checkVec_checkResultVec_dataPosition_6[1];
  wire [3:0]         checkVec_checkResultVec_2_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_51[1]}}, {2{_checkVec_checkResultVec_accessMask_T_51[0]}}};
  wire [1:0]         checkVec_checkResultVec_2_1_1 = {checkVec_checkResultVec_dataPosition_6[1], 1'h0};
  wire [1:0]         checkVec_checkResultVec_2_2_1 = checkVec_checkResultVec_dataPosition_6[3:2];
  wire [8:0]         checkVec_checkResultVec_dataGroup_6 = checkVec_checkResultVec_dataPosition_6[12:4];
  wire [5:0]         checkVec_checkResultVec_2_3_1 = checkVec_checkResultVec_dataGroup_6[5:0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_6 = checkVec_checkResultVec_dataGroup_6[8:6];
  wire [2:0]         checkVec_checkResultVec_2_4_1 = checkVec_checkResultVec_accessRegGrowth_6;
  wire [7:0]         checkVec_checkResultVec_decimalProportion_6 = {checkVec_checkResultVec_2_3_1, checkVec_checkResultVec_2_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_6 = checkVec_checkResultVec_decimalProportion_6[7:5];
  wire               checkVec_checkResultVec_overlap_6 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_6 >= checkVec_checkResultVec_intLMULInput_6[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_6} >= checkVec_checkResultVec_intLMULInput_6, source_2[31:13]};
  wire               checkVec_checkResultVec_2_5_1 = checkVec_checkResultVec_overlap_6 | ~checkVec_checkResultVec_2_6_1;
  wire               checkVec_checkResultVec_3_6_1 = checkVec_validVec_1[3];
  wire [12:0]        checkVec_checkResultVec_dataPosition_7 = {source_3[11:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_59 = 2'h1 << checkVec_checkResultVec_dataPosition_7[1];
  wire [3:0]         checkVec_checkResultVec_3_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_59[1]}}, {2{_checkVec_checkResultVec_accessMask_T_59[0]}}};
  wire [1:0]         checkVec_checkResultVec_3_1_1 = {checkVec_checkResultVec_dataPosition_7[1], 1'h0};
  wire [1:0]         checkVec_checkResultVec_3_2_1 = checkVec_checkResultVec_dataPosition_7[3:2];
  wire [8:0]         checkVec_checkResultVec_dataGroup_7 = checkVec_checkResultVec_dataPosition_7[12:4];
  wire [5:0]         checkVec_checkResultVec_3_3_1 = checkVec_checkResultVec_dataGroup_7[5:0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_7 = checkVec_checkResultVec_dataGroup_7[8:6];
  wire [2:0]         checkVec_checkResultVec_3_4_1 = checkVec_checkResultVec_accessRegGrowth_7;
  wire [7:0]         checkVec_checkResultVec_decimalProportion_7 = {checkVec_checkResultVec_3_3_1, checkVec_checkResultVec_3_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_7 = checkVec_checkResultVec_decimalProportion_7[7:5];
  wire               checkVec_checkResultVec_overlap_7 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_7 >= checkVec_checkResultVec_intLMULInput_7[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_7} >= checkVec_checkResultVec_intLMULInput_7, source_3[31:13]};
  wire               checkVec_checkResultVec_3_5_1 = checkVec_checkResultVec_overlap_7 | ~checkVec_checkResultVec_3_6_1;
  wire [7:0]         checkVec_checkResult_lo_7 = {checkVec_checkResultVec_1_0_1, checkVec_checkResultVec_0_0_1};
  wire [7:0]         checkVec_checkResult_hi_7 = {checkVec_checkResultVec_3_0_1, checkVec_checkResultVec_2_0_1};
  wire [15:0]        checkVec_1_0 = {checkVec_checkResult_hi_7, checkVec_checkResult_lo_7};
  wire [3:0]         checkVec_checkResult_lo_8 = {checkVec_checkResultVec_1_1_1, checkVec_checkResultVec_0_1_1};
  wire [3:0]         checkVec_checkResult_hi_8 = {checkVec_checkResultVec_3_1_1, checkVec_checkResultVec_2_1_1};
  wire [7:0]         checkVec_1_1 = {checkVec_checkResult_hi_8, checkVec_checkResult_lo_8};
  wire [3:0]         checkVec_checkResult_lo_9 = {checkVec_checkResultVec_1_2_1, checkVec_checkResultVec_0_2_1};
  wire [3:0]         checkVec_checkResult_hi_9 = {checkVec_checkResultVec_3_2_1, checkVec_checkResultVec_2_2_1};
  wire [7:0]         checkVec_1_2 = {checkVec_checkResult_hi_9, checkVec_checkResult_lo_9};
  wire [11:0]        checkVec_checkResult_lo_10 = {checkVec_checkResultVec_1_3_1, checkVec_checkResultVec_0_3_1};
  wire [11:0]        checkVec_checkResult_hi_10 = {checkVec_checkResultVec_3_3_1, checkVec_checkResultVec_2_3_1};
  wire [23:0]        checkVec_1_3 = {checkVec_checkResult_hi_10, checkVec_checkResult_lo_10};
  wire [5:0]         checkVec_checkResult_lo_11 = {checkVec_checkResultVec_1_4_1, checkVec_checkResultVec_0_4_1};
  wire [5:0]         checkVec_checkResult_hi_11 = {checkVec_checkResultVec_3_4_1, checkVec_checkResultVec_2_4_1};
  wire [11:0]        checkVec_1_4 = {checkVec_checkResult_hi_11, checkVec_checkResult_lo_11};
  wire [1:0]         checkVec_checkResult_lo_12 = {checkVec_checkResultVec_1_5_1, checkVec_checkResultVec_0_5_1};
  wire [1:0]         checkVec_checkResult_hi_12 = {checkVec_checkResultVec_3_5_1, checkVec_checkResultVec_2_5_1};
  wire [3:0]         checkVec_1_5 = {checkVec_checkResult_hi_12, checkVec_checkResult_lo_12};
  wire [1:0]         checkVec_checkResult_lo_13 = {checkVec_checkResultVec_1_6_1, checkVec_checkResultVec_0_6_1};
  wire [1:0]         checkVec_checkResult_hi_13 = {checkVec_checkResultVec_3_6_1, checkVec_checkResultVec_2_6_1};
  wire [3:0]         checkVec_1_6 = {checkVec_checkResult_hi_13, checkVec_checkResult_lo_13};
  wire               checkVec_checkResultVec_0_6_2 = checkVec_validVec_2[0];
  wire [12:0]        checkVec_checkResultVec_dataPosition_8 = {source_0[10:0], 2'h0};
  wire [1:0]         checkVec_checkResultVec_0_2_2 = checkVec_checkResultVec_dataPosition_8[3:2];
  wire [8:0]         checkVec_checkResultVec_dataGroup_8 = checkVec_checkResultVec_dataPosition_8[12:4];
  wire [5:0]         checkVec_checkResultVec_0_3_2 = checkVec_checkResultVec_dataGroup_8[5:0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_8 = checkVec_checkResultVec_dataGroup_8[8:6];
  wire [2:0]         checkVec_checkResultVec_0_4_2 = checkVec_checkResultVec_accessRegGrowth_8;
  wire [7:0]         checkVec_checkResultVec_decimalProportion_8 = {checkVec_checkResultVec_0_3_2, checkVec_checkResultVec_0_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_8 = checkVec_checkResultVec_decimalProportion_8[7:5];
  wire               checkVec_checkResultVec_overlap_8 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_8 >= checkVec_checkResultVec_intLMULInput_8[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_8} >= checkVec_checkResultVec_intLMULInput_8, source_0[31:13]};
  wire               checkVec_checkResultVec_0_5_2 = checkVec_checkResultVec_overlap_8 | ~checkVec_checkResultVec_0_6_2;
  wire               checkVec_checkResultVec_1_6_2 = checkVec_validVec_2[1];
  wire [12:0]        checkVec_checkResultVec_dataPosition_9 = {source_1[10:0], 2'h0};
  wire [1:0]         checkVec_checkResultVec_1_2_2 = checkVec_checkResultVec_dataPosition_9[3:2];
  wire [8:0]         checkVec_checkResultVec_dataGroup_9 = checkVec_checkResultVec_dataPosition_9[12:4];
  wire [5:0]         checkVec_checkResultVec_1_3_2 = checkVec_checkResultVec_dataGroup_9[5:0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_9 = checkVec_checkResultVec_dataGroup_9[8:6];
  wire [2:0]         checkVec_checkResultVec_1_4_2 = checkVec_checkResultVec_accessRegGrowth_9;
  wire [7:0]         checkVec_checkResultVec_decimalProportion_9 = {checkVec_checkResultVec_1_3_2, checkVec_checkResultVec_1_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_9 = checkVec_checkResultVec_decimalProportion_9[7:5];
  wire               checkVec_checkResultVec_overlap_9 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_9 >= checkVec_checkResultVec_intLMULInput_9[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_9} >= checkVec_checkResultVec_intLMULInput_9, source_1[31:13]};
  wire               checkVec_checkResultVec_1_5_2 = checkVec_checkResultVec_overlap_9 | ~checkVec_checkResultVec_1_6_2;
  wire               checkVec_checkResultVec_2_6_2 = checkVec_validVec_2[2];
  wire [12:0]        checkVec_checkResultVec_dataPosition_10 = {source_2[10:0], 2'h0};
  wire [1:0]         checkVec_checkResultVec_2_2_2 = checkVec_checkResultVec_dataPosition_10[3:2];
  wire [8:0]         checkVec_checkResultVec_dataGroup_10 = checkVec_checkResultVec_dataPosition_10[12:4];
  wire [5:0]         checkVec_checkResultVec_2_3_2 = checkVec_checkResultVec_dataGroup_10[5:0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_10 = checkVec_checkResultVec_dataGroup_10[8:6];
  wire [2:0]         checkVec_checkResultVec_2_4_2 = checkVec_checkResultVec_accessRegGrowth_10;
  wire [7:0]         checkVec_checkResultVec_decimalProportion_10 = {checkVec_checkResultVec_2_3_2, checkVec_checkResultVec_2_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_10 = checkVec_checkResultVec_decimalProportion_10[7:5];
  wire               checkVec_checkResultVec_overlap_10 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_10 >= checkVec_checkResultVec_intLMULInput_10[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_10} >= checkVec_checkResultVec_intLMULInput_10,
      source_2[31:13]};
  wire               checkVec_checkResultVec_2_5_2 = checkVec_checkResultVec_overlap_10 | ~checkVec_checkResultVec_2_6_2;
  wire               checkVec_checkResultVec_3_6_2 = checkVec_validVec_2[3];
  wire [12:0]        checkVec_checkResultVec_dataPosition_11 = {source_3[10:0], 2'h0};
  wire [1:0]         checkVec_checkResultVec_3_2_2 = checkVec_checkResultVec_dataPosition_11[3:2];
  wire [8:0]         checkVec_checkResultVec_dataGroup_11 = checkVec_checkResultVec_dataPosition_11[12:4];
  wire [5:0]         checkVec_checkResultVec_3_3_2 = checkVec_checkResultVec_dataGroup_11[5:0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_11 = checkVec_checkResultVec_dataGroup_11[8:6];
  wire [2:0]         checkVec_checkResultVec_3_4_2 = checkVec_checkResultVec_accessRegGrowth_11;
  wire [7:0]         checkVec_checkResultVec_decimalProportion_11 = {checkVec_checkResultVec_3_3_2, checkVec_checkResultVec_3_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_11 = checkVec_checkResultVec_decimalProportion_11[7:5];
  wire               checkVec_checkResultVec_overlap_11 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_11 >= checkVec_checkResultVec_intLMULInput_11[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_11} >= checkVec_checkResultVec_intLMULInput_11,
      source_3[31:13]};
  wire               checkVec_checkResultVec_3_5_2 = checkVec_checkResultVec_overlap_11 | ~checkVec_checkResultVec_3_6_2;
  wire [3:0]         checkVec_checkResult_lo_16 = {checkVec_checkResultVec_1_2_2, checkVec_checkResultVec_0_2_2};
  wire [3:0]         checkVec_checkResult_hi_16 = {checkVec_checkResultVec_3_2_2, checkVec_checkResultVec_2_2_2};
  wire [7:0]         checkVec_2_2 = {checkVec_checkResult_hi_16, checkVec_checkResult_lo_16};
  wire [11:0]        checkVec_checkResult_lo_17 = {checkVec_checkResultVec_1_3_2, checkVec_checkResultVec_0_3_2};
  wire [11:0]        checkVec_checkResult_hi_17 = {checkVec_checkResultVec_3_3_2, checkVec_checkResultVec_2_3_2};
  wire [23:0]        checkVec_2_3 = {checkVec_checkResult_hi_17, checkVec_checkResult_lo_17};
  wire [5:0]         checkVec_checkResult_lo_18 = {checkVec_checkResultVec_1_4_2, checkVec_checkResultVec_0_4_2};
  wire [5:0]         checkVec_checkResult_hi_18 = {checkVec_checkResultVec_3_4_2, checkVec_checkResultVec_2_4_2};
  wire [11:0]        checkVec_2_4 = {checkVec_checkResult_hi_18, checkVec_checkResult_lo_18};
  wire [1:0]         checkVec_checkResult_lo_19 = {checkVec_checkResultVec_1_5_2, checkVec_checkResultVec_0_5_2};
  wire [1:0]         checkVec_checkResult_hi_19 = {checkVec_checkResultVec_3_5_2, checkVec_checkResultVec_2_5_2};
  wire [3:0]         checkVec_2_5 = {checkVec_checkResult_hi_19, checkVec_checkResult_lo_19};
  wire [1:0]         checkVec_checkResult_lo_20 = {checkVec_checkResultVec_1_6_2, checkVec_checkResultVec_0_6_2};
  wire [1:0]         checkVec_checkResult_hi_20 = {checkVec_checkResultVec_3_6_2, checkVec_checkResultVec_2_6_2};
  wire [3:0]         checkVec_2_6 = {checkVec_checkResult_hi_20, checkVec_checkResult_lo_20};
  wire [7:0]         dataOffsetSelect = (sew1H[0] ? checkVec_0_1 : 8'h0) | (sew1H[1] ? checkVec_1_1 : 8'h0);
  wire [7:0]         accessLaneSelect = (sew1H[0] ? checkVec_0_2 : 8'h0) | (sew1H[1] ? checkVec_1_2 : 8'h0) | (sew1H[2] ? checkVec_2_2 : 8'h0);
  wire [23:0]        offsetSelect = (sew1H[0] ? checkVec_0_3 : 24'h0) | (sew1H[1] ? checkVec_1_3 : 24'h0) | (sew1H[2] ? checkVec_2_3 : 24'h0);
  wire [11:0]        growthSelect = (sew1H[0] ? checkVec_0_4 : 12'h0) | (sew1H[1] ? checkVec_1_4 : 12'h0) | (sew1H[2] ? checkVec_2_4 : 12'h0);
  wire [3:0]         notReadSelect = (sew1H[0] ? checkVec_0_5 : 4'h0) | (sew1H[1] ? checkVec_1_5 : 4'h0) | (sew1H[2] ? checkVec_2_5 : 4'h0);
  wire [3:0]         elementValidSelect = (sew1H[0] ? checkVec_0_6 : 4'h0) | (sew1H[1] ? checkVec_1_6 : 4'h0) | (sew1H[2] ? checkVec_2_6 : 4'h0);
  wire               readTypeRequestDeq;
  wire               waiteStageEnqReady;
  wire               readWaitQueue_deq_valid;
  assign readWaitQueue_deq_valid = ~_readWaitQueue_fifo_empty;
  wire [11:0]        readWaitQueue_dataOut_executeGroup;
  wire [3:0]         readWaitQueue_dataOut_sourceValid;
  wire [3:0]         readWaitQueue_dataOut_replaceVs1;
  wire [3:0]         readWaitQueue_dataOut_needRead;
  wire               readWaitQueue_dataOut_last;
  wire [4:0]         readWaitQueue_dataIn_lo = {readWaitQueue_enq_bits_needRead, readWaitQueue_enq_bits_last};
  wire [15:0]        readWaitQueue_dataIn_hi_hi = {readWaitQueue_enq_bits_executeGroup, readWaitQueue_enq_bits_sourceValid};
  wire [19:0]        readWaitQueue_dataIn_hi = {readWaitQueue_dataIn_hi_hi, readWaitQueue_enq_bits_replaceVs1};
  wire [24:0]        readWaitQueue_dataIn = {readWaitQueue_dataIn_hi, readWaitQueue_dataIn_lo};
  assign readWaitQueue_dataOut_last = _readWaitQueue_fifo_data_out[0];
  assign readWaitQueue_dataOut_needRead = _readWaitQueue_fifo_data_out[4:1];
  assign readWaitQueue_dataOut_replaceVs1 = _readWaitQueue_fifo_data_out[8:5];
  assign readWaitQueue_dataOut_sourceValid = _readWaitQueue_fifo_data_out[12:9];
  assign readWaitQueue_dataOut_executeGroup = _readWaitQueue_fifo_data_out[24:13];
  wire [11:0]        readWaitQueue_deq_bits_executeGroup = readWaitQueue_dataOut_executeGroup;
  wire [3:0]         readWaitQueue_deq_bits_sourceValid = readWaitQueue_dataOut_sourceValid;
  wire [3:0]         readWaitQueue_deq_bits_replaceVs1 = readWaitQueue_dataOut_replaceVs1;
  wire [3:0]         readWaitQueue_deq_bits_needRead = readWaitQueue_dataOut_needRead;
  wire               readWaitQueue_deq_bits_last = readWaitQueue_dataOut_last;
  wire               readWaitQueue_enq_ready = ~_readWaitQueue_fifo_full;
  wire               readWaitQueue_enq_valid;
  wire               readWaitQueue_deq_ready;
  wire               _GEN_165 = lastExecuteGroupDeq | viota;
  assign exeRequestQueue_0_deq_ready = ~exeReqReg_0_valid | _GEN_165;
  assign exeRequestQueue_1_deq_ready = ~exeReqReg_1_valid | _GEN_165;
  assign exeRequestQueue_2_deq_ready = ~exeReqReg_2_valid | _GEN_165;
  assign exeRequestQueue_3_deq_ready = ~exeReqReg_3_valid | _GEN_165;
  wire               isLastExecuteGroup = executeIndex == lastExecuteIndex;
  wire               allDataValid = (exeReqReg_0_valid | ~(groupDataNeed[0])) & (exeReqReg_1_valid | ~(groupDataNeed[1])) & (exeReqReg_2_valid | ~(groupDataNeed[2])) & (exeReqReg_3_valid | ~(groupDataNeed[3]));
  wire               anyDataValid = exeReqReg_0_valid | exeReqReg_1_valid | exeReqReg_2_valid | exeReqReg_3_valid;
  wire               _GEN_166 = compress | mvRd;
  wire               readVs1Valid = (unitType[2] | _GEN_166) & ~readVS1Reg_requestSend | gatherSRead;
  wire [4:0]         readVS1Req_vs = compress ? instReg_vs1 + {4'h0, readVS1Reg_readIndex[8]} : gatherSRead ? instReg_vs1 + {2'h0, gatherGrowth} : instReg_vs1;
  wire [5:0]         readVS1Req_offset = compress ? readVS1Reg_readIndex[7:2] : gatherSRead ? gatherOffset : 6'h0;
  wire [1:0]         readVS1Req_readLane = compress ? readVS1Reg_readIndex[1:0] : gatherSRead ? gatherLane : 2'h0;
  wire [1:0]         readVS1Req_dataOffset = compress | ~gatherSRead ? 2'h0 : gatherDatOffset;
  wire [5:0]         selectExecuteReq_1_bits_offset = readIssueStageState_readOffset[11:6];
  wire [5:0]         selectExecuteReq_2_bits_offset = readIssueStageState_readOffset[17:12];
  wire [5:0]         selectExecuteReq_3_bits_offset = readIssueStageState_readOffset[23:18];
  wire [1:0]         selectExecuteReq_1_bits_dataOffset = readIssueStageState_readDataOffset[3:2];
  wire [1:0]         selectExecuteReq_2_bits_dataOffset = readIssueStageState_readDataOffset[5:4];
  wire [1:0]         selectExecuteReq_3_bits_dataOffset = readIssueStageState_readDataOffset[7:6];
  wire               selectExecuteReq_0_valid = readVs1Valid | readIssueStageValid & ~(readIssueStageState_groupReadState[0]) & readIssueStageState_needRead[0] & readType;
  wire [4:0]         selectExecuteReq_0_bits_vs = readVs1Valid ? readVS1Req_vs : instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_0};
  wire [5:0]         selectExecuteReq_0_bits_offset = readVs1Valid ? readVS1Req_offset : readIssueStageState_readOffset[5:0];
  wire [1:0]         selectExecuteReq_0_bits_readLane = readVs1Valid ? readVS1Req_readLane : readIssueStageState_accessLane_0;
  wire [1:0]         selectExecuteReq_0_bits_dataOffset = readVs1Valid ? readVS1Req_dataOffset : readIssueStageState_readDataOffset[1:0];
  wire               _tokenCheck_T = _readCrossBar_input_0_ready & readCrossBar_input_0_valid;
  wire               pipeReadFire_0 = ~readVs1Valid & _tokenCheck_T;
  wire [4:0]         selectExecuteReq_1_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_1};
  wire               selectExecuteReq_1_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[1]) & readIssueStageState_needRead[1] & readType;
  wire               pipeReadFire_1 = _readCrossBar_input_1_ready & readCrossBar_input_1_valid;
  wire [4:0]         selectExecuteReq_2_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_2};
  wire               selectExecuteReq_2_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[2]) & readIssueStageState_needRead[2] & readType;
  wire               pipeReadFire_2 = _readCrossBar_input_2_ready & readCrossBar_input_2_valid;
  wire [4:0]         selectExecuteReq_3_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_3};
  wire               selectExecuteReq_3_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[3]) & readIssueStageState_needRead[3] & readType;
  wire               pipeReadFire_3 = _readCrossBar_input_3_ready & readCrossBar_input_3_valid;
  reg  [3:0]         tokenCheck_counter;
  wire [3:0]         tokenCheck_counterChange = _tokenCheck_T ? 4'h1 : 4'hF;
  wire               tokenCheck = ~(tokenCheck_counter[3]);
  assign readCrossBar_input_0_valid = selectExecuteReq_0_valid & tokenCheck;
  reg  [3:0]         tokenCheck_counter_1;
  wire [3:0]         tokenCheck_counterChange_1 = pipeReadFire_1 ? 4'h1 : 4'hF;
  wire               tokenCheck_1 = ~(tokenCheck_counter_1[3]);
  assign readCrossBar_input_1_valid = selectExecuteReq_1_valid & tokenCheck_1;
  reg  [3:0]         tokenCheck_counter_2;
  wire [3:0]         tokenCheck_counterChange_2 = pipeReadFire_2 ? 4'h1 : 4'hF;
  wire               tokenCheck_2 = ~(tokenCheck_counter_2[3]);
  assign readCrossBar_input_2_valid = selectExecuteReq_2_valid & tokenCheck_2;
  reg  [3:0]         tokenCheck_counter_3;
  wire [3:0]         tokenCheck_counterChange_3 = pipeReadFire_3 ? 4'h1 : 4'hF;
  wire               tokenCheck_3 = ~(tokenCheck_counter_3[3]);
  assign readCrossBar_input_3_valid = selectExecuteReq_3_valid & tokenCheck_3;
  wire [1:0]         readFire_lo = {pipeReadFire_1, pipeReadFire_0};
  wire [1:0]         readFire_hi = {pipeReadFire_3, pipeReadFire_2};
  wire [3:0]         readFire = {readFire_hi, readFire_lo};
  wire               anyReadFire = |readFire;
  wire [3:0]         readStateUpdate = readFire | readIssueStageState_groupReadState;
  wire               groupReadFinish = readStateUpdate == readIssueStageState_needRead;
  assign readTypeRequestDeq = anyReadFire & groupReadFinish | readIssueStageValid & readIssueStageState_needRead == 4'h0;
  assign readWaitQueue_enq_valid = readTypeRequestDeq;
  wire [3:0]         compressUnitResultQueue_enq_bits_ffoOutput;
  wire               compressUnitResultQueue_enq_bits_compressValid;
  wire [4:0]         compressUnitResultQueue_dataIn_lo = {compressUnitResultQueue_enq_bits_ffoOutput, compressUnitResultQueue_enq_bits_compressValid};
  wire [127:0]       compressUnitResultQueue_enq_bits_data;
  wire [15:0]        compressUnitResultQueue_enq_bits_mask;
  wire [143:0]       compressUnitResultQueue_dataIn_hi_hi = {compressUnitResultQueue_enq_bits_data, compressUnitResultQueue_enq_bits_mask};
  wire [9:0]         compressUnitResultQueue_enq_bits_groupCounter;
  wire [153:0]       compressUnitResultQueue_dataIn_hi = {compressUnitResultQueue_dataIn_hi_hi, compressUnitResultQueue_enq_bits_groupCounter};
  wire [158:0]       compressUnitResultQueue_dataIn = {compressUnitResultQueue_dataIn_hi, compressUnitResultQueue_dataIn_lo};
  wire               compressUnitResultQueue_dataOut_compressValid = _compressUnitResultQueue_fifo_data_out[0];
  wire [3:0]         compressUnitResultQueue_dataOut_ffoOutput = _compressUnitResultQueue_fifo_data_out[4:1];
  wire [9:0]         compressUnitResultQueue_dataOut_groupCounter = _compressUnitResultQueue_fifo_data_out[14:5];
  wire [15:0]        compressUnitResultQueue_dataOut_mask = _compressUnitResultQueue_fifo_data_out[30:15];
  wire [127:0]       compressUnitResultQueue_dataOut_data = _compressUnitResultQueue_fifo_data_out[158:31];
  wire               compressUnitResultQueue_enq_ready = ~_compressUnitResultQueue_fifo_full;
  wire               compressUnitResultQueue_deq_ready;
  wire               compressUnitResultQueue_enq_valid;
  wire               compressUnitResultQueue_deq_valid = ~_compressUnitResultQueue_fifo_empty | compressUnitResultQueue_enq_valid;
  wire [127:0]       compressUnitResultQueue_deq_bits_data = _compressUnitResultQueue_fifo_empty ? compressUnitResultQueue_enq_bits_data : compressUnitResultQueue_dataOut_data;
  wire [15:0]        compressUnitResultQueue_deq_bits_mask = _compressUnitResultQueue_fifo_empty ? compressUnitResultQueue_enq_bits_mask : compressUnitResultQueue_dataOut_mask;
  wire [9:0]         compressUnitResultQueue_deq_bits_groupCounter = _compressUnitResultQueue_fifo_empty ? compressUnitResultQueue_enq_bits_groupCounter : compressUnitResultQueue_dataOut_groupCounter;
  wire [3:0]         compressUnitResultQueue_deq_bits_ffoOutput = _compressUnitResultQueue_fifo_empty ? compressUnitResultQueue_enq_bits_ffoOutput : compressUnitResultQueue_dataOut_ffoOutput;
  wire               compressUnitResultQueue_deq_bits_compressValid = _compressUnitResultQueue_fifo_empty ? compressUnitResultQueue_enq_bits_compressValid : compressUnitResultQueue_dataOut_compressValid;
  wire               noSourceValid = noSource & counterValid & ((|instReg_vl) | mvRd & ~readVS1Reg_sendToExecution);
  wire               vs1DataValid = readVS1Reg_dataValid | ~(unitType[2] | _GEN_166);
  wire [1:0]         _GEN_167 = {_maskedWrite_in_1_ready, _maskedWrite_in_0_ready};
  wire [1:0]         executeDeqReady_lo;
  assign executeDeqReady_lo = _GEN_167;
  wire [1:0]         compressUnitResultQueue_deq_ready_lo;
  assign compressUnitResultQueue_deq_ready_lo = _GEN_167;
  wire [1:0]         _GEN_168 = {_maskedWrite_in_3_ready, _maskedWrite_in_2_ready};
  wire [1:0]         executeDeqReady_hi;
  assign executeDeqReady_hi = _GEN_168;
  wire [1:0]         compressUnitResultQueue_deq_ready_hi;
  assign compressUnitResultQueue_deq_ready_hi = _GEN_168;
  wire               compressUnitResultQueue_empty;
  wire               executeDeqReady = (&{executeDeqReady_hi, executeDeqReady_lo}) & compressUnitResultQueue_empty;
  wire               otherTypeRequestDeq = (noSource ? noSourceValid : allDataValid) & vs1DataValid & instVlValid & executeDeqReady;
  wire               reorderQueueAllocate;
  wire               _GEN_169 = accessCountQueue_enq_ready & reorderQueueAllocate;
  assign readIssueStageEnq = (allDataValid | _slideAddressGen_indexDeq_valid) & (readTypeRequestDeq | ~readIssueStageValid) & instVlValid & readType & _GEN_169;
  assign accessCountQueue_enq_valid = readIssueStageEnq;
  wire               executeReady;
  wire               requestStageDeq = readType ? readIssueStageEnq : otherTypeRequestDeq & executeReady;
  wire               slideAddressGen_indexDeq_ready = (readTypeRequestDeq | ~readIssueStageValid) & _GEN_169;
  wire               _GEN_170 = slideAddressGen_indexDeq_ready & _slideAddressGen_indexDeq_valid;
  wire               _GEN_171 = readIssueStageEnq & _GEN_170;
  assign accessCountEnq_0 =
    _GEN_171
      ? {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 2'h0 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 2'h0 & _slideAddressGen_indexDeq_bits_needRead[1]}}
        + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 2'h0 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 2'h0 & _slideAddressGen_indexDeq_bits_needRead[3]}}
      : {1'h0, {1'h0, accessLaneSelect[1:0] == 2'h0 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[3:2] == 2'h0 & ~(notReadSelect[1])}}
        + {1'h0, {1'h0, accessLaneSelect[5:4] == 2'h0 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[7:6] == 2'h0 & ~(notReadSelect[3])}};
  assign accessCountEnq_1 =
    _GEN_171
      ? {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 2'h1 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 2'h1 & _slideAddressGen_indexDeq_bits_needRead[1]}}
        + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 2'h1 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 2'h1 & _slideAddressGen_indexDeq_bits_needRead[3]}}
      : {1'h0, {1'h0, accessLaneSelect[1:0] == 2'h1 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[3:2] == 2'h1 & ~(notReadSelect[1])}}
        + {1'h0, {1'h0, accessLaneSelect[5:4] == 2'h1 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[7:6] == 2'h1 & ~(notReadSelect[3])}};
  assign accessCountEnq_2 =
    _GEN_171
      ? {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 2'h2 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 2'h2 & _slideAddressGen_indexDeq_bits_needRead[1]}}
        + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 2'h2 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 2'h2 & _slideAddressGen_indexDeq_bits_needRead[3]}}
      : {1'h0, {1'h0, accessLaneSelect[1:0] == 2'h2 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[3:2] == 2'h2 & ~(notReadSelect[1])}}
        + {1'h0, {1'h0, accessLaneSelect[5:4] == 2'h2 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[7:6] == 2'h2 & ~(notReadSelect[3])}};
  assign accessCountEnq_3 =
    _GEN_171
      ? {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_0) & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_1) & _slideAddressGen_indexDeq_bits_needRead[1]}}
        + {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_2) & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_3) & _slideAddressGen_indexDeq_bits_needRead[3]}}
      : {1'h0, {1'h0, (&(accessLaneSelect[1:0])) & ~(notReadSelect[0])} + {1'h0, (&(accessLaneSelect[3:2])) & ~(notReadSelect[1])}}
        + {1'h0, {1'h0, (&(accessLaneSelect[5:4])) & ~(notReadSelect[2])} + {1'h0, (&(accessLaneSelect[7:6])) & ~(notReadSelect[3])}};
  assign lastExecuteGroupDeq = requestStageDeq & isLastExecuteGroup;
  wire [3:0]         readMessageQueue_deq_bits_readSource;
  wire               deqAllocate;
  wire               reorderQueueVec_0_deq_valid;
  assign reorderQueueVec_0_deq_valid = ~_reorderQueueVec_fifo_empty;
  wire [31:0]        reorderQueueVec_dataOut_data;
  wire [3:0]         reorderQueueVec_dataOut_write1H;
  wire [31:0]        dataAfterReorderCheck_0 = reorderQueueVec_0_deq_bits_data;
  wire [31:0]        reorderQueueVec_0_enq_bits_data;
  wire [3:0]         reorderQueueVec_0_enq_bits_write1H;
  wire [35:0]        reorderQueueVec_dataIn = {reorderQueueVec_0_enq_bits_data, reorderQueueVec_0_enq_bits_write1H};
  assign reorderQueueVec_dataOut_write1H = _reorderQueueVec_fifo_data_out[3:0];
  assign reorderQueueVec_dataOut_data = _reorderQueueVec_fifo_data_out[35:4];
  assign reorderQueueVec_0_deq_bits_data = reorderQueueVec_dataOut_data;
  wire [3:0]         reorderQueueVec_0_deq_bits_write1H = reorderQueueVec_dataOut_write1H;
  wire               reorderQueueVec_0_enq_ready = ~_reorderQueueVec_fifo_full;
  wire               reorderQueueVec_0_deq_ready;
  wire [3:0]         readMessageQueue_1_deq_bits_readSource;
  wire               deqAllocate_1;
  wire               reorderQueueVec_1_deq_valid;
  assign reorderQueueVec_1_deq_valid = ~_reorderQueueVec_fifo_1_empty;
  wire [31:0]        reorderQueueVec_dataOut_1_data;
  wire [3:0]         reorderQueueVec_dataOut_1_write1H;
  wire [31:0]        dataAfterReorderCheck_1 = reorderQueueVec_1_deq_bits_data;
  wire [31:0]        reorderQueueVec_1_enq_bits_data;
  wire [3:0]         reorderQueueVec_1_enq_bits_write1H;
  wire [35:0]        reorderQueueVec_dataIn_1 = {reorderQueueVec_1_enq_bits_data, reorderQueueVec_1_enq_bits_write1H};
  assign reorderQueueVec_dataOut_1_write1H = _reorderQueueVec_fifo_1_data_out[3:0];
  assign reorderQueueVec_dataOut_1_data = _reorderQueueVec_fifo_1_data_out[35:4];
  assign reorderQueueVec_1_deq_bits_data = reorderQueueVec_dataOut_1_data;
  wire [3:0]         reorderQueueVec_1_deq_bits_write1H = reorderQueueVec_dataOut_1_write1H;
  wire               reorderQueueVec_1_enq_ready = ~_reorderQueueVec_fifo_1_full;
  wire               reorderQueueVec_1_deq_ready;
  wire [3:0]         readMessageQueue_2_deq_bits_readSource;
  wire               deqAllocate_2;
  wire               reorderQueueVec_2_deq_valid;
  assign reorderQueueVec_2_deq_valid = ~_reorderQueueVec_fifo_2_empty;
  wire [31:0]        reorderQueueVec_dataOut_2_data;
  wire [3:0]         reorderQueueVec_dataOut_2_write1H;
  wire [31:0]        dataAfterReorderCheck_2 = reorderQueueVec_2_deq_bits_data;
  wire [31:0]        reorderQueueVec_2_enq_bits_data;
  wire [3:0]         reorderQueueVec_2_enq_bits_write1H;
  wire [35:0]        reorderQueueVec_dataIn_2 = {reorderQueueVec_2_enq_bits_data, reorderQueueVec_2_enq_bits_write1H};
  assign reorderQueueVec_dataOut_2_write1H = _reorderQueueVec_fifo_2_data_out[3:0];
  assign reorderQueueVec_dataOut_2_data = _reorderQueueVec_fifo_2_data_out[35:4];
  assign reorderQueueVec_2_deq_bits_data = reorderQueueVec_dataOut_2_data;
  wire [3:0]         reorderQueueVec_2_deq_bits_write1H = reorderQueueVec_dataOut_2_write1H;
  wire               reorderQueueVec_2_enq_ready = ~_reorderQueueVec_fifo_2_full;
  wire               reorderQueueVec_2_deq_ready;
  wire [3:0]         readMessageQueue_3_deq_bits_readSource;
  wire               deqAllocate_3;
  wire               reorderQueueVec_3_deq_valid;
  assign reorderQueueVec_3_deq_valid = ~_reorderQueueVec_fifo_3_empty;
  wire [31:0]        reorderQueueVec_dataOut_3_data;
  wire [3:0]         reorderQueueVec_dataOut_3_write1H;
  wire [31:0]        dataAfterReorderCheck_3 = reorderQueueVec_3_deq_bits_data;
  wire [31:0]        reorderQueueVec_3_enq_bits_data;
  wire [3:0]         reorderQueueVec_3_enq_bits_write1H;
  wire [35:0]        reorderQueueVec_dataIn_3 = {reorderQueueVec_3_enq_bits_data, reorderQueueVec_3_enq_bits_write1H};
  assign reorderQueueVec_dataOut_3_write1H = _reorderQueueVec_fifo_3_data_out[3:0];
  assign reorderQueueVec_dataOut_3_data = _reorderQueueVec_fifo_3_data_out[35:4];
  assign reorderQueueVec_3_deq_bits_data = reorderQueueVec_dataOut_3_data;
  wire [3:0]         reorderQueueVec_3_deq_bits_write1H = reorderQueueVec_dataOut_3_write1H;
  wire               reorderQueueVec_3_enq_ready = ~_reorderQueueVec_fifo_3_full;
  wire               reorderQueueVec_3_deq_ready;
  reg  [3:0]         reorderQueueAllocate_counter;
  reg  [3:0]         reorderQueueAllocate_counterWillUpdate;
  wire               _write1HPipe_0_T = reorderQueueVec_0_deq_ready & reorderQueueVec_0_deq_valid;
  wire               reorderQueueAllocate_release = _write1HPipe_0_T & readValid;
  wire [2:0]         reorderQueueAllocate_allocate = readIssueStageEnq ? accessCountEnq_0 : 3'h0;
  wire [3:0]         reorderQueueAllocate_counterUpdate = reorderQueueAllocate_counter + {1'h0, reorderQueueAllocate_allocate} - {3'h0, reorderQueueAllocate_release};
  reg  [3:0]         reorderQueueAllocate_counter_1;
  reg  [3:0]         reorderQueueAllocate_counterWillUpdate_1;
  wire               _write1HPipe_1_T = reorderQueueVec_1_deq_ready & reorderQueueVec_1_deq_valid;
  wire               reorderQueueAllocate_release_1 = _write1HPipe_1_T & readValid;
  wire [2:0]         reorderQueueAllocate_allocate_1 = readIssueStageEnq ? accessCountEnq_1 : 3'h0;
  wire [3:0]         reorderQueueAllocate_counterUpdate_1 = reorderQueueAllocate_counter_1 + {1'h0, reorderQueueAllocate_allocate_1} - {3'h0, reorderQueueAllocate_release_1};
  reg  [3:0]         reorderQueueAllocate_counter_2;
  reg  [3:0]         reorderQueueAllocate_counterWillUpdate_2;
  wire               _write1HPipe_2_T = reorderQueueVec_2_deq_ready & reorderQueueVec_2_deq_valid;
  wire               reorderQueueAllocate_release_2 = _write1HPipe_2_T & readValid;
  wire [2:0]         reorderQueueAllocate_allocate_2 = readIssueStageEnq ? accessCountEnq_2 : 3'h0;
  wire [3:0]         reorderQueueAllocate_counterUpdate_2 = reorderQueueAllocate_counter_2 + {1'h0, reorderQueueAllocate_allocate_2} - {3'h0, reorderQueueAllocate_release_2};
  reg  [3:0]         reorderQueueAllocate_counter_3;
  reg  [3:0]         reorderQueueAllocate_counterWillUpdate_3;
  wire               _write1HPipe_3_T = reorderQueueVec_3_deq_ready & reorderQueueVec_3_deq_valid;
  wire               reorderQueueAllocate_release_3 = _write1HPipe_3_T & readValid;
  wire [2:0]         reorderQueueAllocate_allocate_3 = readIssueStageEnq ? accessCountEnq_3 : 3'h0;
  wire [3:0]         reorderQueueAllocate_counterUpdate_3 = reorderQueueAllocate_counter_3 + {1'h0, reorderQueueAllocate_allocate_3} - {3'h0, reorderQueueAllocate_release_3};
  assign reorderQueueAllocate = ~(reorderQueueAllocate_counterWillUpdate[3]) & ~(reorderQueueAllocate_counterWillUpdate_1[3]) & ~(reorderQueueAllocate_counterWillUpdate_2[3]) & ~(reorderQueueAllocate_counterWillUpdate_3[3]);
  reg                reorderStageValid;
  reg  [2:0]         reorderStageState_0;
  reg  [2:0]         reorderStageState_1;
  reg  [2:0]         reorderStageState_2;
  reg  [2:0]         reorderStageState_3;
  reg  [2:0]         reorderStageNeed_0;
  reg  [2:0]         reorderStageNeed_1;
  reg  [2:0]         reorderStageNeed_2;
  reg  [2:0]         reorderStageNeed_3;
  wire               stateCheck = reorderStageState_0 == reorderStageNeed_0 & reorderStageState_1 == reorderStageNeed_1 & reorderStageState_2 == reorderStageNeed_2 & reorderStageState_3 == reorderStageNeed_3;
  assign accessCountQueue_deq_ready = ~reorderStageValid | stateCheck;
  wire               reorderStageEnqFire = accessCountQueue_deq_ready & accessCountQueue_deq_valid;
  wire               reorderStageDeqFire = stateCheck & reorderStageValid;
  wire [3:0]         sourceLane;
  wire               readMessageQueue_deq_valid;
  assign readMessageQueue_deq_valid = ~_readMessageQueue_fifo_empty;
  wire [3:0]         readMessageQueue_dataOut_readSource;
  assign reorderQueueVec_0_enq_bits_write1H = readMessageQueue_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_dataOffset;
  wire [3:0]         readMessageQueue_enq_bits_readSource;
  wire [1:0]         readMessageQueue_enq_bits_dataOffset;
  wire [5:0]         readMessageQueue_dataIn = {readMessageQueue_enq_bits_readSource, readMessageQueue_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_dataOffset = _readMessageQueue_fifo_data_out[1:0];
  assign readMessageQueue_dataOut_readSource = _readMessageQueue_fifo_data_out[5:2];
  assign readMessageQueue_deq_bits_readSource = readMessageQueue_dataOut_readSource;
  wire [1:0]         readMessageQueue_deq_bits_dataOffset = readMessageQueue_dataOut_dataOffset;
  wire               readMessageQueue_enq_ready = ~_readMessageQueue_fifo_full;
  wire               readMessageQueue_enq_valid;
  assign deqAllocate = ~readValid | reorderStageValid & reorderStageState_0 != reorderStageNeed_0;
  assign reorderQueueVec_0_deq_ready = deqAllocate;
  assign sourceLane = 4'h1 << _readCrossBar_output_0_bits_writeIndex;
  assign readMessageQueue_enq_bits_readSource = sourceLane;
  wire               readChannel_0_valid_0 = maskDestinationType ? _maskedWrite_readChannel_0_valid : _readCrossBar_output_0_valid & readMessageQueue_enq_ready;
  wire [4:0]         readChannel_0_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_0_bits_vs : _readCrossBar_output_0_bits_vs;
  wire [5:0]         readChannel_0_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_0_bits_offset : _readCrossBar_output_0_bits_offset;
  assign readMessageQueue_enq_valid = readChannel_0_ready_0 & readChannel_0_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_0_enq_bits_data = readResult_0_bits >> {27'h0, readMessageQueue_deq_bits_dataOffset, 3'h0};
  wire [3:0]         write1HPipe_0 = _write1HPipe_0_T & ~maskDestinationType ? reorderQueueVec_0_deq_bits_write1H : 4'h0;
  wire [3:0]         sourceLane_1;
  wire               readMessageQueue_1_deq_valid;
  assign readMessageQueue_1_deq_valid = ~_readMessageQueue_fifo_1_empty;
  wire [3:0]         readMessageQueue_dataOut_1_readSource;
  assign reorderQueueVec_1_enq_bits_write1H = readMessageQueue_1_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_1_dataOffset;
  wire [3:0]         readMessageQueue_1_enq_bits_readSource;
  wire [1:0]         readMessageQueue_1_enq_bits_dataOffset;
  wire [5:0]         readMessageQueue_dataIn_1 = {readMessageQueue_1_enq_bits_readSource, readMessageQueue_1_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_1_dataOffset = _readMessageQueue_fifo_1_data_out[1:0];
  assign readMessageQueue_dataOut_1_readSource = _readMessageQueue_fifo_1_data_out[5:2];
  assign readMessageQueue_1_deq_bits_readSource = readMessageQueue_dataOut_1_readSource;
  wire [1:0]         readMessageQueue_1_deq_bits_dataOffset = readMessageQueue_dataOut_1_dataOffset;
  wire               readMessageQueue_1_enq_ready = ~_readMessageQueue_fifo_1_full;
  wire               readMessageQueue_1_enq_valid;
  assign deqAllocate_1 = ~readValid | reorderStageValid & reorderStageState_1 != reorderStageNeed_1;
  assign reorderQueueVec_1_deq_ready = deqAllocate_1;
  assign sourceLane_1 = 4'h1 << _readCrossBar_output_1_bits_writeIndex;
  assign readMessageQueue_1_enq_bits_readSource = sourceLane_1;
  wire               readChannel_1_valid_0 = maskDestinationType ? _maskedWrite_readChannel_1_valid : _readCrossBar_output_1_valid & readMessageQueue_1_enq_ready;
  wire [4:0]         readChannel_1_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_1_bits_vs : _readCrossBar_output_1_bits_vs;
  wire [5:0]         readChannel_1_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_1_bits_offset : _readCrossBar_output_1_bits_offset;
  assign readMessageQueue_1_enq_valid = readChannel_1_ready_0 & readChannel_1_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_1_enq_bits_data = readResult_1_bits >> {27'h0, readMessageQueue_1_deq_bits_dataOffset, 3'h0};
  wire [3:0]         write1HPipe_1 = _write1HPipe_1_T & ~maskDestinationType ? reorderQueueVec_1_deq_bits_write1H : 4'h0;
  wire [3:0]         sourceLane_2;
  wire               readMessageQueue_2_deq_valid;
  assign readMessageQueue_2_deq_valid = ~_readMessageQueue_fifo_2_empty;
  wire [3:0]         readMessageQueue_dataOut_2_readSource;
  assign reorderQueueVec_2_enq_bits_write1H = readMessageQueue_2_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_2_dataOffset;
  wire [3:0]         readMessageQueue_2_enq_bits_readSource;
  wire [1:0]         readMessageQueue_2_enq_bits_dataOffset;
  wire [5:0]         readMessageQueue_dataIn_2 = {readMessageQueue_2_enq_bits_readSource, readMessageQueue_2_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_2_dataOffset = _readMessageQueue_fifo_2_data_out[1:0];
  assign readMessageQueue_dataOut_2_readSource = _readMessageQueue_fifo_2_data_out[5:2];
  assign readMessageQueue_2_deq_bits_readSource = readMessageQueue_dataOut_2_readSource;
  wire [1:0]         readMessageQueue_2_deq_bits_dataOffset = readMessageQueue_dataOut_2_dataOffset;
  wire               readMessageQueue_2_enq_ready = ~_readMessageQueue_fifo_2_full;
  wire               readMessageQueue_2_enq_valid;
  assign deqAllocate_2 = ~readValid | reorderStageValid & reorderStageState_2 != reorderStageNeed_2;
  assign reorderQueueVec_2_deq_ready = deqAllocate_2;
  assign sourceLane_2 = 4'h1 << _readCrossBar_output_2_bits_writeIndex;
  assign readMessageQueue_2_enq_bits_readSource = sourceLane_2;
  wire               readChannel_2_valid_0 = maskDestinationType ? _maskedWrite_readChannel_2_valid : _readCrossBar_output_2_valid & readMessageQueue_2_enq_ready;
  wire [4:0]         readChannel_2_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_2_bits_vs : _readCrossBar_output_2_bits_vs;
  wire [5:0]         readChannel_2_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_2_bits_offset : _readCrossBar_output_2_bits_offset;
  assign readMessageQueue_2_enq_valid = readChannel_2_ready_0 & readChannel_2_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_2_enq_bits_data = readResult_2_bits >> {27'h0, readMessageQueue_2_deq_bits_dataOffset, 3'h0};
  wire [3:0]         write1HPipe_2 = _write1HPipe_2_T & ~maskDestinationType ? reorderQueueVec_2_deq_bits_write1H : 4'h0;
  wire [3:0]         sourceLane_3;
  wire               readMessageQueue_3_deq_valid;
  assign readMessageQueue_3_deq_valid = ~_readMessageQueue_fifo_3_empty;
  wire [3:0]         readMessageQueue_dataOut_3_readSource;
  assign reorderQueueVec_3_enq_bits_write1H = readMessageQueue_3_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_3_dataOffset;
  wire [3:0]         readMessageQueue_3_enq_bits_readSource;
  wire [1:0]         readMessageQueue_3_enq_bits_dataOffset;
  wire [5:0]         readMessageQueue_dataIn_3 = {readMessageQueue_3_enq_bits_readSource, readMessageQueue_3_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_3_dataOffset = _readMessageQueue_fifo_3_data_out[1:0];
  assign readMessageQueue_dataOut_3_readSource = _readMessageQueue_fifo_3_data_out[5:2];
  assign readMessageQueue_3_deq_bits_readSource = readMessageQueue_dataOut_3_readSource;
  wire [1:0]         readMessageQueue_3_deq_bits_dataOffset = readMessageQueue_dataOut_3_dataOffset;
  wire               readMessageQueue_3_enq_ready = ~_readMessageQueue_fifo_3_full;
  wire               readMessageQueue_3_enq_valid;
  assign deqAllocate_3 = ~readValid | reorderStageValid & reorderStageState_3 != reorderStageNeed_3;
  assign reorderQueueVec_3_deq_ready = deqAllocate_3;
  assign sourceLane_3 = 4'h1 << _readCrossBar_output_3_bits_writeIndex;
  assign readMessageQueue_3_enq_bits_readSource = sourceLane_3;
  wire               readChannel_3_valid_0 = maskDestinationType ? _maskedWrite_readChannel_3_valid : _readCrossBar_output_3_valid & readMessageQueue_3_enq_ready;
  wire [4:0]         readChannel_3_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_3_bits_vs : _readCrossBar_output_3_bits_vs;
  wire [5:0]         readChannel_3_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_3_bits_offset : _readCrossBar_output_3_bits_offset;
  assign readMessageQueue_3_enq_valid = readChannel_3_ready_0 & readChannel_3_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_3_enq_bits_data = readResult_3_bits >> {27'h0, readMessageQueue_3_deq_bits_dataOffset, 3'h0};
  wire [3:0]         write1HPipe_3 = _write1HPipe_3_T & ~maskDestinationType ? reorderQueueVec_3_deq_bits_write1H : 4'h0;
  wire [31:0]        readData_data;
  wire               readData_readDataQueue_enq_ready = ~_readData_readDataQueue_fifo_full;
  wire               readData_readDataQueue_deq_ready;
  wire               readData_readDataQueue_enq_valid;
  wire               readData_readDataQueue_deq_valid = ~_readData_readDataQueue_fifo_empty | readData_readDataQueue_enq_valid;
  wire [31:0]        readData_readDataQueue_enq_bits;
  wire [31:0]        readData_readDataQueue_deq_bits = _readData_readDataQueue_fifo_empty ? readData_readDataQueue_enq_bits : _readData_readDataQueue_fifo_data_out;
  wire [1:0]         readData_readResultSelect_lo = {write1HPipe_1[0], write1HPipe_0[0]};
  wire [1:0]         readData_readResultSelect_hi = {write1HPipe_3[0], write1HPipe_2[0]};
  wire [3:0]         readData_readResultSelect = {readData_readResultSelect_hi, readData_readResultSelect_lo};
  assign readData_data =
    (readData_readResultSelect[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect[3] ? dataAfterReorderCheck_3 : 32'h0);
  assign readData_readDataQueue_enq_bits = readData_data;
  wire               readTokenRelease_0 = readData_readDataQueue_deq_ready & readData_readDataQueue_deq_valid;
  assign readData_readDataQueue_enq_valid = |readData_readResultSelect;
  wire [31:0]        readData_data_1;
  wire               isWaiteForThisData_1;
  wire               readData_readDataQueue_1_enq_ready = ~_readData_readDataQueue_fifo_1_full;
  wire               readData_readDataQueue_1_deq_ready;
  wire               readData_readDataQueue_1_enq_valid;
  wire               readData_readDataQueue_1_deq_valid = ~_readData_readDataQueue_fifo_1_empty | readData_readDataQueue_1_enq_valid;
  wire [31:0]        readData_readDataQueue_1_enq_bits;
  wire [31:0]        readData_readDataQueue_1_deq_bits = _readData_readDataQueue_fifo_1_empty ? readData_readDataQueue_1_enq_bits : _readData_readDataQueue_fifo_1_data_out;
  wire [1:0]         readData_readResultSelect_lo_1 = {write1HPipe_1[1], write1HPipe_0[1]};
  wire [1:0]         readData_readResultSelect_hi_1 = {write1HPipe_3[1], write1HPipe_2[1]};
  wire [3:0]         readData_readResultSelect_1 = {readData_readResultSelect_hi_1, readData_readResultSelect_lo_1};
  assign readData_data_1 =
    (readData_readResultSelect_1[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_1[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_1[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_1[3] ? dataAfterReorderCheck_3 : 32'h0);
  assign readData_readDataQueue_1_enq_bits = readData_data_1;
  wire               readTokenRelease_1 = readData_readDataQueue_1_deq_ready & readData_readDataQueue_1_deq_valid;
  assign readData_readDataQueue_1_enq_valid = |readData_readResultSelect_1;
  wire [31:0]        readData_data_2;
  wire               isWaiteForThisData_2;
  wire               readData_readDataQueue_2_enq_ready = ~_readData_readDataQueue_fifo_2_full;
  wire               readData_readDataQueue_2_deq_ready;
  wire               readData_readDataQueue_2_enq_valid;
  wire               readData_readDataQueue_2_deq_valid = ~_readData_readDataQueue_fifo_2_empty | readData_readDataQueue_2_enq_valid;
  wire [31:0]        readData_readDataQueue_2_enq_bits;
  wire [31:0]        readData_readDataQueue_2_deq_bits = _readData_readDataQueue_fifo_2_empty ? readData_readDataQueue_2_enq_bits : _readData_readDataQueue_fifo_2_data_out;
  wire [1:0]         readData_readResultSelect_lo_2 = {write1HPipe_1[2], write1HPipe_0[2]};
  wire [1:0]         readData_readResultSelect_hi_2 = {write1HPipe_3[2], write1HPipe_2[2]};
  wire [3:0]         readData_readResultSelect_2 = {readData_readResultSelect_hi_2, readData_readResultSelect_lo_2};
  assign readData_data_2 =
    (readData_readResultSelect_2[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_2[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_2[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_2[3] ? dataAfterReorderCheck_3 : 32'h0);
  assign readData_readDataQueue_2_enq_bits = readData_data_2;
  wire               readTokenRelease_2 = readData_readDataQueue_2_deq_ready & readData_readDataQueue_2_deq_valid;
  assign readData_readDataQueue_2_enq_valid = |readData_readResultSelect_2;
  wire [31:0]        readData_data_3;
  wire               isWaiteForThisData_3;
  wire               readData_readDataQueue_3_enq_ready = ~_readData_readDataQueue_fifo_3_full;
  wire               readData_readDataQueue_3_deq_ready;
  wire               readData_readDataQueue_3_enq_valid;
  wire               readData_readDataQueue_3_deq_valid = ~_readData_readDataQueue_fifo_3_empty | readData_readDataQueue_3_enq_valid;
  wire [31:0]        readData_readDataQueue_3_enq_bits;
  wire [31:0]        readData_readDataQueue_3_deq_bits = _readData_readDataQueue_fifo_3_empty ? readData_readDataQueue_3_enq_bits : _readData_readDataQueue_fifo_3_data_out;
  wire [1:0]         readData_readResultSelect_lo_3 = {write1HPipe_1[3], write1HPipe_0[3]};
  wire [1:0]         readData_readResultSelect_hi_3 = {write1HPipe_3[3], write1HPipe_2[3]};
  wire [3:0]         readData_readResultSelect_3 = {readData_readResultSelect_hi_3, readData_readResultSelect_lo_3};
  assign readData_data_3 =
    (readData_readResultSelect_3[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_3[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_3[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_3[3] ? dataAfterReorderCheck_3 : 32'h0);
  assign readData_readDataQueue_3_enq_bits = readData_data_3;
  wire               readTokenRelease_3 = readData_readDataQueue_3_deq_ready & readData_readDataQueue_3_deq_valid;
  assign readData_readDataQueue_3_enq_valid = |readData_readResultSelect_3;
  reg  [11:0]        waiteReadDataPipeReg_executeGroup;
  reg  [3:0]         waiteReadDataPipeReg_sourceValid;
  reg  [3:0]         waiteReadDataPipeReg_replaceVs1;
  reg  [3:0]         waiteReadDataPipeReg_needRead;
  reg                waiteReadDataPipeReg_last;
  reg  [31:0]        waiteReadData_0;
  reg  [31:0]        waiteReadData_1;
  reg  [31:0]        waiteReadData_2;
  reg  [31:0]        waiteReadData_3;
  reg  [3:0]         waiteReadSate;
  reg                waiteReadStageValid;
  wire [1:0]         executeIndexVec_0 = waiteReadDataPipeReg_executeGroup[1:0];
  wire [1:0]         executeIndexVec_1 = {waiteReadDataPipeReg_executeGroup[0], 1'h0};
  wire               writeDataVec_data_dataIsRead = waiteReadDataPipeReg_needRead[0];
  wire               writeDataVec_data_dataIsRead_4 = waiteReadDataPipeReg_needRead[0];
  wire               writeDataVec_data_dataIsRead_8 = waiteReadDataPipeReg_needRead[0];
  wire [31:0]        _GEN_172 = waiteReadDataPipeReg_replaceVs1[0] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData;
  assign writeDataVec_data_unreadData = _GEN_172;
  wire [31:0]        writeDataVec_data_unreadData_4;
  assign writeDataVec_data_unreadData_4 = _GEN_172;
  wire [31:0]        writeDataVec_data_unreadData_8;
  assign writeDataVec_data_unreadData_8 = _GEN_172;
  wire [7:0]         writeDataVec_data_dataElement = writeDataVec_data_dataIsRead ? waiteReadData_0[7:0] : writeDataVec_data_unreadData[7:0];
  wire               writeDataVec_data_dataIsRead_1 = waiteReadDataPipeReg_needRead[1];
  wire               writeDataVec_data_dataIsRead_5 = waiteReadDataPipeReg_needRead[1];
  wire               writeDataVec_data_dataIsRead_9 = waiteReadDataPipeReg_needRead[1];
  wire [31:0]        _GEN_173 = waiteReadDataPipeReg_replaceVs1[1] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_1;
  assign writeDataVec_data_unreadData_1 = _GEN_173;
  wire [31:0]        writeDataVec_data_unreadData_5;
  assign writeDataVec_data_unreadData_5 = _GEN_173;
  wire [31:0]        writeDataVec_data_unreadData_9;
  assign writeDataVec_data_unreadData_9 = _GEN_173;
  wire [7:0]         writeDataVec_data_dataElement_1 = writeDataVec_data_dataIsRead_1 ? waiteReadData_1[7:0] : writeDataVec_data_unreadData_1[7:0];
  wire               writeDataVec_data_dataIsRead_2 = waiteReadDataPipeReg_needRead[2];
  wire               writeDataVec_data_dataIsRead_6 = waiteReadDataPipeReg_needRead[2];
  wire               writeDataVec_data_dataIsRead_10 = waiteReadDataPipeReg_needRead[2];
  wire [31:0]        _GEN_174 = waiteReadDataPipeReg_replaceVs1[2] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_2;
  assign writeDataVec_data_unreadData_2 = _GEN_174;
  wire [31:0]        writeDataVec_data_unreadData_6;
  assign writeDataVec_data_unreadData_6 = _GEN_174;
  wire [31:0]        writeDataVec_data_unreadData_10;
  assign writeDataVec_data_unreadData_10 = _GEN_174;
  wire [7:0]         writeDataVec_data_dataElement_2 = writeDataVec_data_dataIsRead_2 ? waiteReadData_2[7:0] : writeDataVec_data_unreadData_2[7:0];
  wire               writeDataVec_data_dataIsRead_3 = waiteReadDataPipeReg_needRead[3];
  wire               writeDataVec_data_dataIsRead_7 = waiteReadDataPipeReg_needRead[3];
  wire               writeDataVec_data_dataIsRead_11 = waiteReadDataPipeReg_needRead[3];
  wire [31:0]        _GEN_175 = waiteReadDataPipeReg_replaceVs1[3] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_3;
  assign writeDataVec_data_unreadData_3 = _GEN_175;
  wire [31:0]        writeDataVec_data_unreadData_7;
  assign writeDataVec_data_unreadData_7 = _GEN_175;
  wire [31:0]        writeDataVec_data_unreadData_11;
  assign writeDataVec_data_unreadData_11 = _GEN_175;
  wire [7:0]         writeDataVec_data_dataElement_3 = writeDataVec_data_dataIsRead_3 ? waiteReadData_3[7:0] : writeDataVec_data_unreadData_3[7:0];
  wire [15:0]        writeDataVec_data_lo = {writeDataVec_data_dataElement_1, writeDataVec_data_dataElement};
  wire [15:0]        writeDataVec_data_hi = {writeDataVec_data_dataElement_3, writeDataVec_data_dataElement_2};
  wire [31:0]        writeDataVec_data = {writeDataVec_data_hi, writeDataVec_data_lo};
  wire [158:0]       writeDataVec_shifterData = {127'h0, writeDataVec_data} << {152'h0, executeIndexVec_0, 5'h0};
  wire [127:0]       writeDataVec_0 = writeDataVec_shifterData[127:0];
  wire [15:0]        writeDataVec_data_dataElement_4 = writeDataVec_data_dataIsRead_4 ? waiteReadData_0[15:0] : writeDataVec_data_unreadData_4[15:0];
  wire [15:0]        writeDataVec_data_dataElement_5 = writeDataVec_data_dataIsRead_5 ? waiteReadData_1[15:0] : writeDataVec_data_unreadData_5[15:0];
  wire [15:0]        writeDataVec_data_dataElement_6 = writeDataVec_data_dataIsRead_6 ? waiteReadData_2[15:0] : writeDataVec_data_unreadData_6[15:0];
  wire [15:0]        writeDataVec_data_dataElement_7 = writeDataVec_data_dataIsRead_7 ? waiteReadData_3[15:0] : writeDataVec_data_unreadData_7[15:0];
  wire [31:0]        writeDataVec_data_lo_1 = {writeDataVec_data_dataElement_5, writeDataVec_data_dataElement_4};
  wire [31:0]        writeDataVec_data_hi_1 = {writeDataVec_data_dataElement_7, writeDataVec_data_dataElement_6};
  wire [63:0]        writeDataVec_data_1 = {writeDataVec_data_hi_1, writeDataVec_data_lo_1};
  wire [190:0]       writeDataVec_shifterData_1 = {127'h0, writeDataVec_data_1} << {184'h0, executeIndexVec_1, 5'h0};
  wire [127:0]       writeDataVec_1 = writeDataVec_shifterData_1[127:0];
  wire [31:0]        writeDataVec_data_dataElement_8 = writeDataVec_data_dataIsRead_8 ? waiteReadData_0 : writeDataVec_data_unreadData_8;
  wire [31:0]        writeDataVec_data_dataElement_9 = writeDataVec_data_dataIsRead_9 ? waiteReadData_1 : writeDataVec_data_unreadData_9;
  wire [31:0]        writeDataVec_data_dataElement_10 = writeDataVec_data_dataIsRead_10 ? waiteReadData_2 : writeDataVec_data_unreadData_10;
  wire [31:0]        writeDataVec_data_dataElement_11 = writeDataVec_data_dataIsRead_11 ? waiteReadData_3 : writeDataVec_data_unreadData_11;
  wire [63:0]        writeDataVec_data_lo_2 = {writeDataVec_data_dataElement_9, writeDataVec_data_dataElement_8};
  wire [63:0]        writeDataVec_data_hi_2 = {writeDataVec_data_dataElement_11, writeDataVec_data_dataElement_10};
  wire [127:0]       writeDataVec_data_2 = {writeDataVec_data_hi_2, writeDataVec_data_lo_2};
  wire [190:0]       writeDataVec_shifterData_2 = {63'h0, writeDataVec_data_2};
  wire [127:0]       writeDataVec_2 = writeDataVec_shifterData_2[127:0];
  wire [127:0]       writeData = (sew1H[0] ? writeDataVec_0 : 128'h0) | (sew1H[1] ? writeDataVec_1 : 128'h0) | (sew1H[2] ? writeDataVec_2 : 128'h0);
  wire [1:0]         writeMaskVec_mask_lo = waiteReadDataPipeReg_sourceValid[1:0];
  wire [1:0]         writeMaskVec_mask_hi = waiteReadDataPipeReg_sourceValid[3:2];
  wire [3:0]         writeMaskVec_mask = {writeMaskVec_mask_hi, writeMaskVec_mask_lo};
  wire [18:0]        writeMaskVec_shifterMask = {15'h0, writeMaskVec_mask} << {15'h0, executeIndexVec_0, 2'h0};
  wire [15:0]        writeMaskVec_0 = writeMaskVec_shifterMask[15:0];
  wire [3:0]         writeMaskVec_mask_lo_1 = {{2{waiteReadDataPipeReg_sourceValid[1]}}, {2{waiteReadDataPipeReg_sourceValid[0]}}};
  wire [3:0]         writeMaskVec_mask_hi_1 = {{2{waiteReadDataPipeReg_sourceValid[3]}}, {2{waiteReadDataPipeReg_sourceValid[2]}}};
  wire [7:0]         writeMaskVec_mask_1 = {writeMaskVec_mask_hi_1, writeMaskVec_mask_lo_1};
  wire [22:0]        writeMaskVec_shifterMask_1 = {15'h0, writeMaskVec_mask_1} << {19'h0, executeIndexVec_1, 2'h0};
  wire [15:0]        writeMaskVec_1 = writeMaskVec_shifterMask_1[15:0];
  wire [7:0]         writeMaskVec_mask_lo_2 = {{4{waiteReadDataPipeReg_sourceValid[1]}}, {4{waiteReadDataPipeReg_sourceValid[0]}}};
  wire [7:0]         writeMaskVec_mask_hi_2 = {{4{waiteReadDataPipeReg_sourceValid[3]}}, {4{waiteReadDataPipeReg_sourceValid[2]}}};
  wire [15:0]        writeMaskVec_mask_2 = {writeMaskVec_mask_hi_2, writeMaskVec_mask_lo_2};
  wire [22:0]        writeMaskVec_shifterMask_2 = {7'h0, writeMaskVec_mask_2};
  wire [15:0]        writeMaskVec_2 = writeMaskVec_shifterMask_2[15:0];
  wire [15:0]        writeMask = (sew1H[0] ? writeMaskVec_0 : 16'h0) | (sew1H[1] ? writeMaskVec_1 : 16'h0) | (sew1H[2] ? writeMaskVec_2 : 16'h0);
  wire [14:0]        _writeRequest_res_writeData_groupCounter_T_6 = {3'h0, waiteReadDataPipeReg_executeGroup} << instReg_sew;
  wire [9:0]         writeRequest_0_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_6[11:2];
  wire [9:0]         writeRequest_1_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_6[11:2];
  wire [9:0]         writeRequest_2_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_6[11:2];
  wire [9:0]         writeRequest_3_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_6[11:2];
  wire [31:0]        writeRequest_0_writeData_data = writeData[31:0];
  wire [31:0]        writeRequest_1_writeData_data = writeData[63:32];
  wire [31:0]        writeRequest_2_writeData_data = writeData[95:64];
  wire [31:0]        writeRequest_3_writeData_data = writeData[127:96];
  wire [3:0]         writeRequest_0_writeData_mask = writeMask[3:0];
  wire [3:0]         writeRequest_1_writeData_mask = writeMask[7:4];
  wire [3:0]         writeRequest_2_writeData_mask = writeMask[11:8];
  wire [3:0]         writeRequest_3_writeData_mask = writeMask[15:12];
  wire [1:0]         WillWriteLane_lo = {|writeRequest_1_writeData_mask, |writeRequest_0_writeData_mask};
  wire [1:0]         WillWriteLane_hi = {|writeRequest_3_writeData_mask, |writeRequest_2_writeData_mask};
  wire [3:0]         WillWriteLane = {WillWriteLane_hi, WillWriteLane_lo};
  wire               waiteStageDeqValid = waiteReadStageValid & (waiteReadSate == waiteReadDataPipeReg_needRead | waiteReadDataPipeReg_needRead == 4'h0);
  wire               waiteStageDeqReady;
  wire               waiteStageDeqFire = waiteStageDeqValid & waiteStageDeqReady;
  assign waiteStageEnqReady = ~waiteReadStageValid | waiteStageDeqFire;
  assign readWaitQueue_deq_ready = waiteStageEnqReady;
  wire               waiteStageEnqFire = readWaitQueue_deq_valid & waiteStageEnqReady;
  wire               isWaiteForThisData = waiteReadDataPipeReg_needRead[0] & ~(waiteReadSate[0]) & waiteReadStageValid;
  assign readData_readDataQueue_deq_ready = isWaiteForThisData | unitType[2] | compress | gatherWaiteRead | mvRd;
  assign isWaiteForThisData_1 = waiteReadDataPipeReg_needRead[1] & ~(waiteReadSate[1]) & waiteReadStageValid;
  assign readData_readDataQueue_1_deq_ready = isWaiteForThisData_1;
  assign isWaiteForThisData_2 = waiteReadDataPipeReg_needRead[2] & ~(waiteReadSate[2]) & waiteReadStageValid;
  assign readData_readDataQueue_2_deq_ready = isWaiteForThisData_2;
  assign isWaiteForThisData_3 = waiteReadDataPipeReg_needRead[3] & ~(waiteReadSate[3]) & waiteReadStageValid;
  assign readData_readDataQueue_3_deq_ready = isWaiteForThisData_3;
  wire [1:0]         readResultValid_lo = {readTokenRelease_1, readTokenRelease_0};
  wire [1:0]         readResultValid_hi = {readTokenRelease_3, readTokenRelease_2};
  wire [3:0]         readResultValid = {readResultValid_hi, readResultValid_lo};
  wire               executeEnqValid = otherTypeRequestDeq & ~readType;
  wire [63:0]        source2_lo = {exeReqReg_1_bits_source2, exeReqReg_0_bits_source2};
  wire [63:0]        source2_hi = {exeReqReg_3_bits_source2, exeReqReg_2_bits_source2};
  wire [127:0]       source2 = {source2_hi, source2_lo};
  wire [127:0]       source1 = {source1_hi, source1_lo};
  wire               vs1Split_vs1SetIndex = requestCounter[0];
  wire               vs1Split_0_2 = vs1Split_vs1SetIndex;
  wire [1:0]         vs1Split_vs1SetIndex_1 = requestCounter[1:0];
  wire               vs1Split_1_2 = &vs1Split_vs1SetIndex_1;
  wire [2:0]         vs1Split_vs1SetIndex_2 = requestCounter[2:0];
  wire               vs1Split_2_2 = &vs1Split_vs1SetIndex_2;
  wire [15:0]        _compressSource1_T_3 = sew1H[0] ? (vs1Split_vs1SetIndex ? readVS1Reg_data[31:16] : readVS1Reg_data[15:0]) : 16'h0;
  wire [3:0][7:0]    _GEN_176 = {{readVS1Reg_data[31:24]}, {readVS1Reg_data[23:16]}, {readVS1Reg_data[15:8]}, {readVS1Reg_data[7:0]}};
  wire [7:0][3:0]    _GEN_180 = {{readVS1Reg_data[31:28]}, {readVS1Reg_data[27:24]}, {readVS1Reg_data[23:20]}, {readVS1Reg_data[19:16]}, {readVS1Reg_data[15:12]}, {readVS1Reg_data[11:8]}, {readVS1Reg_data[7:4]}, {readVS1Reg_data[3:0]}};
  wire [7:0]         _GEN_181 = _compressSource1_T_3[7:0] | (sew1H[1] ? _GEN_176[vs1Split_vs1SetIndex_1] : 8'h0);
  wire [15:0]        compressSource1 = {_compressSource1_T_3[15:8], _GEN_181[7:4], _GEN_181[3:0] | (sew1H[2] ? _GEN_180[vs1Split_vs1SetIndex_2] : 4'h0)};
  wire [31:0]        source1Select = mv ? readVS1Reg_data : {16'h0, compressSource1};
  wire               source1Change = sew1H[0] & vs1Split_0_2 | sew1H[1] & vs1Split_1_2 | sew1H[2] & vs1Split_2_2;
  assign viotaCounterAdd = executeEnqValid & unitType[1];
  wire [1:0]         view__in_bits_ffoInput_lo = {exeReqReg_1_bits_ffo, exeReqReg_0_bits_ffo};
  wire [1:0]         view__in_bits_ffoInput_hi = {exeReqReg_3_bits_ffo, exeReqReg_2_bits_ffo};
  wire               reduceUnit_in_valid = executeEnqValid & unitType[2];
  wire               _view__firstGroup_T_1 = _reduceUnit_in_ready & reduceUnit_in_valid;
  wire [11:0]        extendGroupCount = extendType ? (subType[2] ? _extendGroupCount_T_1 : {1'h0, requestCounter, executeIndex[1]}) : {2'h0, requestCounter};
  wire [127:0]       _executeResult_T_4 = unitType[1] ? compressUnitResultQueue_deq_bits_data : 128'h0;
  wire [127:0]       executeResult = {_executeResult_T_4[127:32], _executeResult_T_4[31:0] | (unitType[2] ? _reduceUnit_out_bits_data : 32'h0)} | (unitType[3] ? _extendUnit_out : 128'h0);
  assign executeReady = readType | unitType[1] | unitType[2] & _reduceUnit_in_ready & readVS1Reg_dataValid | unitType[3] & executeEnqValid;
  assign compressUnitResultQueue_deq_ready = &{compressUnitResultQueue_deq_ready_hi, compressUnitResultQueue_deq_ready_lo};
  wire               compressDeq = compressUnitResultQueue_deq_ready & compressUnitResultQueue_deq_valid;
  wire               executeValid = unitType[1] & compressDeq | unitType[3] & executeEnqValid;
  assign executeGroupCounter = (unitType[1] | unitType[2] ? requestCounter : 10'h0) | (unitType[3] ? extendGroupCount[9:0] : 10'h0);
  wire [11:0]        executeDeqGroupCounter = {2'h0, (unitType[1] ? compressUnitResultQueue_deq_bits_groupCounter : 10'h0) | (unitType[2] ? requestCounter : 10'h0)} | (unitType[3] ? extendGroupCount : 12'h0);
  wire [15:0]        executeWriteByteMask = compress | ffo | mvVd ? compressUnitResultQueue_deq_bits_mask : executeByteMask;
  wire               maskFilter = |{~maskDestinationType, currentMaskGroupForDestination[31:0]};
  wire               maskFilter_1 = |{~maskDestinationType, currentMaskGroupForDestination[63:32]};
  wire               maskFilter_2 = |{~maskDestinationType, currentMaskGroupForDestination[95:64]};
  wire               maskFilter_3 = |{~maskDestinationType, currentMaskGroupForDestination[127:96]};
  assign writeQueue_0_deq_valid = ~_writeQueue_fifo_empty;
  wire               exeResp_0_valid_0 = writeQueue_0_deq_valid;
  wire               writeQueue_dataOut_ffoByOther;
  wire [31:0]        writeQueue_dataOut_writeData_data;
  wire [31:0]        exeResp_0_bits_data_0 = writeQueue_0_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_writeData_mask;
  wire [3:0]         exeResp_0_bits_mask_0 = writeQueue_0_deq_bits_writeData_mask;
  wire [9:0]         writeQueue_dataOut_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_writeData_vd;
  wire [2:0]         writeQueue_dataOut_index;
  wire [9:0]         writeQueue_0_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_0_enq_bits_writeData_vd;
  wire [14:0]        writeQueue_dataIn_lo = {writeQueue_0_enq_bits_writeData_groupCounter, writeQueue_0_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_0_enq_bits_writeData_data;
  wire [3:0]         writeQueue_0_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi = {writeQueue_0_enq_bits_writeData_data, writeQueue_0_enq_bits_writeData_mask};
  wire               writeQueue_0_enq_bits_ffoByOther;
  wire [51:0]        writeQueue_dataIn_hi_1 = {writeQueue_0_enq_bits_ffoByOther, writeQueue_dataIn_hi, writeQueue_dataIn_lo};
  wire [54:0]        writeQueue_dataIn = {writeQueue_dataIn_hi_1, writeQueue_0_enq_bits_index};
  assign writeQueue_dataOut_index = _writeQueue_fifo_data_out[2:0];
  assign writeQueue_dataOut_writeData_vd = _writeQueue_fifo_data_out[7:3];
  assign writeQueue_dataOut_writeData_groupCounter = _writeQueue_fifo_data_out[17:8];
  assign writeQueue_dataOut_writeData_mask = _writeQueue_fifo_data_out[21:18];
  assign writeQueue_dataOut_writeData_data = _writeQueue_fifo_data_out[53:22];
  assign writeQueue_dataOut_ffoByOther = _writeQueue_fifo_data_out[54];
  wire               writeQueue_0_deq_bits_ffoByOther = writeQueue_dataOut_ffoByOther;
  assign writeQueue_0_deq_bits_writeData_data = writeQueue_dataOut_writeData_data;
  assign writeQueue_0_deq_bits_writeData_mask = writeQueue_dataOut_writeData_mask;
  wire [9:0]         writeQueue_0_deq_bits_writeData_groupCounter = writeQueue_dataOut_writeData_groupCounter;
  wire [4:0]         writeQueue_0_deq_bits_writeData_vd = writeQueue_dataOut_writeData_vd;
  wire [2:0]         writeQueue_0_deq_bits_index = writeQueue_dataOut_index;
  wire               writeQueue_0_enq_ready = ~_writeQueue_fifo_full;
  wire               writeQueue_0_enq_valid;
  assign writeQueue_1_deq_valid = ~_writeQueue_fifo_1_empty;
  wire               exeResp_1_valid_0 = writeQueue_1_deq_valid;
  wire               writeQueue_dataOut_1_ffoByOther;
  wire [31:0]        writeQueue_dataOut_1_writeData_data;
  wire [31:0]        exeResp_1_bits_data_0 = writeQueue_1_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_1_writeData_mask;
  wire [3:0]         exeResp_1_bits_mask_0 = writeQueue_1_deq_bits_writeData_mask;
  wire [9:0]         writeQueue_dataOut_1_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_1_writeData_vd;
  wire [2:0]         writeQueue_dataOut_1_index;
  wire [9:0]         writeQueue_1_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_1_enq_bits_writeData_vd;
  wire [14:0]        writeQueue_dataIn_lo_1 = {writeQueue_1_enq_bits_writeData_groupCounter, writeQueue_1_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_1_enq_bits_writeData_data;
  wire [3:0]         writeQueue_1_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_2 = {writeQueue_1_enq_bits_writeData_data, writeQueue_1_enq_bits_writeData_mask};
  wire               writeQueue_1_enq_bits_ffoByOther;
  wire [51:0]        writeQueue_dataIn_hi_3 = {writeQueue_1_enq_bits_ffoByOther, writeQueue_dataIn_hi_2, writeQueue_dataIn_lo_1};
  wire [54:0]        writeQueue_dataIn_1 = {writeQueue_dataIn_hi_3, writeQueue_1_enq_bits_index};
  assign writeQueue_dataOut_1_index = _writeQueue_fifo_1_data_out[2:0];
  assign writeQueue_dataOut_1_writeData_vd = _writeQueue_fifo_1_data_out[7:3];
  assign writeQueue_dataOut_1_writeData_groupCounter = _writeQueue_fifo_1_data_out[17:8];
  assign writeQueue_dataOut_1_writeData_mask = _writeQueue_fifo_1_data_out[21:18];
  assign writeQueue_dataOut_1_writeData_data = _writeQueue_fifo_1_data_out[53:22];
  assign writeQueue_dataOut_1_ffoByOther = _writeQueue_fifo_1_data_out[54];
  wire               writeQueue_1_deq_bits_ffoByOther = writeQueue_dataOut_1_ffoByOther;
  assign writeQueue_1_deq_bits_writeData_data = writeQueue_dataOut_1_writeData_data;
  assign writeQueue_1_deq_bits_writeData_mask = writeQueue_dataOut_1_writeData_mask;
  wire [9:0]         writeQueue_1_deq_bits_writeData_groupCounter = writeQueue_dataOut_1_writeData_groupCounter;
  wire [4:0]         writeQueue_1_deq_bits_writeData_vd = writeQueue_dataOut_1_writeData_vd;
  wire [2:0]         writeQueue_1_deq_bits_index = writeQueue_dataOut_1_index;
  wire               writeQueue_1_enq_ready = ~_writeQueue_fifo_1_full;
  wire               writeQueue_1_enq_valid;
  assign writeQueue_2_deq_valid = ~_writeQueue_fifo_2_empty;
  wire               exeResp_2_valid_0 = writeQueue_2_deq_valid;
  wire               writeQueue_dataOut_2_ffoByOther;
  wire [31:0]        writeQueue_dataOut_2_writeData_data;
  wire [31:0]        exeResp_2_bits_data_0 = writeQueue_2_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_2_writeData_mask;
  wire [3:0]         exeResp_2_bits_mask_0 = writeQueue_2_deq_bits_writeData_mask;
  wire [9:0]         writeQueue_dataOut_2_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_2_writeData_vd;
  wire [2:0]         writeQueue_dataOut_2_index;
  wire [9:0]         writeQueue_2_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_2_enq_bits_writeData_vd;
  wire [14:0]        writeQueue_dataIn_lo_2 = {writeQueue_2_enq_bits_writeData_groupCounter, writeQueue_2_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_2_enq_bits_writeData_data;
  wire [3:0]         writeQueue_2_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_4 = {writeQueue_2_enq_bits_writeData_data, writeQueue_2_enq_bits_writeData_mask};
  wire               writeQueue_2_enq_bits_ffoByOther;
  wire [51:0]        writeQueue_dataIn_hi_5 = {writeQueue_2_enq_bits_ffoByOther, writeQueue_dataIn_hi_4, writeQueue_dataIn_lo_2};
  wire [54:0]        writeQueue_dataIn_2 = {writeQueue_dataIn_hi_5, writeQueue_2_enq_bits_index};
  assign writeQueue_dataOut_2_index = _writeQueue_fifo_2_data_out[2:0];
  assign writeQueue_dataOut_2_writeData_vd = _writeQueue_fifo_2_data_out[7:3];
  assign writeQueue_dataOut_2_writeData_groupCounter = _writeQueue_fifo_2_data_out[17:8];
  assign writeQueue_dataOut_2_writeData_mask = _writeQueue_fifo_2_data_out[21:18];
  assign writeQueue_dataOut_2_writeData_data = _writeQueue_fifo_2_data_out[53:22];
  assign writeQueue_dataOut_2_ffoByOther = _writeQueue_fifo_2_data_out[54];
  wire               writeQueue_2_deq_bits_ffoByOther = writeQueue_dataOut_2_ffoByOther;
  assign writeQueue_2_deq_bits_writeData_data = writeQueue_dataOut_2_writeData_data;
  assign writeQueue_2_deq_bits_writeData_mask = writeQueue_dataOut_2_writeData_mask;
  wire [9:0]         writeQueue_2_deq_bits_writeData_groupCounter = writeQueue_dataOut_2_writeData_groupCounter;
  wire [4:0]         writeQueue_2_deq_bits_writeData_vd = writeQueue_dataOut_2_writeData_vd;
  wire [2:0]         writeQueue_2_deq_bits_index = writeQueue_dataOut_2_index;
  wire               writeQueue_2_enq_ready = ~_writeQueue_fifo_2_full;
  wire               writeQueue_2_enq_valid;
  assign writeQueue_3_deq_valid = ~_writeQueue_fifo_3_empty;
  wire               exeResp_3_valid_0 = writeQueue_3_deq_valid;
  wire               writeQueue_dataOut_3_ffoByOther;
  wire [31:0]        writeQueue_dataOut_3_writeData_data;
  wire [31:0]        exeResp_3_bits_data_0 = writeQueue_3_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_3_writeData_mask;
  wire [3:0]         exeResp_3_bits_mask_0 = writeQueue_3_deq_bits_writeData_mask;
  wire [9:0]         writeQueue_dataOut_3_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_3_writeData_vd;
  wire [2:0]         writeQueue_dataOut_3_index;
  wire [9:0]         writeQueue_3_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_3_enq_bits_writeData_vd;
  wire [14:0]        writeQueue_dataIn_lo_3 = {writeQueue_3_enq_bits_writeData_groupCounter, writeQueue_3_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_3_enq_bits_writeData_data;
  wire [3:0]         writeQueue_3_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_6 = {writeQueue_3_enq_bits_writeData_data, writeQueue_3_enq_bits_writeData_mask};
  wire               writeQueue_3_enq_bits_ffoByOther;
  wire [51:0]        writeQueue_dataIn_hi_7 = {writeQueue_3_enq_bits_ffoByOther, writeQueue_dataIn_hi_6, writeQueue_dataIn_lo_3};
  wire [54:0]        writeQueue_dataIn_3 = {writeQueue_dataIn_hi_7, writeQueue_3_enq_bits_index};
  assign writeQueue_dataOut_3_index = _writeQueue_fifo_3_data_out[2:0];
  assign writeQueue_dataOut_3_writeData_vd = _writeQueue_fifo_3_data_out[7:3];
  assign writeQueue_dataOut_3_writeData_groupCounter = _writeQueue_fifo_3_data_out[17:8];
  assign writeQueue_dataOut_3_writeData_mask = _writeQueue_fifo_3_data_out[21:18];
  assign writeQueue_dataOut_3_writeData_data = _writeQueue_fifo_3_data_out[53:22];
  assign writeQueue_dataOut_3_ffoByOther = _writeQueue_fifo_3_data_out[54];
  wire               writeQueue_3_deq_bits_ffoByOther = writeQueue_dataOut_3_ffoByOther;
  assign writeQueue_3_deq_bits_writeData_data = writeQueue_dataOut_3_writeData_data;
  assign writeQueue_3_deq_bits_writeData_mask = writeQueue_dataOut_3_writeData_mask;
  wire [9:0]         writeQueue_3_deq_bits_writeData_groupCounter = writeQueue_dataOut_3_writeData_groupCounter;
  wire [4:0]         writeQueue_3_deq_bits_writeData_vd = writeQueue_dataOut_3_writeData_vd;
  wire [2:0]         writeQueue_3_deq_bits_index = writeQueue_dataOut_3_index;
  wire               writeQueue_3_enq_ready = ~_writeQueue_fifo_3_full;
  wire               writeQueue_3_enq_valid;
  wire               dataNotInShifter_readTypeWriteVrf = waiteStageDeqFire & WillWriteLane[0];
  assign writeQueue_0_enq_valid = _maskedWrite_out_0_valid | dataNotInShifter_readTypeWriteVrf;
  assign writeQueue_0_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf ? writeRequest_0_writeData_vd : 5'h0;
  assign writeQueue_0_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf ? writeRequest_0_writeData_groupCounter : _maskedWrite_out_0_bits_writeData_groupCounter;
  assign writeQueue_0_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf ? writeRequest_0_writeData_mask : _maskedWrite_out_0_bits_writeData_mask;
  assign writeQueue_0_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf ? writeRequest_0_writeData_data : _maskedWrite_out_0_bits_writeData_data;
  assign writeQueue_0_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf & _maskedWrite_out_0_bits_ffoByOther;
  wire [4:0]         exeResp_0_bits_vd_0 = instReg_vd + {1'h0, writeQueue_0_deq_bits_writeData_groupCounter[9:6]};
  wire [5:0]         exeResp_0_bits_offset_0 = writeQueue_0_deq_bits_writeData_groupCounter[5:0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter;
  wire               _dataNotInShifter_T = exeResp_0_ready_0 & exeResp_0_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange = _dataNotInShifter_T ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_1 = waiteStageDeqFire & WillWriteLane[1];
  assign writeQueue_1_enq_valid = _maskedWrite_out_1_valid | dataNotInShifter_readTypeWriteVrf_1;
  assign writeQueue_1_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_1 ? writeRequest_1_writeData_vd : 5'h0;
  assign writeQueue_1_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_1 ? writeRequest_1_writeData_groupCounter : _maskedWrite_out_1_bits_writeData_groupCounter;
  assign writeQueue_1_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_1 ? writeRequest_1_writeData_mask : _maskedWrite_out_1_bits_writeData_mask;
  assign writeQueue_1_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_1 ? writeRequest_1_writeData_data : _maskedWrite_out_1_bits_writeData_data;
  assign writeQueue_1_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_1 & _maskedWrite_out_1_bits_ffoByOther;
  wire [4:0]         exeResp_1_bits_vd_0 = instReg_vd + {1'h0, writeQueue_1_deq_bits_writeData_groupCounter[9:6]};
  wire [5:0]         exeResp_1_bits_offset_0 = writeQueue_1_deq_bits_writeData_groupCounter[5:0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_1;
  wire               _dataNotInShifter_T_3 = exeResp_1_ready_0 & exeResp_1_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_1 = _dataNotInShifter_T_3 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_2 = waiteStageDeqFire & WillWriteLane[2];
  assign writeQueue_2_enq_valid = _maskedWrite_out_2_valid | dataNotInShifter_readTypeWriteVrf_2;
  assign writeQueue_2_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_2 ? writeRequest_2_writeData_vd : 5'h0;
  assign writeQueue_2_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_2 ? writeRequest_2_writeData_groupCounter : _maskedWrite_out_2_bits_writeData_groupCounter;
  assign writeQueue_2_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_2 ? writeRequest_2_writeData_mask : _maskedWrite_out_2_bits_writeData_mask;
  assign writeQueue_2_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_2 ? writeRequest_2_writeData_data : _maskedWrite_out_2_bits_writeData_data;
  assign writeQueue_2_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_2 & _maskedWrite_out_2_bits_ffoByOther;
  wire [4:0]         exeResp_2_bits_vd_0 = instReg_vd + {1'h0, writeQueue_2_deq_bits_writeData_groupCounter[9:6]};
  wire [5:0]         exeResp_2_bits_offset_0 = writeQueue_2_deq_bits_writeData_groupCounter[5:0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_2;
  wire               _dataNotInShifter_T_6 = exeResp_2_ready_0 & exeResp_2_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_2 = _dataNotInShifter_T_6 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_3 = waiteStageDeqFire & WillWriteLane[3];
  assign writeQueue_3_enq_valid = _maskedWrite_out_3_valid | dataNotInShifter_readTypeWriteVrf_3;
  assign writeQueue_3_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_3 ? writeRequest_3_writeData_vd : 5'h0;
  assign writeQueue_3_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_3 ? writeRequest_3_writeData_groupCounter : _maskedWrite_out_3_bits_writeData_groupCounter;
  assign writeQueue_3_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_3 ? writeRequest_3_writeData_mask : _maskedWrite_out_3_bits_writeData_mask;
  assign writeQueue_3_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_3 ? writeRequest_3_writeData_data : _maskedWrite_out_3_bits_writeData_data;
  assign writeQueue_3_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_3 & _maskedWrite_out_3_bits_ffoByOther;
  wire [4:0]         exeResp_3_bits_vd_0 = instReg_vd + {1'h0, writeQueue_3_deq_bits_writeData_groupCounter[9:6]};
  wire [5:0]         exeResp_3_bits_offset_0 = writeQueue_3_deq_bits_writeData_groupCounter[5:0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_3;
  wire               _dataNotInShifter_T_9 = exeResp_3_ready_0 & exeResp_3_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_3 = _dataNotInShifter_T_9 ? 3'h1 : 3'h7;
  wire               dataNotInShifter = dataNotInShifter_writeTokenCounter == 3'h0 & dataNotInShifter_writeTokenCounter_1 == 3'h0 & dataNotInShifter_writeTokenCounter_2 == 3'h0 & dataNotInShifter_writeTokenCounter_3 == 3'h0;
  assign waiteStageDeqReady = (~(WillWriteLane[0]) | writeQueue_0_enq_ready) & (~(WillWriteLane[1]) | writeQueue_1_enq_ready) & (~(WillWriteLane[2]) | writeQueue_2_enq_ready) & (~(WillWriteLane[3]) | writeQueue_3_enq_ready);
  reg                waiteLastRequest;
  reg                waitQueueClear;
  wire               lastReportValid = waitQueueClear & ~(writeQueue_0_deq_valid | writeQueue_1_deq_valid | writeQueue_2_deq_valid | writeQueue_3_deq_valid) & dataNotInShifter;
  wire               executeStageInvalid = unitType[1] & ~compressUnitResultQueue_deq_valid & ~_compressUnit_stageValid | unitType[2] & _reduceUnit_in_ready | unitType[3];
  wire               executeStageClean = readType ? waiteStageDeqFire & waiteReadDataPipeReg_last : waiteLastRequest & _maskedWrite_stageClear & executeStageInvalid;
  wire               invalidEnq = instReq_valid & instReq_bits_vl == 14'h0 & ~enqMvRD;
  wire [7:0]         _lastReport_output = lastReportValid ? 8'h1 << instReg_instructionIndex : 8'h0;
  wire [31:0]        gatherData_bits_0 = readVS1Reg_dataValid ? readVS1Reg_data : 32'h0;
  always @(posedge clock) begin
    if (reset) begin
      v0_0 <= 32'h0;
      v0_1 <= 32'h0;
      v0_2 <= 32'h0;
      v0_3 <= 32'h0;
      v0_4 <= 32'h0;
      v0_5 <= 32'h0;
      v0_6 <= 32'h0;
      v0_7 <= 32'h0;
      v0_8 <= 32'h0;
      v0_9 <= 32'h0;
      v0_10 <= 32'h0;
      v0_11 <= 32'h0;
      v0_12 <= 32'h0;
      v0_13 <= 32'h0;
      v0_14 <= 32'h0;
      v0_15 <= 32'h0;
      v0_16 <= 32'h0;
      v0_17 <= 32'h0;
      v0_18 <= 32'h0;
      v0_19 <= 32'h0;
      v0_20 <= 32'h0;
      v0_21 <= 32'h0;
      v0_22 <= 32'h0;
      v0_23 <= 32'h0;
      v0_24 <= 32'h0;
      v0_25 <= 32'h0;
      v0_26 <= 32'h0;
      v0_27 <= 32'h0;
      v0_28 <= 32'h0;
      v0_29 <= 32'h0;
      v0_30 <= 32'h0;
      v0_31 <= 32'h0;
      v0_32 <= 32'h0;
      v0_33 <= 32'h0;
      v0_34 <= 32'h0;
      v0_35 <= 32'h0;
      v0_36 <= 32'h0;
      v0_37 <= 32'h0;
      v0_38 <= 32'h0;
      v0_39 <= 32'h0;
      v0_40 <= 32'h0;
      v0_41 <= 32'h0;
      v0_42 <= 32'h0;
      v0_43 <= 32'h0;
      v0_44 <= 32'h0;
      v0_45 <= 32'h0;
      v0_46 <= 32'h0;
      v0_47 <= 32'h0;
      v0_48 <= 32'h0;
      v0_49 <= 32'h0;
      v0_50 <= 32'h0;
      v0_51 <= 32'h0;
      v0_52 <= 32'h0;
      v0_53 <= 32'h0;
      v0_54 <= 32'h0;
      v0_55 <= 32'h0;
      v0_56 <= 32'h0;
      v0_57 <= 32'h0;
      v0_58 <= 32'h0;
      v0_59 <= 32'h0;
      v0_60 <= 32'h0;
      v0_61 <= 32'h0;
      v0_62 <= 32'h0;
      v0_63 <= 32'h0;
      v0_64 <= 32'h0;
      v0_65 <= 32'h0;
      v0_66 <= 32'h0;
      v0_67 <= 32'h0;
      v0_68 <= 32'h0;
      v0_69 <= 32'h0;
      v0_70 <= 32'h0;
      v0_71 <= 32'h0;
      v0_72 <= 32'h0;
      v0_73 <= 32'h0;
      v0_74 <= 32'h0;
      v0_75 <= 32'h0;
      v0_76 <= 32'h0;
      v0_77 <= 32'h0;
      v0_78 <= 32'h0;
      v0_79 <= 32'h0;
      v0_80 <= 32'h0;
      v0_81 <= 32'h0;
      v0_82 <= 32'h0;
      v0_83 <= 32'h0;
      v0_84 <= 32'h0;
      v0_85 <= 32'h0;
      v0_86 <= 32'h0;
      v0_87 <= 32'h0;
      v0_88 <= 32'h0;
      v0_89 <= 32'h0;
      v0_90 <= 32'h0;
      v0_91 <= 32'h0;
      v0_92 <= 32'h0;
      v0_93 <= 32'h0;
      v0_94 <= 32'h0;
      v0_95 <= 32'h0;
      v0_96 <= 32'h0;
      v0_97 <= 32'h0;
      v0_98 <= 32'h0;
      v0_99 <= 32'h0;
      v0_100 <= 32'h0;
      v0_101 <= 32'h0;
      v0_102 <= 32'h0;
      v0_103 <= 32'h0;
      v0_104 <= 32'h0;
      v0_105 <= 32'h0;
      v0_106 <= 32'h0;
      v0_107 <= 32'h0;
      v0_108 <= 32'h0;
      v0_109 <= 32'h0;
      v0_110 <= 32'h0;
      v0_111 <= 32'h0;
      v0_112 <= 32'h0;
      v0_113 <= 32'h0;
      v0_114 <= 32'h0;
      v0_115 <= 32'h0;
      v0_116 <= 32'h0;
      v0_117 <= 32'h0;
      v0_118 <= 32'h0;
      v0_119 <= 32'h0;
      v0_120 <= 32'h0;
      v0_121 <= 32'h0;
      v0_122 <= 32'h0;
      v0_123 <= 32'h0;
      v0_124 <= 32'h0;
      v0_125 <= 32'h0;
      v0_126 <= 32'h0;
      v0_127 <= 32'h0;
      v0_128 <= 32'h0;
      v0_129 <= 32'h0;
      v0_130 <= 32'h0;
      v0_131 <= 32'h0;
      v0_132 <= 32'h0;
      v0_133 <= 32'h0;
      v0_134 <= 32'h0;
      v0_135 <= 32'h0;
      v0_136 <= 32'h0;
      v0_137 <= 32'h0;
      v0_138 <= 32'h0;
      v0_139 <= 32'h0;
      v0_140 <= 32'h0;
      v0_141 <= 32'h0;
      v0_142 <= 32'h0;
      v0_143 <= 32'h0;
      v0_144 <= 32'h0;
      v0_145 <= 32'h0;
      v0_146 <= 32'h0;
      v0_147 <= 32'h0;
      v0_148 <= 32'h0;
      v0_149 <= 32'h0;
      v0_150 <= 32'h0;
      v0_151 <= 32'h0;
      v0_152 <= 32'h0;
      v0_153 <= 32'h0;
      v0_154 <= 32'h0;
      v0_155 <= 32'h0;
      v0_156 <= 32'h0;
      v0_157 <= 32'h0;
      v0_158 <= 32'h0;
      v0_159 <= 32'h0;
      v0_160 <= 32'h0;
      v0_161 <= 32'h0;
      v0_162 <= 32'h0;
      v0_163 <= 32'h0;
      v0_164 <= 32'h0;
      v0_165 <= 32'h0;
      v0_166 <= 32'h0;
      v0_167 <= 32'h0;
      v0_168 <= 32'h0;
      v0_169 <= 32'h0;
      v0_170 <= 32'h0;
      v0_171 <= 32'h0;
      v0_172 <= 32'h0;
      v0_173 <= 32'h0;
      v0_174 <= 32'h0;
      v0_175 <= 32'h0;
      v0_176 <= 32'h0;
      v0_177 <= 32'h0;
      v0_178 <= 32'h0;
      v0_179 <= 32'h0;
      v0_180 <= 32'h0;
      v0_181 <= 32'h0;
      v0_182 <= 32'h0;
      v0_183 <= 32'h0;
      v0_184 <= 32'h0;
      v0_185 <= 32'h0;
      v0_186 <= 32'h0;
      v0_187 <= 32'h0;
      v0_188 <= 32'h0;
      v0_189 <= 32'h0;
      v0_190 <= 32'h0;
      v0_191 <= 32'h0;
      v0_192 <= 32'h0;
      v0_193 <= 32'h0;
      v0_194 <= 32'h0;
      v0_195 <= 32'h0;
      v0_196 <= 32'h0;
      v0_197 <= 32'h0;
      v0_198 <= 32'h0;
      v0_199 <= 32'h0;
      v0_200 <= 32'h0;
      v0_201 <= 32'h0;
      v0_202 <= 32'h0;
      v0_203 <= 32'h0;
      v0_204 <= 32'h0;
      v0_205 <= 32'h0;
      v0_206 <= 32'h0;
      v0_207 <= 32'h0;
      v0_208 <= 32'h0;
      v0_209 <= 32'h0;
      v0_210 <= 32'h0;
      v0_211 <= 32'h0;
      v0_212 <= 32'h0;
      v0_213 <= 32'h0;
      v0_214 <= 32'h0;
      v0_215 <= 32'h0;
      v0_216 <= 32'h0;
      v0_217 <= 32'h0;
      v0_218 <= 32'h0;
      v0_219 <= 32'h0;
      v0_220 <= 32'h0;
      v0_221 <= 32'h0;
      v0_222 <= 32'h0;
      v0_223 <= 32'h0;
      v0_224 <= 32'h0;
      v0_225 <= 32'h0;
      v0_226 <= 32'h0;
      v0_227 <= 32'h0;
      v0_228 <= 32'h0;
      v0_229 <= 32'h0;
      v0_230 <= 32'h0;
      v0_231 <= 32'h0;
      v0_232 <= 32'h0;
      v0_233 <= 32'h0;
      v0_234 <= 32'h0;
      v0_235 <= 32'h0;
      v0_236 <= 32'h0;
      v0_237 <= 32'h0;
      v0_238 <= 32'h0;
      v0_239 <= 32'h0;
      v0_240 <= 32'h0;
      v0_241 <= 32'h0;
      v0_242 <= 32'h0;
      v0_243 <= 32'h0;
      v0_244 <= 32'h0;
      v0_245 <= 32'h0;
      v0_246 <= 32'h0;
      v0_247 <= 32'h0;
      v0_248 <= 32'h0;
      v0_249 <= 32'h0;
      v0_250 <= 32'h0;
      v0_251 <= 32'h0;
      v0_252 <= 32'h0;
      v0_253 <= 32'h0;
      v0_254 <= 32'h0;
      v0_255 <= 32'h0;
      gatherReadState <= 2'h0;
      gatherDatOffset <= 2'h0;
      gatherLane <= 2'h0;
      gatherOffset <= 6'h0;
      gatherGrowth <= 3'h0;
      instReg_instructionIndex <= 3'h0;
      instReg_decodeResult_specialSlot <= 1'h0;
      instReg_decodeResult_topUop <= 5'h0;
      instReg_decodeResult_popCount <= 1'h0;
      instReg_decodeResult_ffo <= 1'h0;
      instReg_decodeResult_average <= 1'h0;
      instReg_decodeResult_reverse <= 1'h0;
      instReg_decodeResult_dontNeedExecuteInLane <= 1'h0;
      instReg_decodeResult_scheduler <= 1'h0;
      instReg_decodeResult_sReadVD <= 1'h0;
      instReg_decodeResult_vtype <= 1'h0;
      instReg_decodeResult_sWrite <= 1'h0;
      instReg_decodeResult_crossRead <= 1'h0;
      instReg_decodeResult_crossWrite <= 1'h0;
      instReg_decodeResult_maskUnit <= 1'h0;
      instReg_decodeResult_special <= 1'h0;
      instReg_decodeResult_saturate <= 1'h0;
      instReg_decodeResult_vwmacc <= 1'h0;
      instReg_decodeResult_readOnly <= 1'h0;
      instReg_decodeResult_maskSource <= 1'h0;
      instReg_decodeResult_maskDestination <= 1'h0;
      instReg_decodeResult_maskLogic <= 1'h0;
      instReg_decodeResult_uop <= 4'h0;
      instReg_decodeResult_iota <= 1'h0;
      instReg_decodeResult_mv <= 1'h0;
      instReg_decodeResult_extend <= 1'h0;
      instReg_decodeResult_unOrderWrite <= 1'h0;
      instReg_decodeResult_compress <= 1'h0;
      instReg_decodeResult_gather16 <= 1'h0;
      instReg_decodeResult_gather <= 1'h0;
      instReg_decodeResult_slid <= 1'h0;
      instReg_decodeResult_targetRd <= 1'h0;
      instReg_decodeResult_widenReduce <= 1'h0;
      instReg_decodeResult_red <= 1'h0;
      instReg_decodeResult_nr <= 1'h0;
      instReg_decodeResult_itype <= 1'h0;
      instReg_decodeResult_unsigned1 <= 1'h0;
      instReg_decodeResult_unsigned0 <= 1'h0;
      instReg_decodeResult_other <= 1'h0;
      instReg_decodeResult_multiCycle <= 1'h0;
      instReg_decodeResult_divider <= 1'h0;
      instReg_decodeResult_multiplier <= 1'h0;
      instReg_decodeResult_shift <= 1'h0;
      instReg_decodeResult_adder <= 1'h0;
      instReg_decodeResult_logic <= 1'h0;
      instReg_readFromScala <= 32'h0;
      instReg_sew <= 2'h0;
      instReg_vlmul <= 3'h0;
      instReg_maskType <= 1'h0;
      instReg_vxrm <= 3'h0;
      instReg_vs2 <= 5'h0;
      instReg_vs1 <= 5'h0;
      instReg_vd <= 5'h0;
      instReg_vl <= 14'h0;
      instVlValid <= 1'h0;
      readVS1Reg_dataValid <= 1'h0;
      readVS1Reg_requestSend <= 1'h0;
      readVS1Reg_sendToExecution <= 1'h0;
      readVS1Reg_data <= 32'h0;
      readVS1Reg_readIndex <= 9'h0;
      exeReqReg_0_valid <= 1'h0;
      exeReqReg_0_bits_source1 <= 32'h0;
      exeReqReg_0_bits_source2 <= 32'h0;
      exeReqReg_0_bits_index <= 3'h0;
      exeReqReg_0_bits_ffo <= 1'h0;
      exeReqReg_1_valid <= 1'h0;
      exeReqReg_1_bits_source1 <= 32'h0;
      exeReqReg_1_bits_source2 <= 32'h0;
      exeReqReg_1_bits_index <= 3'h0;
      exeReqReg_1_bits_ffo <= 1'h0;
      exeReqReg_2_valid <= 1'h0;
      exeReqReg_2_bits_source1 <= 32'h0;
      exeReqReg_2_bits_source2 <= 32'h0;
      exeReqReg_2_bits_index <= 3'h0;
      exeReqReg_2_bits_ffo <= 1'h0;
      exeReqReg_3_valid <= 1'h0;
      exeReqReg_3_bits_source1 <= 32'h0;
      exeReqReg_3_bits_source2 <= 32'h0;
      exeReqReg_3_bits_index <= 3'h0;
      exeReqReg_3_bits_ffo <= 1'h0;
      requestCounter <= 10'h0;
      executeIndex <= 2'h0;
      readIssueStageState_groupReadState <= 4'h0;
      readIssueStageState_needRead <= 4'h0;
      readIssueStageState_elementValid <= 4'h0;
      readIssueStageState_replaceVs1 <= 4'h0;
      readIssueStageState_readOffset <= 24'h0;
      readIssueStageState_accessLane_0 <= 2'h0;
      readIssueStageState_accessLane_1 <= 2'h0;
      readIssueStageState_accessLane_2 <= 2'h0;
      readIssueStageState_accessLane_3 <= 2'h0;
      readIssueStageState_vsGrowth_0 <= 3'h0;
      readIssueStageState_vsGrowth_1 <= 3'h0;
      readIssueStageState_vsGrowth_2 <= 3'h0;
      readIssueStageState_vsGrowth_3 <= 3'h0;
      readIssueStageState_executeGroup <= 12'h0;
      readIssueStageState_readDataOffset <= 8'h0;
      readIssueStageState_last <= 1'h0;
      readIssueStageValid <= 1'h0;
      tokenCheck_counter <= 4'h0;
      tokenCheck_counter_1 <= 4'h0;
      tokenCheck_counter_2 <= 4'h0;
      tokenCheck_counter_3 <= 4'h0;
      reorderQueueAllocate_counter <= 4'h0;
      reorderQueueAllocate_counterWillUpdate <= 4'h0;
      reorderQueueAllocate_counter_1 <= 4'h0;
      reorderQueueAllocate_counterWillUpdate_1 <= 4'h0;
      reorderQueueAllocate_counter_2 <= 4'h0;
      reorderQueueAllocate_counterWillUpdate_2 <= 4'h0;
      reorderQueueAllocate_counter_3 <= 4'h0;
      reorderQueueAllocate_counterWillUpdate_3 <= 4'h0;
      reorderStageValid <= 1'h0;
      reorderStageState_0 <= 3'h0;
      reorderStageState_1 <= 3'h0;
      reorderStageState_2 <= 3'h0;
      reorderStageState_3 <= 3'h0;
      reorderStageNeed_0 <= 3'h0;
      reorderStageNeed_1 <= 3'h0;
      reorderStageNeed_2 <= 3'h0;
      reorderStageNeed_3 <= 3'h0;
      waiteReadDataPipeReg_executeGroup <= 12'h0;
      waiteReadDataPipeReg_sourceValid <= 4'h0;
      waiteReadDataPipeReg_replaceVs1 <= 4'h0;
      waiteReadDataPipeReg_needRead <= 4'h0;
      waiteReadDataPipeReg_last <= 1'h0;
      waiteReadData_0 <= 32'h0;
      waiteReadData_1 <= 32'h0;
      waiteReadData_2 <= 32'h0;
      waiteReadData_3 <= 32'h0;
      waiteReadSate <= 4'h0;
      waiteReadStageValid <= 1'h0;
      dataNotInShifter_writeTokenCounter <= 3'h0;
      dataNotInShifter_writeTokenCounter_1 <= 3'h0;
      dataNotInShifter_writeTokenCounter_2 <= 3'h0;
      dataNotInShifter_writeTokenCounter_3 <= 3'h0;
      waiteLastRequest <= 1'h0;
      waitQueueClear <= 1'h0;
    end
    else begin
      automatic logic _GEN_177 = instReq_valid & (viotaReq | enqMvRD) | gatherRequestFire;
      automatic logic _GEN_178;
      automatic logic _GEN_179 = source1Change & viotaCounterAdd;
      _GEN_178 = instReq_valid | gatherRequestFire;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h0)
        v0_0 <= v0_0 & ~maskExt | maskExt & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h0)
        v0_1 <= v0_1 & ~maskExt_1 | maskExt_1 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h0)
        v0_2 <= v0_2 & ~maskExt_2 | maskExt_2 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h0)
        v0_3 <= v0_3 & ~maskExt_3 | maskExt_3 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h1)
        v0_4 <= v0_4 & ~maskExt_4 | maskExt_4 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h1)
        v0_5 <= v0_5 & ~maskExt_5 | maskExt_5 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h1)
        v0_6 <= v0_6 & ~maskExt_6 | maskExt_6 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h1)
        v0_7 <= v0_7 & ~maskExt_7 | maskExt_7 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h2)
        v0_8 <= v0_8 & ~maskExt_8 | maskExt_8 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h2)
        v0_9 <= v0_9 & ~maskExt_9 | maskExt_9 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h2)
        v0_10 <= v0_10 & ~maskExt_10 | maskExt_10 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h2)
        v0_11 <= v0_11 & ~maskExt_11 | maskExt_11 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h3)
        v0_12 <= v0_12 & ~maskExt_12 | maskExt_12 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h3)
        v0_13 <= v0_13 & ~maskExt_13 | maskExt_13 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h3)
        v0_14 <= v0_14 & ~maskExt_14 | maskExt_14 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h3)
        v0_15 <= v0_15 & ~maskExt_15 | maskExt_15 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h4)
        v0_16 <= v0_16 & ~maskExt_16 | maskExt_16 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h4)
        v0_17 <= v0_17 & ~maskExt_17 | maskExt_17 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h4)
        v0_18 <= v0_18 & ~maskExt_18 | maskExt_18 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h4)
        v0_19 <= v0_19 & ~maskExt_19 | maskExt_19 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h5)
        v0_20 <= v0_20 & ~maskExt_20 | maskExt_20 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h5)
        v0_21 <= v0_21 & ~maskExt_21 | maskExt_21 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h5)
        v0_22 <= v0_22 & ~maskExt_22 | maskExt_22 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h5)
        v0_23 <= v0_23 & ~maskExt_23 | maskExt_23 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h6)
        v0_24 <= v0_24 & ~maskExt_24 | maskExt_24 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h6)
        v0_25 <= v0_25 & ~maskExt_25 | maskExt_25 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h6)
        v0_26 <= v0_26 & ~maskExt_26 | maskExt_26 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h6)
        v0_27 <= v0_27 & ~maskExt_27 | maskExt_27 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h7)
        v0_28 <= v0_28 & ~maskExt_28 | maskExt_28 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h7)
        v0_29 <= v0_29 & ~maskExt_29 | maskExt_29 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h7)
        v0_30 <= v0_30 & ~maskExt_30 | maskExt_30 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h7)
        v0_31 <= v0_31 & ~maskExt_31 | maskExt_31 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h8)
        v0_32 <= v0_32 & ~maskExt_32 | maskExt_32 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h8)
        v0_33 <= v0_33 & ~maskExt_33 | maskExt_33 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h8)
        v0_34 <= v0_34 & ~maskExt_34 | maskExt_34 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h8)
        v0_35 <= v0_35 & ~maskExt_35 | maskExt_35 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h9)
        v0_36 <= v0_36 & ~maskExt_36 | maskExt_36 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h9)
        v0_37 <= v0_37 & ~maskExt_37 | maskExt_37 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h9)
        v0_38 <= v0_38 & ~maskExt_38 | maskExt_38 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h9)
        v0_39 <= v0_39 & ~maskExt_39 | maskExt_39 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'hA)
        v0_40 <= v0_40 & ~maskExt_40 | maskExt_40 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'hA)
        v0_41 <= v0_41 & ~maskExt_41 | maskExt_41 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'hA)
        v0_42 <= v0_42 & ~maskExt_42 | maskExt_42 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'hA)
        v0_43 <= v0_43 & ~maskExt_43 | maskExt_43 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'hB)
        v0_44 <= v0_44 & ~maskExt_44 | maskExt_44 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'hB)
        v0_45 <= v0_45 & ~maskExt_45 | maskExt_45 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'hB)
        v0_46 <= v0_46 & ~maskExt_46 | maskExt_46 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'hB)
        v0_47 <= v0_47 & ~maskExt_47 | maskExt_47 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'hC)
        v0_48 <= v0_48 & ~maskExt_48 | maskExt_48 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'hC)
        v0_49 <= v0_49 & ~maskExt_49 | maskExt_49 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'hC)
        v0_50 <= v0_50 & ~maskExt_50 | maskExt_50 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'hC)
        v0_51 <= v0_51 & ~maskExt_51 | maskExt_51 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'hD)
        v0_52 <= v0_52 & ~maskExt_52 | maskExt_52 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'hD)
        v0_53 <= v0_53 & ~maskExt_53 | maskExt_53 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'hD)
        v0_54 <= v0_54 & ~maskExt_54 | maskExt_54 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'hD)
        v0_55 <= v0_55 & ~maskExt_55 | maskExt_55 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'hE)
        v0_56 <= v0_56 & ~maskExt_56 | maskExt_56 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'hE)
        v0_57 <= v0_57 & ~maskExt_57 | maskExt_57 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'hE)
        v0_58 <= v0_58 & ~maskExt_58 | maskExt_58 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'hE)
        v0_59 <= v0_59 & ~maskExt_59 | maskExt_59 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'hF)
        v0_60 <= v0_60 & ~maskExt_60 | maskExt_60 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'hF)
        v0_61 <= v0_61 & ~maskExt_61 | maskExt_61 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'hF)
        v0_62 <= v0_62 & ~maskExt_62 | maskExt_62 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'hF)
        v0_63 <= v0_63 & ~maskExt_63 | maskExt_63 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h10)
        v0_64 <= v0_64 & ~maskExt_64 | maskExt_64 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h10)
        v0_65 <= v0_65 & ~maskExt_65 | maskExt_65 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h10)
        v0_66 <= v0_66 & ~maskExt_66 | maskExt_66 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h10)
        v0_67 <= v0_67 & ~maskExt_67 | maskExt_67 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h11)
        v0_68 <= v0_68 & ~maskExt_68 | maskExt_68 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h11)
        v0_69 <= v0_69 & ~maskExt_69 | maskExt_69 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h11)
        v0_70 <= v0_70 & ~maskExt_70 | maskExt_70 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h11)
        v0_71 <= v0_71 & ~maskExt_71 | maskExt_71 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h12)
        v0_72 <= v0_72 & ~maskExt_72 | maskExt_72 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h12)
        v0_73 <= v0_73 & ~maskExt_73 | maskExt_73 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h12)
        v0_74 <= v0_74 & ~maskExt_74 | maskExt_74 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h12)
        v0_75 <= v0_75 & ~maskExt_75 | maskExt_75 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h13)
        v0_76 <= v0_76 & ~maskExt_76 | maskExt_76 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h13)
        v0_77 <= v0_77 & ~maskExt_77 | maskExt_77 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h13)
        v0_78 <= v0_78 & ~maskExt_78 | maskExt_78 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h13)
        v0_79 <= v0_79 & ~maskExt_79 | maskExt_79 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h14)
        v0_80 <= v0_80 & ~maskExt_80 | maskExt_80 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h14)
        v0_81 <= v0_81 & ~maskExt_81 | maskExt_81 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h14)
        v0_82 <= v0_82 & ~maskExt_82 | maskExt_82 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h14)
        v0_83 <= v0_83 & ~maskExt_83 | maskExt_83 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h15)
        v0_84 <= v0_84 & ~maskExt_84 | maskExt_84 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h15)
        v0_85 <= v0_85 & ~maskExt_85 | maskExt_85 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h15)
        v0_86 <= v0_86 & ~maskExt_86 | maskExt_86 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h15)
        v0_87 <= v0_87 & ~maskExt_87 | maskExt_87 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h16)
        v0_88 <= v0_88 & ~maskExt_88 | maskExt_88 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h16)
        v0_89 <= v0_89 & ~maskExt_89 | maskExt_89 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h16)
        v0_90 <= v0_90 & ~maskExt_90 | maskExt_90 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h16)
        v0_91 <= v0_91 & ~maskExt_91 | maskExt_91 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h17)
        v0_92 <= v0_92 & ~maskExt_92 | maskExt_92 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h17)
        v0_93 <= v0_93 & ~maskExt_93 | maskExt_93 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h17)
        v0_94 <= v0_94 & ~maskExt_94 | maskExt_94 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h17)
        v0_95 <= v0_95 & ~maskExt_95 | maskExt_95 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h18)
        v0_96 <= v0_96 & ~maskExt_96 | maskExt_96 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h18)
        v0_97 <= v0_97 & ~maskExt_97 | maskExt_97 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h18)
        v0_98 <= v0_98 & ~maskExt_98 | maskExt_98 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h18)
        v0_99 <= v0_99 & ~maskExt_99 | maskExt_99 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h19)
        v0_100 <= v0_100 & ~maskExt_100 | maskExt_100 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h19)
        v0_101 <= v0_101 & ~maskExt_101 | maskExt_101 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h19)
        v0_102 <= v0_102 & ~maskExt_102 | maskExt_102 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h19)
        v0_103 <= v0_103 & ~maskExt_103 | maskExt_103 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h1A)
        v0_104 <= v0_104 & ~maskExt_104 | maskExt_104 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h1A)
        v0_105 <= v0_105 & ~maskExt_105 | maskExt_105 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h1A)
        v0_106 <= v0_106 & ~maskExt_106 | maskExt_106 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h1A)
        v0_107 <= v0_107 & ~maskExt_107 | maskExt_107 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h1B)
        v0_108 <= v0_108 & ~maskExt_108 | maskExt_108 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h1B)
        v0_109 <= v0_109 & ~maskExt_109 | maskExt_109 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h1B)
        v0_110 <= v0_110 & ~maskExt_110 | maskExt_110 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h1B)
        v0_111 <= v0_111 & ~maskExt_111 | maskExt_111 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h1C)
        v0_112 <= v0_112 & ~maskExt_112 | maskExt_112 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h1C)
        v0_113 <= v0_113 & ~maskExt_113 | maskExt_113 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h1C)
        v0_114 <= v0_114 & ~maskExt_114 | maskExt_114 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h1C)
        v0_115 <= v0_115 & ~maskExt_115 | maskExt_115 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h1D)
        v0_116 <= v0_116 & ~maskExt_116 | maskExt_116 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h1D)
        v0_117 <= v0_117 & ~maskExt_117 | maskExt_117 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h1D)
        v0_118 <= v0_118 & ~maskExt_118 | maskExt_118 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h1D)
        v0_119 <= v0_119 & ~maskExt_119 | maskExt_119 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h1E)
        v0_120 <= v0_120 & ~maskExt_120 | maskExt_120 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h1E)
        v0_121 <= v0_121 & ~maskExt_121 | maskExt_121 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h1E)
        v0_122 <= v0_122 & ~maskExt_122 | maskExt_122 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h1E)
        v0_123 <= v0_123 & ~maskExt_123 | maskExt_123 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h1F)
        v0_124 <= v0_124 & ~maskExt_124 | maskExt_124 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h1F)
        v0_125 <= v0_125 & ~maskExt_125 | maskExt_125 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h1F)
        v0_126 <= v0_126 & ~maskExt_126 | maskExt_126 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h1F)
        v0_127 <= v0_127 & ~maskExt_127 | maskExt_127 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h20)
        v0_128 <= v0_128 & ~maskExt_128 | maskExt_128 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h20)
        v0_129 <= v0_129 & ~maskExt_129 | maskExt_129 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h20)
        v0_130 <= v0_130 & ~maskExt_130 | maskExt_130 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h20)
        v0_131 <= v0_131 & ~maskExt_131 | maskExt_131 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h21)
        v0_132 <= v0_132 & ~maskExt_132 | maskExt_132 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h21)
        v0_133 <= v0_133 & ~maskExt_133 | maskExt_133 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h21)
        v0_134 <= v0_134 & ~maskExt_134 | maskExt_134 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h21)
        v0_135 <= v0_135 & ~maskExt_135 | maskExt_135 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h22)
        v0_136 <= v0_136 & ~maskExt_136 | maskExt_136 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h22)
        v0_137 <= v0_137 & ~maskExt_137 | maskExt_137 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h22)
        v0_138 <= v0_138 & ~maskExt_138 | maskExt_138 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h22)
        v0_139 <= v0_139 & ~maskExt_139 | maskExt_139 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h23)
        v0_140 <= v0_140 & ~maskExt_140 | maskExt_140 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h23)
        v0_141 <= v0_141 & ~maskExt_141 | maskExt_141 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h23)
        v0_142 <= v0_142 & ~maskExt_142 | maskExt_142 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h23)
        v0_143 <= v0_143 & ~maskExt_143 | maskExt_143 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h24)
        v0_144 <= v0_144 & ~maskExt_144 | maskExt_144 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h24)
        v0_145 <= v0_145 & ~maskExt_145 | maskExt_145 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h24)
        v0_146 <= v0_146 & ~maskExt_146 | maskExt_146 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h24)
        v0_147 <= v0_147 & ~maskExt_147 | maskExt_147 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h25)
        v0_148 <= v0_148 & ~maskExt_148 | maskExt_148 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h25)
        v0_149 <= v0_149 & ~maskExt_149 | maskExt_149 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h25)
        v0_150 <= v0_150 & ~maskExt_150 | maskExt_150 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h25)
        v0_151 <= v0_151 & ~maskExt_151 | maskExt_151 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h26)
        v0_152 <= v0_152 & ~maskExt_152 | maskExt_152 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h26)
        v0_153 <= v0_153 & ~maskExt_153 | maskExt_153 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h26)
        v0_154 <= v0_154 & ~maskExt_154 | maskExt_154 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h26)
        v0_155 <= v0_155 & ~maskExt_155 | maskExt_155 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h27)
        v0_156 <= v0_156 & ~maskExt_156 | maskExt_156 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h27)
        v0_157 <= v0_157 & ~maskExt_157 | maskExt_157 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h27)
        v0_158 <= v0_158 & ~maskExt_158 | maskExt_158 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h27)
        v0_159 <= v0_159 & ~maskExt_159 | maskExt_159 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h28)
        v0_160 <= v0_160 & ~maskExt_160 | maskExt_160 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h28)
        v0_161 <= v0_161 & ~maskExt_161 | maskExt_161 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h28)
        v0_162 <= v0_162 & ~maskExt_162 | maskExt_162 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h28)
        v0_163 <= v0_163 & ~maskExt_163 | maskExt_163 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h29)
        v0_164 <= v0_164 & ~maskExt_164 | maskExt_164 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h29)
        v0_165 <= v0_165 & ~maskExt_165 | maskExt_165 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h29)
        v0_166 <= v0_166 & ~maskExt_166 | maskExt_166 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h29)
        v0_167 <= v0_167 & ~maskExt_167 | maskExt_167 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h2A)
        v0_168 <= v0_168 & ~maskExt_168 | maskExt_168 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h2A)
        v0_169 <= v0_169 & ~maskExt_169 | maskExt_169 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h2A)
        v0_170 <= v0_170 & ~maskExt_170 | maskExt_170 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h2A)
        v0_171 <= v0_171 & ~maskExt_171 | maskExt_171 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h2B)
        v0_172 <= v0_172 & ~maskExt_172 | maskExt_172 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h2B)
        v0_173 <= v0_173 & ~maskExt_173 | maskExt_173 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h2B)
        v0_174 <= v0_174 & ~maskExt_174 | maskExt_174 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h2B)
        v0_175 <= v0_175 & ~maskExt_175 | maskExt_175 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h2C)
        v0_176 <= v0_176 & ~maskExt_176 | maskExt_176 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h2C)
        v0_177 <= v0_177 & ~maskExt_177 | maskExt_177 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h2C)
        v0_178 <= v0_178 & ~maskExt_178 | maskExt_178 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h2C)
        v0_179 <= v0_179 & ~maskExt_179 | maskExt_179 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h2D)
        v0_180 <= v0_180 & ~maskExt_180 | maskExt_180 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h2D)
        v0_181 <= v0_181 & ~maskExt_181 | maskExt_181 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h2D)
        v0_182 <= v0_182 & ~maskExt_182 | maskExt_182 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h2D)
        v0_183 <= v0_183 & ~maskExt_183 | maskExt_183 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h2E)
        v0_184 <= v0_184 & ~maskExt_184 | maskExt_184 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h2E)
        v0_185 <= v0_185 & ~maskExt_185 | maskExt_185 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h2E)
        v0_186 <= v0_186 & ~maskExt_186 | maskExt_186 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h2E)
        v0_187 <= v0_187 & ~maskExt_187 | maskExt_187 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h2F)
        v0_188 <= v0_188 & ~maskExt_188 | maskExt_188 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h2F)
        v0_189 <= v0_189 & ~maskExt_189 | maskExt_189 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h2F)
        v0_190 <= v0_190 & ~maskExt_190 | maskExt_190 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h2F)
        v0_191 <= v0_191 & ~maskExt_191 | maskExt_191 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h30)
        v0_192 <= v0_192 & ~maskExt_192 | maskExt_192 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h30)
        v0_193 <= v0_193 & ~maskExt_193 | maskExt_193 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h30)
        v0_194 <= v0_194 & ~maskExt_194 | maskExt_194 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h30)
        v0_195 <= v0_195 & ~maskExt_195 | maskExt_195 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h31)
        v0_196 <= v0_196 & ~maskExt_196 | maskExt_196 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h31)
        v0_197 <= v0_197 & ~maskExt_197 | maskExt_197 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h31)
        v0_198 <= v0_198 & ~maskExt_198 | maskExt_198 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h31)
        v0_199 <= v0_199 & ~maskExt_199 | maskExt_199 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h32)
        v0_200 <= v0_200 & ~maskExt_200 | maskExt_200 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h32)
        v0_201 <= v0_201 & ~maskExt_201 | maskExt_201 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h32)
        v0_202 <= v0_202 & ~maskExt_202 | maskExt_202 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h32)
        v0_203 <= v0_203 & ~maskExt_203 | maskExt_203 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h33)
        v0_204 <= v0_204 & ~maskExt_204 | maskExt_204 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h33)
        v0_205 <= v0_205 & ~maskExt_205 | maskExt_205 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h33)
        v0_206 <= v0_206 & ~maskExt_206 | maskExt_206 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h33)
        v0_207 <= v0_207 & ~maskExt_207 | maskExt_207 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h34)
        v0_208 <= v0_208 & ~maskExt_208 | maskExt_208 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h34)
        v0_209 <= v0_209 & ~maskExt_209 | maskExt_209 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h34)
        v0_210 <= v0_210 & ~maskExt_210 | maskExt_210 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h34)
        v0_211 <= v0_211 & ~maskExt_211 | maskExt_211 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h35)
        v0_212 <= v0_212 & ~maskExt_212 | maskExt_212 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h35)
        v0_213 <= v0_213 & ~maskExt_213 | maskExt_213 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h35)
        v0_214 <= v0_214 & ~maskExt_214 | maskExt_214 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h35)
        v0_215 <= v0_215 & ~maskExt_215 | maskExt_215 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h36)
        v0_216 <= v0_216 & ~maskExt_216 | maskExt_216 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h36)
        v0_217 <= v0_217 & ~maskExt_217 | maskExt_217 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h36)
        v0_218 <= v0_218 & ~maskExt_218 | maskExt_218 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h36)
        v0_219 <= v0_219 & ~maskExt_219 | maskExt_219 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h37)
        v0_220 <= v0_220 & ~maskExt_220 | maskExt_220 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h37)
        v0_221 <= v0_221 & ~maskExt_221 | maskExt_221 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h37)
        v0_222 <= v0_222 & ~maskExt_222 | maskExt_222 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h37)
        v0_223 <= v0_223 & ~maskExt_223 | maskExt_223 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h38)
        v0_224 <= v0_224 & ~maskExt_224 | maskExt_224 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h38)
        v0_225 <= v0_225 & ~maskExt_225 | maskExt_225 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h38)
        v0_226 <= v0_226 & ~maskExt_226 | maskExt_226 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h38)
        v0_227 <= v0_227 & ~maskExt_227 | maskExt_227 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h39)
        v0_228 <= v0_228 & ~maskExt_228 | maskExt_228 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h39)
        v0_229 <= v0_229 & ~maskExt_229 | maskExt_229 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h39)
        v0_230 <= v0_230 & ~maskExt_230 | maskExt_230 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h39)
        v0_231 <= v0_231 & ~maskExt_231 | maskExt_231 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h3A)
        v0_232 <= v0_232 & ~maskExt_232 | maskExt_232 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h3A)
        v0_233 <= v0_233 & ~maskExt_233 | maskExt_233 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h3A)
        v0_234 <= v0_234 & ~maskExt_234 | maskExt_234 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h3A)
        v0_235 <= v0_235 & ~maskExt_235 | maskExt_235 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h3B)
        v0_236 <= v0_236 & ~maskExt_236 | maskExt_236 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h3B)
        v0_237 <= v0_237 & ~maskExt_237 | maskExt_237 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h3B)
        v0_238 <= v0_238 & ~maskExt_238 | maskExt_238 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h3B)
        v0_239 <= v0_239 & ~maskExt_239 | maskExt_239 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h3C)
        v0_240 <= v0_240 & ~maskExt_240 | maskExt_240 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h3C)
        v0_241 <= v0_241 & ~maskExt_241 | maskExt_241 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h3C)
        v0_242 <= v0_242 & ~maskExt_242 | maskExt_242 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h3C)
        v0_243 <= v0_243 & ~maskExt_243 | maskExt_243 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h3D)
        v0_244 <= v0_244 & ~maskExt_244 | maskExt_244 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h3D)
        v0_245 <= v0_245 & ~maskExt_245 | maskExt_245 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h3D)
        v0_246 <= v0_246 & ~maskExt_246 | maskExt_246 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h3D)
        v0_247 <= v0_247 & ~maskExt_247 | maskExt_247 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 6'h3E)
        v0_248 <= v0_248 & ~maskExt_248 | maskExt_248 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 6'h3E)
        v0_249 <= v0_249 & ~maskExt_249 | maskExt_249 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 6'h3E)
        v0_250 <= v0_250 & ~maskExt_250 | maskExt_250 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 6'h3E)
        v0_251 <= v0_251 & ~maskExt_251 | maskExt_251 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & (&v0UpdateVec_0_bits_offset))
        v0_252 <= v0_252 & ~maskExt_252 | maskExt_252 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & (&v0UpdateVec_1_bits_offset))
        v0_253 <= v0_253 & ~maskExt_253 | maskExt_253 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & (&v0UpdateVec_2_bits_offset))
        v0_254 <= v0_254 & ~maskExt_254 | maskExt_254 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & (&v0UpdateVec_3_bits_offset))
        v0_255 <= v0_255 & ~maskExt_255 | maskExt_255 & v0UpdateVec_3_bits_data;
      if (gatherData_ready_0 & gatherData_valid_0)
        gatherReadState <= 2'h0;
      else if (_tokenCheck_T & gatherSRead)
        gatherReadState <= 2'h2;
      else if (gatherRequestFire)
        gatherReadState <= {notNeedRead, 1'h1};
      else if (readTokenRelease_0 & gatherWaiteRead)
        gatherReadState <= 2'h3;
      if (gatherRequestFire) begin
        gatherDatOffset <= dataOffset;
        gatherLane <= accessLane;
        gatherOffset <= offset;
        gatherGrowth <= reallyGrowth;
      end
      if (_GEN_177 | instReq_valid)
        instReg_instructionIndex <= instReq_bits_instructionIndex;
      if (instReq_valid) begin
        instReg_decodeResult_specialSlot <= instReq_bits_decodeResult_specialSlot;
        instReg_decodeResult_topUop <= instReq_bits_decodeResult_topUop;
        instReg_decodeResult_popCount <= instReq_bits_decodeResult_popCount;
        instReg_decodeResult_ffo <= instReq_bits_decodeResult_ffo;
        instReg_decodeResult_average <= instReq_bits_decodeResult_average;
        instReg_decodeResult_reverse <= instReq_bits_decodeResult_reverse;
        instReg_decodeResult_dontNeedExecuteInLane <= instReq_bits_decodeResult_dontNeedExecuteInLane;
        instReg_decodeResult_scheduler <= instReq_bits_decodeResult_scheduler;
        instReg_decodeResult_sReadVD <= instReq_bits_decodeResult_sReadVD;
        instReg_decodeResult_vtype <= instReq_bits_decodeResult_vtype;
        instReg_decodeResult_sWrite <= instReq_bits_decodeResult_sWrite;
        instReg_decodeResult_crossRead <= instReq_bits_decodeResult_crossRead;
        instReg_decodeResult_crossWrite <= instReq_bits_decodeResult_crossWrite;
        instReg_decodeResult_maskUnit <= instReq_bits_decodeResult_maskUnit;
        instReg_decodeResult_special <= instReq_bits_decodeResult_special;
        instReg_decodeResult_saturate <= instReq_bits_decodeResult_saturate;
        instReg_decodeResult_vwmacc <= instReq_bits_decodeResult_vwmacc;
        instReg_decodeResult_readOnly <= instReq_bits_decodeResult_readOnly;
        instReg_decodeResult_maskSource <= instReq_bits_decodeResult_maskSource;
        instReg_decodeResult_maskDestination <= instReq_bits_decodeResult_maskDestination;
        instReg_decodeResult_maskLogic <= instReq_bits_decodeResult_maskLogic;
        instReg_decodeResult_uop <= instReq_bits_decodeResult_uop;
        instReg_decodeResult_iota <= instReq_bits_decodeResult_iota;
        instReg_decodeResult_mv <= instReq_bits_decodeResult_mv;
        instReg_decodeResult_extend <= instReq_bits_decodeResult_extend;
        instReg_decodeResult_unOrderWrite <= instReq_bits_decodeResult_unOrderWrite;
        instReg_decodeResult_compress <= instReq_bits_decodeResult_compress;
        instReg_decodeResult_gather16 <= instReq_bits_decodeResult_gather16;
        instReg_decodeResult_gather <= instReq_bits_decodeResult_gather;
        instReg_decodeResult_slid <= instReq_bits_decodeResult_slid;
        instReg_decodeResult_targetRd <= instReq_bits_decodeResult_targetRd;
        instReg_decodeResult_widenReduce <= instReq_bits_decodeResult_widenReduce;
        instReg_decodeResult_red <= instReq_bits_decodeResult_red;
        instReg_decodeResult_nr <= instReq_bits_decodeResult_nr;
        instReg_decodeResult_itype <= instReq_bits_decodeResult_itype;
        instReg_decodeResult_unsigned1 <= instReq_bits_decodeResult_unsigned1;
        instReg_decodeResult_unsigned0 <= instReq_bits_decodeResult_unsigned0;
        instReg_decodeResult_other <= instReq_bits_decodeResult_other;
        instReg_decodeResult_multiCycle <= instReq_bits_decodeResult_multiCycle;
        instReg_decodeResult_divider <= instReq_bits_decodeResult_divider;
        instReg_decodeResult_multiplier <= instReq_bits_decodeResult_multiplier;
        instReg_decodeResult_shift <= instReq_bits_decodeResult_shift;
        instReg_decodeResult_adder <= instReq_bits_decodeResult_adder;
        instReg_decodeResult_logic <= instReq_bits_decodeResult_logic;
        instReg_readFromScala <= instReq_bits_readFromScala;
        instReg_sew <= instReq_bits_sew;
        instReg_vlmul <= instReq_bits_vlmul;
        instReg_maskType <= instReq_bits_maskType;
        instReg_vxrm <= instReq_bits_vxrm;
        instReg_vs2 <= instReq_bits_vs2;
        instReg_vd <= instReq_bits_vd;
        instReg_vl <= instReq_bits_vl;
      end
      if (_GEN_177)
        instReg_vs1 <= instReq_bits_vs2;
      else if (instReq_valid)
        instReg_vs1 <= instReq_bits_vs1;
      if (|{instReq_valid, _lastReport_output})
        instVlValid <= ((|instReq_bits_vl) | enqMvRD) & instReq_valid;
      readVS1Reg_dataValid <= ~_GEN_179 & (readTokenRelease_0 | ~_GEN_178 & readVS1Reg_dataValid);
      readVS1Reg_requestSend <= ~_GEN_179 & (_tokenCheck_T | ~_GEN_178 & readVS1Reg_requestSend);
      readVS1Reg_sendToExecution <= _view__firstGroup_T_1 | viotaCounterAdd | ~_GEN_178 & readVS1Reg_sendToExecution;
      if (readTokenRelease_0) begin
        readVS1Reg_data <= readData_readDataQueue_deq_bits;
        waiteReadData_0 <= readData_readDataQueue_deq_bits;
      end
      if (_GEN_179)
        readVS1Reg_readIndex <= readVS1Reg_readIndex + 9'h1;
      else if (_GEN_178)
        readVS1Reg_readIndex <= 9'h0;
      if (tokenIO_0_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_0_valid <= tokenIO_0_maskRequestRelease_0 & ~viota;
      if (tokenIO_0_maskRequestRelease_0) begin
        exeReqReg_0_bits_source1 <= exeRequestQueue_0_deq_bits_source1;
        exeReqReg_0_bits_source2 <= exeRequestQueue_0_deq_bits_source2;
        exeReqReg_0_bits_index <= exeRequestQueue_0_deq_bits_index;
        exeReqReg_0_bits_ffo <= exeRequestQueue_0_deq_bits_ffo;
      end
      if (tokenIO_1_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_1_valid <= tokenIO_1_maskRequestRelease_0 & ~viota;
      if (tokenIO_1_maskRequestRelease_0) begin
        exeReqReg_1_bits_source1 <= exeRequestQueue_1_deq_bits_source1;
        exeReqReg_1_bits_source2 <= exeRequestQueue_1_deq_bits_source2;
        exeReqReg_1_bits_index <= exeRequestQueue_1_deq_bits_index;
        exeReqReg_1_bits_ffo <= exeRequestQueue_1_deq_bits_ffo;
      end
      if (tokenIO_2_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_2_valid <= tokenIO_2_maskRequestRelease_0 & ~viota;
      if (tokenIO_2_maskRequestRelease_0) begin
        exeReqReg_2_bits_source1 <= exeRequestQueue_2_deq_bits_source1;
        exeReqReg_2_bits_source2 <= exeRequestQueue_2_deq_bits_source2;
        exeReqReg_2_bits_index <= exeRequestQueue_2_deq_bits_index;
        exeReqReg_2_bits_ffo <= exeRequestQueue_2_deq_bits_ffo;
      end
      if (tokenIO_3_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_3_valid <= tokenIO_3_maskRequestRelease_0 & ~viota;
      if (tokenIO_3_maskRequestRelease_0) begin
        exeReqReg_3_bits_source1 <= exeRequestQueue_3_deq_bits_source1;
        exeReqReg_3_bits_source2 <= exeRequestQueue_3_deq_bits_source2;
        exeReqReg_3_bits_index <= exeRequestQueue_3_deq_bits_index;
        exeReqReg_3_bits_ffo <= exeRequestQueue_3_deq_bits_ffo;
      end
      if (instReq_valid | groupCounterAdd)
        requestCounter <= instReq_valid ? 10'h0 : requestCounter + 10'h1;
      if (requestStageDeq & anyDataValid)
        executeIndex <= executeIndex + executeIndexGrowth[1:0];
      if (readIssueStageEnq) begin
        readIssueStageState_groupReadState <= 4'h0;
        readIssueStageState_needRead <= _GEN_170 ? _slideAddressGen_indexDeq_bits_needRead : ~notReadSelect;
        readIssueStageState_elementValid <= _GEN_170 ? _slideAddressGen_indexDeq_bits_elementValid : elementValidSelect;
        readIssueStageState_replaceVs1 <= _GEN_170 ? _slideAddressGen_indexDeq_bits_replaceVs1 : 4'h0;
        readIssueStageState_readOffset <= _GEN_170 ? _slideAddressGen_indexDeq_bits_readOffset : offsetSelect;
        readIssueStageState_accessLane_0 <= _GEN_170 ? _slideAddressGen_indexDeq_bits_accessLane_0 : accessLaneSelect[1:0];
        readIssueStageState_accessLane_1 <= _GEN_170 ? _slideAddressGen_indexDeq_bits_accessLane_1 : accessLaneSelect[3:2];
        readIssueStageState_accessLane_2 <= _GEN_170 ? _slideAddressGen_indexDeq_bits_accessLane_2 : accessLaneSelect[5:4];
        readIssueStageState_accessLane_3 <= _GEN_170 ? _slideAddressGen_indexDeq_bits_accessLane_3 : accessLaneSelect[7:6];
        readIssueStageState_vsGrowth_0 <= _GEN_170 ? _slideAddressGen_indexDeq_bits_vsGrowth_0 : growthSelect[2:0];
        readIssueStageState_vsGrowth_1 <= _GEN_170 ? _slideAddressGen_indexDeq_bits_vsGrowth_1 : growthSelect[5:3];
        readIssueStageState_vsGrowth_2 <= _GEN_170 ? _slideAddressGen_indexDeq_bits_vsGrowth_2 : growthSelect[8:6];
        readIssueStageState_vsGrowth_3 <= _GEN_170 ? _slideAddressGen_indexDeq_bits_vsGrowth_3 : growthSelect[11:9];
        readIssueStageState_executeGroup <= _GEN_170 ? _slideAddressGen_indexDeq_bits_executeGroup : executeGroup;
        readIssueStageState_readDataOffset <= _GEN_170 ? _slideAddressGen_indexDeq_bits_readDataOffset : dataOffsetSelect;
        readIssueStageState_last <= _GEN_170 ? _slideAddressGen_indexDeq_bits_last : isVlBoundary;
      end
      else if (anyReadFire)
        readIssueStageState_groupReadState <= readStateUpdate;
      if (readTypeRequestDeq ^ readIssueStageEnq)
        readIssueStageValid <= readIssueStageEnq;
      if (_tokenCheck_T ^ readTokenRelease_0)
        tokenCheck_counter <= tokenCheck_counter + tokenCheck_counterChange;
      if (pipeReadFire_1 ^ readTokenRelease_1)
        tokenCheck_counter_1 <= tokenCheck_counter_1 + tokenCheck_counterChange_1;
      if (pipeReadFire_2 ^ readTokenRelease_2)
        tokenCheck_counter_2 <= tokenCheck_counter_2 + tokenCheck_counterChange_2;
      if (pipeReadFire_3 ^ readTokenRelease_3)
        tokenCheck_counter_3 <= tokenCheck_counter_3 + tokenCheck_counterChange_3;
      if (reorderQueueAllocate_release | readIssueStageEnq) begin
        reorderQueueAllocate_counter <= reorderQueueAllocate_counterUpdate;
        reorderQueueAllocate_counterWillUpdate <= reorderQueueAllocate_counterUpdate + 4'h4;
      end
      if (reorderQueueAllocate_release_1 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_1 <= reorderQueueAllocate_counterUpdate_1;
        reorderQueueAllocate_counterWillUpdate_1 <= reorderQueueAllocate_counterUpdate_1 + 4'h4;
      end
      if (reorderQueueAllocate_release_2 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_2 <= reorderQueueAllocate_counterUpdate_2;
        reorderQueueAllocate_counterWillUpdate_2 <= reorderQueueAllocate_counterUpdate_2 + 4'h4;
      end
      if (reorderQueueAllocate_release_3 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_3 <= reorderQueueAllocate_counterUpdate_3;
        reorderQueueAllocate_counterWillUpdate_3 <= reorderQueueAllocate_counterUpdate_3 + 4'h4;
      end
      if (reorderStageEnqFire ^ reorderStageDeqFire)
        reorderStageValid <= reorderStageEnqFire;
      if (_write1HPipe_0_T & readType)
        reorderStageState_0 <= reorderStageState_0 + 3'h1;
      else if (reorderStageEnqFire)
        reorderStageState_0 <= 3'h0;
      if (_write1HPipe_1_T & readType)
        reorderStageState_1 <= reorderStageState_1 + 3'h1;
      else if (reorderStageEnqFire)
        reorderStageState_1 <= 3'h0;
      if (_write1HPipe_2_T & readType)
        reorderStageState_2 <= reorderStageState_2 + 3'h1;
      else if (reorderStageEnqFire)
        reorderStageState_2 <= 3'h0;
      if (_write1HPipe_3_T & readType)
        reorderStageState_3 <= reorderStageState_3 + 3'h1;
      else if (reorderStageEnqFire)
        reorderStageState_3 <= 3'h0;
      if (reorderStageEnqFire) begin
        reorderStageNeed_0 <= accessCountQueue_deq_bits_0;
        reorderStageNeed_1 <= accessCountQueue_deq_bits_1;
        reorderStageNeed_2 <= accessCountQueue_deq_bits_2;
        reorderStageNeed_3 <= accessCountQueue_deq_bits_3;
      end
      if (waiteStageEnqFire) begin
        waiteReadDataPipeReg_executeGroup <= readWaitQueue_deq_bits_executeGroup;
        waiteReadDataPipeReg_sourceValid <= readWaitQueue_deq_bits_sourceValid;
        waiteReadDataPipeReg_replaceVs1 <= readWaitQueue_deq_bits_replaceVs1;
        waiteReadDataPipeReg_needRead <= readWaitQueue_deq_bits_needRead;
        waiteReadDataPipeReg_last <= readWaitQueue_deq_bits_last;
      end
      if (readTokenRelease_1)
        waiteReadData_1 <= readData_readDataQueue_1_deq_bits;
      if (readTokenRelease_2)
        waiteReadData_2 <= readData_readDataQueue_2_deq_bits;
      if (readTokenRelease_3)
        waiteReadData_3 <= readData_readDataQueue_3_deq_bits;
      if (waiteStageEnqFire & (|readResultValid))
        waiteReadSate <= readResultValid;
      else if (|readResultValid)
        waiteReadSate <= waiteReadSate | readResultValid;
      else if (waiteStageEnqFire)
        waiteReadSate <= 4'h0;
      if (waiteStageDeqFire ^ waiteStageEnqFire)
        waiteReadStageValid <= waiteStageEnqFire;
      if (_dataNotInShifter_T ^ writeRelease_0)
        dataNotInShifter_writeTokenCounter <= dataNotInShifter_writeTokenCounter + dataNotInShifter_writeTokenChange;
      if (_dataNotInShifter_T_3 ^ writeRelease_1)
        dataNotInShifter_writeTokenCounter_1 <= dataNotInShifter_writeTokenCounter_1 + dataNotInShifter_writeTokenChange_1;
      if (_dataNotInShifter_T_6 ^ writeRelease_2)
        dataNotInShifter_writeTokenCounter_2 <= dataNotInShifter_writeTokenCounter_2 + dataNotInShifter_writeTokenChange_2;
      if (_dataNotInShifter_T_9 ^ writeRelease_3)
        dataNotInShifter_writeTokenCounter_3 <= dataNotInShifter_writeTokenCounter_3 + dataNotInShifter_writeTokenChange_3;
      waiteLastRequest <= ~readType & requestStageDeq & lastGroup | ~lastReportValid & waiteLastRequest;
      waitQueueClear <= executeStageClean | invalidEnq | ~lastReportValid & waitQueueClear;
    end
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:281];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [8:0] i = 9'h0; i < 9'h11A; i += 9'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        v0_0 = _RANDOM[9'h0];
        v0_1 = _RANDOM[9'h1];
        v0_2 = _RANDOM[9'h2];
        v0_3 = _RANDOM[9'h3];
        v0_4 = _RANDOM[9'h4];
        v0_5 = _RANDOM[9'h5];
        v0_6 = _RANDOM[9'h6];
        v0_7 = _RANDOM[9'h7];
        v0_8 = _RANDOM[9'h8];
        v0_9 = _RANDOM[9'h9];
        v0_10 = _RANDOM[9'hA];
        v0_11 = _RANDOM[9'hB];
        v0_12 = _RANDOM[9'hC];
        v0_13 = _RANDOM[9'hD];
        v0_14 = _RANDOM[9'hE];
        v0_15 = _RANDOM[9'hF];
        v0_16 = _RANDOM[9'h10];
        v0_17 = _RANDOM[9'h11];
        v0_18 = _RANDOM[9'h12];
        v0_19 = _RANDOM[9'h13];
        v0_20 = _RANDOM[9'h14];
        v0_21 = _RANDOM[9'h15];
        v0_22 = _RANDOM[9'h16];
        v0_23 = _RANDOM[9'h17];
        v0_24 = _RANDOM[9'h18];
        v0_25 = _RANDOM[9'h19];
        v0_26 = _RANDOM[9'h1A];
        v0_27 = _RANDOM[9'h1B];
        v0_28 = _RANDOM[9'h1C];
        v0_29 = _RANDOM[9'h1D];
        v0_30 = _RANDOM[9'h1E];
        v0_31 = _RANDOM[9'h1F];
        v0_32 = _RANDOM[9'h20];
        v0_33 = _RANDOM[9'h21];
        v0_34 = _RANDOM[9'h22];
        v0_35 = _RANDOM[9'h23];
        v0_36 = _RANDOM[9'h24];
        v0_37 = _RANDOM[9'h25];
        v0_38 = _RANDOM[9'h26];
        v0_39 = _RANDOM[9'h27];
        v0_40 = _RANDOM[9'h28];
        v0_41 = _RANDOM[9'h29];
        v0_42 = _RANDOM[9'h2A];
        v0_43 = _RANDOM[9'h2B];
        v0_44 = _RANDOM[9'h2C];
        v0_45 = _RANDOM[9'h2D];
        v0_46 = _RANDOM[9'h2E];
        v0_47 = _RANDOM[9'h2F];
        v0_48 = _RANDOM[9'h30];
        v0_49 = _RANDOM[9'h31];
        v0_50 = _RANDOM[9'h32];
        v0_51 = _RANDOM[9'h33];
        v0_52 = _RANDOM[9'h34];
        v0_53 = _RANDOM[9'h35];
        v0_54 = _RANDOM[9'h36];
        v0_55 = _RANDOM[9'h37];
        v0_56 = _RANDOM[9'h38];
        v0_57 = _RANDOM[9'h39];
        v0_58 = _RANDOM[9'h3A];
        v0_59 = _RANDOM[9'h3B];
        v0_60 = _RANDOM[9'h3C];
        v0_61 = _RANDOM[9'h3D];
        v0_62 = _RANDOM[9'h3E];
        v0_63 = _RANDOM[9'h3F];
        v0_64 = _RANDOM[9'h40];
        v0_65 = _RANDOM[9'h41];
        v0_66 = _RANDOM[9'h42];
        v0_67 = _RANDOM[9'h43];
        v0_68 = _RANDOM[9'h44];
        v0_69 = _RANDOM[9'h45];
        v0_70 = _RANDOM[9'h46];
        v0_71 = _RANDOM[9'h47];
        v0_72 = _RANDOM[9'h48];
        v0_73 = _RANDOM[9'h49];
        v0_74 = _RANDOM[9'h4A];
        v0_75 = _RANDOM[9'h4B];
        v0_76 = _RANDOM[9'h4C];
        v0_77 = _RANDOM[9'h4D];
        v0_78 = _RANDOM[9'h4E];
        v0_79 = _RANDOM[9'h4F];
        v0_80 = _RANDOM[9'h50];
        v0_81 = _RANDOM[9'h51];
        v0_82 = _RANDOM[9'h52];
        v0_83 = _RANDOM[9'h53];
        v0_84 = _RANDOM[9'h54];
        v0_85 = _RANDOM[9'h55];
        v0_86 = _RANDOM[9'h56];
        v0_87 = _RANDOM[9'h57];
        v0_88 = _RANDOM[9'h58];
        v0_89 = _RANDOM[9'h59];
        v0_90 = _RANDOM[9'h5A];
        v0_91 = _RANDOM[9'h5B];
        v0_92 = _RANDOM[9'h5C];
        v0_93 = _RANDOM[9'h5D];
        v0_94 = _RANDOM[9'h5E];
        v0_95 = _RANDOM[9'h5F];
        v0_96 = _RANDOM[9'h60];
        v0_97 = _RANDOM[9'h61];
        v0_98 = _RANDOM[9'h62];
        v0_99 = _RANDOM[9'h63];
        v0_100 = _RANDOM[9'h64];
        v0_101 = _RANDOM[9'h65];
        v0_102 = _RANDOM[9'h66];
        v0_103 = _RANDOM[9'h67];
        v0_104 = _RANDOM[9'h68];
        v0_105 = _RANDOM[9'h69];
        v0_106 = _RANDOM[9'h6A];
        v0_107 = _RANDOM[9'h6B];
        v0_108 = _RANDOM[9'h6C];
        v0_109 = _RANDOM[9'h6D];
        v0_110 = _RANDOM[9'h6E];
        v0_111 = _RANDOM[9'h6F];
        v0_112 = _RANDOM[9'h70];
        v0_113 = _RANDOM[9'h71];
        v0_114 = _RANDOM[9'h72];
        v0_115 = _RANDOM[9'h73];
        v0_116 = _RANDOM[9'h74];
        v0_117 = _RANDOM[9'h75];
        v0_118 = _RANDOM[9'h76];
        v0_119 = _RANDOM[9'h77];
        v0_120 = _RANDOM[9'h78];
        v0_121 = _RANDOM[9'h79];
        v0_122 = _RANDOM[9'h7A];
        v0_123 = _RANDOM[9'h7B];
        v0_124 = _RANDOM[9'h7C];
        v0_125 = _RANDOM[9'h7D];
        v0_126 = _RANDOM[9'h7E];
        v0_127 = _RANDOM[9'h7F];
        v0_128 = _RANDOM[9'h80];
        v0_129 = _RANDOM[9'h81];
        v0_130 = _RANDOM[9'h82];
        v0_131 = _RANDOM[9'h83];
        v0_132 = _RANDOM[9'h84];
        v0_133 = _RANDOM[9'h85];
        v0_134 = _RANDOM[9'h86];
        v0_135 = _RANDOM[9'h87];
        v0_136 = _RANDOM[9'h88];
        v0_137 = _RANDOM[9'h89];
        v0_138 = _RANDOM[9'h8A];
        v0_139 = _RANDOM[9'h8B];
        v0_140 = _RANDOM[9'h8C];
        v0_141 = _RANDOM[9'h8D];
        v0_142 = _RANDOM[9'h8E];
        v0_143 = _RANDOM[9'h8F];
        v0_144 = _RANDOM[9'h90];
        v0_145 = _RANDOM[9'h91];
        v0_146 = _RANDOM[9'h92];
        v0_147 = _RANDOM[9'h93];
        v0_148 = _RANDOM[9'h94];
        v0_149 = _RANDOM[9'h95];
        v0_150 = _RANDOM[9'h96];
        v0_151 = _RANDOM[9'h97];
        v0_152 = _RANDOM[9'h98];
        v0_153 = _RANDOM[9'h99];
        v0_154 = _RANDOM[9'h9A];
        v0_155 = _RANDOM[9'h9B];
        v0_156 = _RANDOM[9'h9C];
        v0_157 = _RANDOM[9'h9D];
        v0_158 = _RANDOM[9'h9E];
        v0_159 = _RANDOM[9'h9F];
        v0_160 = _RANDOM[9'hA0];
        v0_161 = _RANDOM[9'hA1];
        v0_162 = _RANDOM[9'hA2];
        v0_163 = _RANDOM[9'hA3];
        v0_164 = _RANDOM[9'hA4];
        v0_165 = _RANDOM[9'hA5];
        v0_166 = _RANDOM[9'hA6];
        v0_167 = _RANDOM[9'hA7];
        v0_168 = _RANDOM[9'hA8];
        v0_169 = _RANDOM[9'hA9];
        v0_170 = _RANDOM[9'hAA];
        v0_171 = _RANDOM[9'hAB];
        v0_172 = _RANDOM[9'hAC];
        v0_173 = _RANDOM[9'hAD];
        v0_174 = _RANDOM[9'hAE];
        v0_175 = _RANDOM[9'hAF];
        v0_176 = _RANDOM[9'hB0];
        v0_177 = _RANDOM[9'hB1];
        v0_178 = _RANDOM[9'hB2];
        v0_179 = _RANDOM[9'hB3];
        v0_180 = _RANDOM[9'hB4];
        v0_181 = _RANDOM[9'hB5];
        v0_182 = _RANDOM[9'hB6];
        v0_183 = _RANDOM[9'hB7];
        v0_184 = _RANDOM[9'hB8];
        v0_185 = _RANDOM[9'hB9];
        v0_186 = _RANDOM[9'hBA];
        v0_187 = _RANDOM[9'hBB];
        v0_188 = _RANDOM[9'hBC];
        v0_189 = _RANDOM[9'hBD];
        v0_190 = _RANDOM[9'hBE];
        v0_191 = _RANDOM[9'hBF];
        v0_192 = _RANDOM[9'hC0];
        v0_193 = _RANDOM[9'hC1];
        v0_194 = _RANDOM[9'hC2];
        v0_195 = _RANDOM[9'hC3];
        v0_196 = _RANDOM[9'hC4];
        v0_197 = _RANDOM[9'hC5];
        v0_198 = _RANDOM[9'hC6];
        v0_199 = _RANDOM[9'hC7];
        v0_200 = _RANDOM[9'hC8];
        v0_201 = _RANDOM[9'hC9];
        v0_202 = _RANDOM[9'hCA];
        v0_203 = _RANDOM[9'hCB];
        v0_204 = _RANDOM[9'hCC];
        v0_205 = _RANDOM[9'hCD];
        v0_206 = _RANDOM[9'hCE];
        v0_207 = _RANDOM[9'hCF];
        v0_208 = _RANDOM[9'hD0];
        v0_209 = _RANDOM[9'hD1];
        v0_210 = _RANDOM[9'hD2];
        v0_211 = _RANDOM[9'hD3];
        v0_212 = _RANDOM[9'hD4];
        v0_213 = _RANDOM[9'hD5];
        v0_214 = _RANDOM[9'hD6];
        v0_215 = _RANDOM[9'hD7];
        v0_216 = _RANDOM[9'hD8];
        v0_217 = _RANDOM[9'hD9];
        v0_218 = _RANDOM[9'hDA];
        v0_219 = _RANDOM[9'hDB];
        v0_220 = _RANDOM[9'hDC];
        v0_221 = _RANDOM[9'hDD];
        v0_222 = _RANDOM[9'hDE];
        v0_223 = _RANDOM[9'hDF];
        v0_224 = _RANDOM[9'hE0];
        v0_225 = _RANDOM[9'hE1];
        v0_226 = _RANDOM[9'hE2];
        v0_227 = _RANDOM[9'hE3];
        v0_228 = _RANDOM[9'hE4];
        v0_229 = _RANDOM[9'hE5];
        v0_230 = _RANDOM[9'hE6];
        v0_231 = _RANDOM[9'hE7];
        v0_232 = _RANDOM[9'hE8];
        v0_233 = _RANDOM[9'hE9];
        v0_234 = _RANDOM[9'hEA];
        v0_235 = _RANDOM[9'hEB];
        v0_236 = _RANDOM[9'hEC];
        v0_237 = _RANDOM[9'hED];
        v0_238 = _RANDOM[9'hEE];
        v0_239 = _RANDOM[9'hEF];
        v0_240 = _RANDOM[9'hF0];
        v0_241 = _RANDOM[9'hF1];
        v0_242 = _RANDOM[9'hF2];
        v0_243 = _RANDOM[9'hF3];
        v0_244 = _RANDOM[9'hF4];
        v0_245 = _RANDOM[9'hF5];
        v0_246 = _RANDOM[9'hF6];
        v0_247 = _RANDOM[9'hF7];
        v0_248 = _RANDOM[9'hF8];
        v0_249 = _RANDOM[9'hF9];
        v0_250 = _RANDOM[9'hFA];
        v0_251 = _RANDOM[9'hFB];
        v0_252 = _RANDOM[9'hFC];
        v0_253 = _RANDOM[9'hFD];
        v0_254 = _RANDOM[9'hFE];
        v0_255 = _RANDOM[9'hFF];
        gatherReadState = _RANDOM[9'h100][1:0];
        gatherDatOffset = _RANDOM[9'h100][3:2];
        gatherLane = _RANDOM[9'h100][5:4];
        gatherOffset = _RANDOM[9'h100][11:6];
        gatherGrowth = _RANDOM[9'h100][14:12];
        instReg_instructionIndex = _RANDOM[9'h100][17:15];
        instReg_decodeResult_specialSlot = _RANDOM[9'h100][18];
        instReg_decodeResult_topUop = _RANDOM[9'h100][23:19];
        instReg_decodeResult_popCount = _RANDOM[9'h100][24];
        instReg_decodeResult_ffo = _RANDOM[9'h100][25];
        instReg_decodeResult_average = _RANDOM[9'h100][26];
        instReg_decodeResult_reverse = _RANDOM[9'h100][27];
        instReg_decodeResult_dontNeedExecuteInLane = _RANDOM[9'h100][28];
        instReg_decodeResult_scheduler = _RANDOM[9'h100][29];
        instReg_decodeResult_sReadVD = _RANDOM[9'h100][30];
        instReg_decodeResult_vtype = _RANDOM[9'h100][31];
        instReg_decodeResult_sWrite = _RANDOM[9'h101][0];
        instReg_decodeResult_crossRead = _RANDOM[9'h101][1];
        instReg_decodeResult_crossWrite = _RANDOM[9'h101][2];
        instReg_decodeResult_maskUnit = _RANDOM[9'h101][3];
        instReg_decodeResult_special = _RANDOM[9'h101][4];
        instReg_decodeResult_saturate = _RANDOM[9'h101][5];
        instReg_decodeResult_vwmacc = _RANDOM[9'h101][6];
        instReg_decodeResult_readOnly = _RANDOM[9'h101][7];
        instReg_decodeResult_maskSource = _RANDOM[9'h101][8];
        instReg_decodeResult_maskDestination = _RANDOM[9'h101][9];
        instReg_decodeResult_maskLogic = _RANDOM[9'h101][10];
        instReg_decodeResult_uop = _RANDOM[9'h101][14:11];
        instReg_decodeResult_iota = _RANDOM[9'h101][15];
        instReg_decodeResult_mv = _RANDOM[9'h101][16];
        instReg_decodeResult_extend = _RANDOM[9'h101][17];
        instReg_decodeResult_unOrderWrite = _RANDOM[9'h101][18];
        instReg_decodeResult_compress = _RANDOM[9'h101][19];
        instReg_decodeResult_gather16 = _RANDOM[9'h101][20];
        instReg_decodeResult_gather = _RANDOM[9'h101][21];
        instReg_decodeResult_slid = _RANDOM[9'h101][22];
        instReg_decodeResult_targetRd = _RANDOM[9'h101][23];
        instReg_decodeResult_widenReduce = _RANDOM[9'h101][24];
        instReg_decodeResult_red = _RANDOM[9'h101][25];
        instReg_decodeResult_nr = _RANDOM[9'h101][26];
        instReg_decodeResult_itype = _RANDOM[9'h101][27];
        instReg_decodeResult_unsigned1 = _RANDOM[9'h101][28];
        instReg_decodeResult_unsigned0 = _RANDOM[9'h101][29];
        instReg_decodeResult_other = _RANDOM[9'h101][30];
        instReg_decodeResult_multiCycle = _RANDOM[9'h101][31];
        instReg_decodeResult_divider = _RANDOM[9'h102][0];
        instReg_decodeResult_multiplier = _RANDOM[9'h102][1];
        instReg_decodeResult_shift = _RANDOM[9'h102][2];
        instReg_decodeResult_adder = _RANDOM[9'h102][3];
        instReg_decodeResult_logic = _RANDOM[9'h102][4];
        instReg_readFromScala = {_RANDOM[9'h102][31:5], _RANDOM[9'h103][4:0]};
        instReg_sew = _RANDOM[9'h103][6:5];
        instReg_vlmul = _RANDOM[9'h103][9:7];
        instReg_maskType = _RANDOM[9'h103][10];
        instReg_vxrm = _RANDOM[9'h103][13:11];
        instReg_vs2 = _RANDOM[9'h103][18:14];
        instReg_vs1 = _RANDOM[9'h103][23:19];
        instReg_vd = _RANDOM[9'h103][28:24];
        instReg_vl = {_RANDOM[9'h103][31:29], _RANDOM[9'h104][10:0]};
        instVlValid = _RANDOM[9'h104][11];
        readVS1Reg_dataValid = _RANDOM[9'h104][12];
        readVS1Reg_requestSend = _RANDOM[9'h104][13];
        readVS1Reg_sendToExecution = _RANDOM[9'h104][14];
        readVS1Reg_data = {_RANDOM[9'h104][31:15], _RANDOM[9'h105][14:0]};
        readVS1Reg_readIndex = _RANDOM[9'h105][23:15];
        exeReqReg_0_valid = _RANDOM[9'h105][28];
        exeReqReg_0_bits_source1 = {_RANDOM[9'h105][31:29], _RANDOM[9'h106][28:0]};
        exeReqReg_0_bits_source2 = {_RANDOM[9'h106][31:29], _RANDOM[9'h107][28:0]};
        exeReqReg_0_bits_index = _RANDOM[9'h107][31:29];
        exeReqReg_0_bits_ffo = _RANDOM[9'h108][0];
        exeReqReg_1_valid = _RANDOM[9'h108][1];
        exeReqReg_1_bits_source1 = {_RANDOM[9'h108][31:2], _RANDOM[9'h109][1:0]};
        exeReqReg_1_bits_source2 = {_RANDOM[9'h109][31:2], _RANDOM[9'h10A][1:0]};
        exeReqReg_1_bits_index = _RANDOM[9'h10A][4:2];
        exeReqReg_1_bits_ffo = _RANDOM[9'h10A][5];
        exeReqReg_2_valid = _RANDOM[9'h10A][6];
        exeReqReg_2_bits_source1 = {_RANDOM[9'h10A][31:7], _RANDOM[9'h10B][6:0]};
        exeReqReg_2_bits_source2 = {_RANDOM[9'h10B][31:7], _RANDOM[9'h10C][6:0]};
        exeReqReg_2_bits_index = _RANDOM[9'h10C][9:7];
        exeReqReg_2_bits_ffo = _RANDOM[9'h10C][10];
        exeReqReg_3_valid = _RANDOM[9'h10C][11];
        exeReqReg_3_bits_source1 = {_RANDOM[9'h10C][31:12], _RANDOM[9'h10D][11:0]};
        exeReqReg_3_bits_source2 = {_RANDOM[9'h10D][31:12], _RANDOM[9'h10E][11:0]};
        exeReqReg_3_bits_index = _RANDOM[9'h10E][14:12];
        exeReqReg_3_bits_ffo = _RANDOM[9'h10E][15];
        requestCounter = _RANDOM[9'h10E][25:16];
        executeIndex = _RANDOM[9'h10E][27:26];
        readIssueStageState_groupReadState = _RANDOM[9'h10E][31:28];
        readIssueStageState_needRead = _RANDOM[9'h10F][3:0];
        readIssueStageState_elementValid = _RANDOM[9'h10F][7:4];
        readIssueStageState_replaceVs1 = _RANDOM[9'h10F][11:8];
        readIssueStageState_readOffset = {_RANDOM[9'h10F][31:12], _RANDOM[9'h110][3:0]};
        readIssueStageState_accessLane_0 = _RANDOM[9'h110][5:4];
        readIssueStageState_accessLane_1 = _RANDOM[9'h110][7:6];
        readIssueStageState_accessLane_2 = _RANDOM[9'h110][9:8];
        readIssueStageState_accessLane_3 = _RANDOM[9'h110][11:10];
        readIssueStageState_vsGrowth_0 = _RANDOM[9'h110][14:12];
        readIssueStageState_vsGrowth_1 = _RANDOM[9'h110][17:15];
        readIssueStageState_vsGrowth_2 = _RANDOM[9'h110][20:18];
        readIssueStageState_vsGrowth_3 = _RANDOM[9'h110][23:21];
        readIssueStageState_executeGroup = {_RANDOM[9'h110][31:24], _RANDOM[9'h111][3:0]};
        readIssueStageState_readDataOffset = _RANDOM[9'h111][11:4];
        readIssueStageState_last = _RANDOM[9'h111][12];
        readIssueStageValid = _RANDOM[9'h111][13];
        tokenCheck_counter = _RANDOM[9'h111][17:14];
        tokenCheck_counter_1 = _RANDOM[9'h111][21:18];
        tokenCheck_counter_2 = _RANDOM[9'h111][25:22];
        tokenCheck_counter_3 = _RANDOM[9'h111][29:26];
        reorderQueueAllocate_counter = {_RANDOM[9'h111][31:30], _RANDOM[9'h112][1:0]};
        reorderQueueAllocate_counterWillUpdate = _RANDOM[9'h112][5:2];
        reorderQueueAllocate_counter_1 = _RANDOM[9'h112][9:6];
        reorderQueueAllocate_counterWillUpdate_1 = _RANDOM[9'h112][13:10];
        reorderQueueAllocate_counter_2 = _RANDOM[9'h112][17:14];
        reorderQueueAllocate_counterWillUpdate_2 = _RANDOM[9'h112][21:18];
        reorderQueueAllocate_counter_3 = _RANDOM[9'h112][25:22];
        reorderQueueAllocate_counterWillUpdate_3 = _RANDOM[9'h112][29:26];
        reorderStageValid = _RANDOM[9'h112][30];
        reorderStageState_0 = {_RANDOM[9'h112][31], _RANDOM[9'h113][1:0]};
        reorderStageState_1 = _RANDOM[9'h113][4:2];
        reorderStageState_2 = _RANDOM[9'h113][7:5];
        reorderStageState_3 = _RANDOM[9'h113][10:8];
        reorderStageNeed_0 = _RANDOM[9'h113][13:11];
        reorderStageNeed_1 = _RANDOM[9'h113][16:14];
        reorderStageNeed_2 = _RANDOM[9'h113][19:17];
        reorderStageNeed_3 = _RANDOM[9'h113][22:20];
        waiteReadDataPipeReg_executeGroup = {_RANDOM[9'h113][31:23], _RANDOM[9'h114][2:0]};
        waiteReadDataPipeReg_sourceValid = _RANDOM[9'h114][6:3];
        waiteReadDataPipeReg_replaceVs1 = _RANDOM[9'h114][10:7];
        waiteReadDataPipeReg_needRead = _RANDOM[9'h114][14:11];
        waiteReadDataPipeReg_last = _RANDOM[9'h114][15];
        waiteReadData_0 = {_RANDOM[9'h114][31:16], _RANDOM[9'h115][15:0]};
        waiteReadData_1 = {_RANDOM[9'h115][31:16], _RANDOM[9'h116][15:0]};
        waiteReadData_2 = {_RANDOM[9'h116][31:16], _RANDOM[9'h117][15:0]};
        waiteReadData_3 = {_RANDOM[9'h117][31:16], _RANDOM[9'h118][15:0]};
        waiteReadSate = _RANDOM[9'h118][19:16];
        waiteReadStageValid = _RANDOM[9'h118][20];
        dataNotInShifter_writeTokenCounter = _RANDOM[9'h118][23:21];
        dataNotInShifter_writeTokenCounter_1 = _RANDOM[9'h118][26:24];
        dataNotInShifter_writeTokenCounter_2 = _RANDOM[9'h118][29:27];
        dataNotInShifter_writeTokenCounter_3 = {_RANDOM[9'h118][31:30], _RANDOM[9'h119][0]};
        waiteLastRequest = _RANDOM[9'h119][1];
        waitQueueClear = _RANDOM[9'h119][2];
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  wire               exeRequestQueue_0_empty;
  assign exeRequestQueue_0_empty = _exeRequestQueue_queue_fifo_empty;
  wire               exeRequestQueue_0_full;
  assign exeRequestQueue_0_full = _exeRequestQueue_queue_fifo_full;
  wire               exeRequestQueue_1_empty;
  assign exeRequestQueue_1_empty = _exeRequestQueue_queue_fifo_1_empty;
  wire               exeRequestQueue_1_full;
  assign exeRequestQueue_1_full = _exeRequestQueue_queue_fifo_1_full;
  wire               exeRequestQueue_2_empty;
  assign exeRequestQueue_2_empty = _exeRequestQueue_queue_fifo_2_empty;
  wire               exeRequestQueue_2_full;
  assign exeRequestQueue_2_full = _exeRequestQueue_queue_fifo_2_full;
  wire               exeRequestQueue_3_empty;
  assign exeRequestQueue_3_empty = _exeRequestQueue_queue_fifo_3_empty;
  wire               exeRequestQueue_3_full;
  assign exeRequestQueue_3_full = _exeRequestQueue_queue_fifo_3_full;
  wire               accessCountQueue_empty;
  assign accessCountQueue_empty = _accessCountQueue_fifo_empty;
  wire               accessCountQueue_full;
  assign accessCountQueue_full = _accessCountQueue_fifo_full;
  wire               readWaitQueue_empty;
  assign readWaitQueue_empty = _readWaitQueue_fifo_empty;
  wire               readWaitQueue_full;
  assign readWaitQueue_full = _readWaitQueue_fifo_full;
  assign compressUnitResultQueue_empty = _compressUnitResultQueue_fifo_empty;
  wire               compressUnitResultQueue_full;
  assign compressUnitResultQueue_full = _compressUnitResultQueue_fifo_full;
  wire               reorderQueueVec_0_empty;
  assign reorderQueueVec_0_empty = _reorderQueueVec_fifo_empty;
  wire               reorderQueueVec_0_full;
  assign reorderQueueVec_0_full = _reorderQueueVec_fifo_full;
  wire               reorderQueueVec_1_empty;
  assign reorderQueueVec_1_empty = _reorderQueueVec_fifo_1_empty;
  wire               reorderQueueVec_1_full;
  assign reorderQueueVec_1_full = _reorderQueueVec_fifo_1_full;
  wire               reorderQueueVec_2_empty;
  assign reorderQueueVec_2_empty = _reorderQueueVec_fifo_2_empty;
  wire               reorderQueueVec_2_full;
  assign reorderQueueVec_2_full = _reorderQueueVec_fifo_2_full;
  wire               reorderQueueVec_3_empty;
  assign reorderQueueVec_3_empty = _reorderQueueVec_fifo_3_empty;
  wire               reorderQueueVec_3_full;
  assign reorderQueueVec_3_full = _reorderQueueVec_fifo_3_full;
  wire               readMessageQueue_empty;
  assign readMessageQueue_empty = _readMessageQueue_fifo_empty;
  wire               readMessageQueue_full;
  assign readMessageQueue_full = _readMessageQueue_fifo_full;
  wire               readMessageQueue_1_empty;
  assign readMessageQueue_1_empty = _readMessageQueue_fifo_1_empty;
  wire               readMessageQueue_1_full;
  assign readMessageQueue_1_full = _readMessageQueue_fifo_1_full;
  wire               readMessageQueue_2_empty;
  assign readMessageQueue_2_empty = _readMessageQueue_fifo_2_empty;
  wire               readMessageQueue_2_full;
  assign readMessageQueue_2_full = _readMessageQueue_fifo_2_full;
  wire               readMessageQueue_3_empty;
  assign readMessageQueue_3_empty = _readMessageQueue_fifo_3_empty;
  wire               readMessageQueue_3_full;
  assign readMessageQueue_3_full = _readMessageQueue_fifo_3_full;
  wire               readData_readDataQueue_empty;
  assign readData_readDataQueue_empty = _readData_readDataQueue_fifo_empty;
  wire               readData_readDataQueue_full;
  assign readData_readDataQueue_full = _readData_readDataQueue_fifo_full;
  wire               readData_readDataQueue_1_empty;
  assign readData_readDataQueue_1_empty = _readData_readDataQueue_fifo_1_empty;
  wire               readData_readDataQueue_1_full;
  assign readData_readDataQueue_1_full = _readData_readDataQueue_fifo_1_full;
  wire               readData_readDataQueue_2_empty;
  assign readData_readDataQueue_2_empty = _readData_readDataQueue_fifo_2_empty;
  wire               readData_readDataQueue_2_full;
  assign readData_readDataQueue_2_full = _readData_readDataQueue_fifo_2_full;
  wire               readData_readDataQueue_3_empty;
  assign readData_readDataQueue_3_empty = _readData_readDataQueue_fifo_3_empty;
  wire               readData_readDataQueue_3_full;
  assign readData_readDataQueue_3_full = _readData_readDataQueue_fifo_3_full;
  assign compressUnitResultQueue_enq_valid = _compressUnit_out_compressValid;
  assign compressUnitResultQueue_enq_bits_compressValid = _compressUnit_out_compressValid;
  wire               writeQueue_0_empty;
  assign writeQueue_0_empty = _writeQueue_fifo_empty;
  wire               writeQueue_0_full;
  assign writeQueue_0_full = _writeQueue_fifo_full;
  wire               writeQueue_1_empty;
  assign writeQueue_1_empty = _writeQueue_fifo_1_empty;
  wire               writeQueue_1_full;
  assign writeQueue_1_full = _writeQueue_fifo_1_full;
  wire               writeQueue_2_empty;
  assign writeQueue_2_empty = _writeQueue_fifo_2_empty;
  wire               writeQueue_2_full;
  assign writeQueue_2_full = _writeQueue_fifo_2_full;
  wire               writeQueue_3_empty;
  assign writeQueue_3_empty = _writeQueue_fifo_3_empty;
  wire               writeQueue_3_full;
  assign writeQueue_3_full = _writeQueue_fifo_3_full;
  BitLevelMaskWrite maskedWrite (
    .clock                             (clock),
    .reset                             (reset),
    .needWAR                           (maskDestinationType),
    .vd                                (instReg_vd),
    .in_0_ready                        (_maskedWrite_in_0_ready),
    .in_0_valid                        (unitType[2] ? _reduceUnit_out_valid : executeValid & maskFilter),
    .in_0_bits_data                    (unitType[2] ? _reduceUnit_out_bits_data : executeResult[31:0]),
    .in_0_bits_bitMask                 (currentMaskGroupForDestination[31:0]),
    .in_0_bits_mask                    (unitType[2] ? _reduceUnit_out_bits_mask : executeWriteByteMask[3:0]),
    .in_0_bits_groupCounter            (unitType[2] ? 10'h0 : executeDeqGroupCounter[9:0]),
    .in_0_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[0] & ffo),
    .in_1_ready                        (_maskedWrite_in_1_ready),
    .in_1_valid                        (executeValid & maskFilter_1),
    .in_1_bits_data                    (executeResult[63:32]),
    .in_1_bits_bitMask                 (currentMaskGroupForDestination[63:32]),
    .in_1_bits_mask                    (executeWriteByteMask[7:4]),
    .in_1_bits_groupCounter            (executeDeqGroupCounter[9:0]),
    .in_1_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[1] & ffo),
    .in_2_ready                        (_maskedWrite_in_2_ready),
    .in_2_valid                        (executeValid & maskFilter_2),
    .in_2_bits_data                    (executeResult[95:64]),
    .in_2_bits_bitMask                 (currentMaskGroupForDestination[95:64]),
    .in_2_bits_mask                    (executeWriteByteMask[11:8]),
    .in_2_bits_groupCounter            (executeDeqGroupCounter[9:0]),
    .in_2_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[2] & ffo),
    .in_3_ready                        (_maskedWrite_in_3_ready),
    .in_3_valid                        (executeValid & maskFilter_3),
    .in_3_bits_data                    (executeResult[127:96]),
    .in_3_bits_bitMask                 (currentMaskGroupForDestination[127:96]),
    .in_3_bits_mask                    (executeWriteByteMask[15:12]),
    .in_3_bits_groupCounter            (executeDeqGroupCounter[9:0]),
    .in_3_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[3] & ffo),
    .out_0_ready                       (writeQueue_0_enq_ready),
    .out_0_valid                       (_maskedWrite_out_0_valid),
    .out_0_bits_ffoByOther             (_maskedWrite_out_0_bits_ffoByOther),
    .out_0_bits_writeData_data         (_maskedWrite_out_0_bits_writeData_data),
    .out_0_bits_writeData_mask         (_maskedWrite_out_0_bits_writeData_mask),
    .out_0_bits_writeData_groupCounter (_maskedWrite_out_0_bits_writeData_groupCounter),
    .out_1_ready                       (writeQueue_1_enq_ready),
    .out_1_valid                       (_maskedWrite_out_1_valid),
    .out_1_bits_ffoByOther             (_maskedWrite_out_1_bits_ffoByOther),
    .out_1_bits_writeData_data         (_maskedWrite_out_1_bits_writeData_data),
    .out_1_bits_writeData_mask         (_maskedWrite_out_1_bits_writeData_mask),
    .out_1_bits_writeData_groupCounter (_maskedWrite_out_1_bits_writeData_groupCounter),
    .out_2_ready                       (writeQueue_2_enq_ready),
    .out_2_valid                       (_maskedWrite_out_2_valid),
    .out_2_bits_ffoByOther             (_maskedWrite_out_2_bits_ffoByOther),
    .out_2_bits_writeData_data         (_maskedWrite_out_2_bits_writeData_data),
    .out_2_bits_writeData_mask         (_maskedWrite_out_2_bits_writeData_mask),
    .out_2_bits_writeData_groupCounter (_maskedWrite_out_2_bits_writeData_groupCounter),
    .out_3_ready                       (writeQueue_3_enq_ready),
    .out_3_valid                       (_maskedWrite_out_3_valid),
    .out_3_bits_ffoByOther             (_maskedWrite_out_3_bits_ffoByOther),
    .out_3_bits_writeData_data         (_maskedWrite_out_3_bits_writeData_data),
    .out_3_bits_writeData_mask         (_maskedWrite_out_3_bits_writeData_mask),
    .out_3_bits_writeData_groupCounter (_maskedWrite_out_3_bits_writeData_groupCounter),
    .readChannel_0_ready               (readChannel_0_ready_0),
    .readChannel_0_valid               (_maskedWrite_readChannel_0_valid),
    .readChannel_0_bits_vs             (_maskedWrite_readChannel_0_bits_vs),
    .readChannel_0_bits_offset         (_maskedWrite_readChannel_0_bits_offset),
    .readChannel_1_ready               (readChannel_1_ready_0),
    .readChannel_1_valid               (_maskedWrite_readChannel_1_valid),
    .readChannel_1_bits_vs             (_maskedWrite_readChannel_1_bits_vs),
    .readChannel_1_bits_offset         (_maskedWrite_readChannel_1_bits_offset),
    .readChannel_2_ready               (readChannel_2_ready_0),
    .readChannel_2_valid               (_maskedWrite_readChannel_2_valid),
    .readChannel_2_bits_vs             (_maskedWrite_readChannel_2_bits_vs),
    .readChannel_2_bits_offset         (_maskedWrite_readChannel_2_bits_offset),
    .readChannel_3_ready               (readChannel_3_ready_0),
    .readChannel_3_valid               (_maskedWrite_readChannel_3_valid),
    .readChannel_3_bits_vs             (_maskedWrite_readChannel_3_bits_vs),
    .readChannel_3_bits_offset         (_maskedWrite_readChannel_3_bits_offset),
    .readResult_0_valid                (readResult_0_valid),
    .readResult_0_bits                 (readResult_0_bits),
    .readResult_1_valid                (readResult_1_valid),
    .readResult_1_bits                 (readResult_1_bits),
    .readResult_2_valid                (readResult_2_valid),
    .readResult_2_bits                 (readResult_2_bits),
    .readResult_3_valid                (readResult_3_valid),
    .readResult_3_bits                 (readResult_3_bits),
    .stageClear                        (_maskedWrite_stageClear)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_0_enq_ready & exeRequestQueue_0_enq_valid & ~(_exeRequestQueue_queue_fifo_empty & exeRequestQueue_0_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_0_deq_ready & ~_exeRequestQueue_queue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn),
    .empty        (_exeRequestQueue_queue_fifo_empty),
    .almost_empty (exeRequestQueue_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_0_almostFull),
    .full         (_exeRequestQueue_queue_fifo_full),
    .error        (_exeRequestQueue_queue_fifo_error),
    .data_out     (_exeRequestQueue_queue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_1_enq_ready & exeRequestQueue_1_enq_valid & ~(_exeRequestQueue_queue_fifo_1_empty & exeRequestQueue_1_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_1_deq_ready & ~_exeRequestQueue_queue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_1),
    .empty        (_exeRequestQueue_queue_fifo_1_empty),
    .almost_empty (exeRequestQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_1_almostFull),
    .full         (_exeRequestQueue_queue_fifo_1_full),
    .error        (_exeRequestQueue_queue_fifo_1_error),
    .data_out     (_exeRequestQueue_queue_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_2_enq_ready & exeRequestQueue_2_enq_valid & ~(_exeRequestQueue_queue_fifo_2_empty & exeRequestQueue_2_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_2_deq_ready & ~_exeRequestQueue_queue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_2),
    .empty        (_exeRequestQueue_queue_fifo_2_empty),
    .almost_empty (exeRequestQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_2_almostFull),
    .full         (_exeRequestQueue_queue_fifo_2_full),
    .error        (_exeRequestQueue_queue_fifo_2_error),
    .data_out     (_exeRequestQueue_queue_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_3_enq_ready & exeRequestQueue_3_enq_valid & ~(_exeRequestQueue_queue_fifo_3_empty & exeRequestQueue_3_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_3_deq_ready & ~_exeRequestQueue_queue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_3),
    .empty        (_exeRequestQueue_queue_fifo_3_empty),
    .almost_empty (exeRequestQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_3_almostFull),
    .full         (_exeRequestQueue_queue_fifo_3_full),
    .error        (_exeRequestQueue_queue_fifo_3_error),
    .data_out     (_exeRequestQueue_queue_fifo_3_data_out)
  );
  SlideIndexGen slideAddressGen (
    .clock                              (clock),
    .reset                              (reset),
    .newInstruction                     (instReq_valid & (|instReq_bits_vl)),
    .instructionReq_decodeResult_topUop (instReg_decodeResult_topUop),
    .instructionReq_readFromScala       (instReg_readFromScala),
    .instructionReq_sew                 (instReg_sew),
    .instructionReq_vlmul               (instReg_vlmul),
    .instructionReq_maskType            (instReg_maskType),
    .instructionReq_vl                  (instReg_vl),
    .indexDeq_ready                     (slideAddressGen_indexDeq_ready),
    .indexDeq_valid                     (_slideAddressGen_indexDeq_valid),
    .indexDeq_bits_needRead             (_slideAddressGen_indexDeq_bits_needRead),
    .indexDeq_bits_elementValid         (_slideAddressGen_indexDeq_bits_elementValid),
    .indexDeq_bits_replaceVs1           (_slideAddressGen_indexDeq_bits_replaceVs1),
    .indexDeq_bits_readOffset           (_slideAddressGen_indexDeq_bits_readOffset),
    .indexDeq_bits_accessLane_0         (_slideAddressGen_indexDeq_bits_accessLane_0),
    .indexDeq_bits_accessLane_1         (_slideAddressGen_indexDeq_bits_accessLane_1),
    .indexDeq_bits_accessLane_2         (_slideAddressGen_indexDeq_bits_accessLane_2),
    .indexDeq_bits_accessLane_3         (_slideAddressGen_indexDeq_bits_accessLane_3),
    .indexDeq_bits_vsGrowth_0           (_slideAddressGen_indexDeq_bits_vsGrowth_0),
    .indexDeq_bits_vsGrowth_1           (_slideAddressGen_indexDeq_bits_vsGrowth_1),
    .indexDeq_bits_vsGrowth_2           (_slideAddressGen_indexDeq_bits_vsGrowth_2),
    .indexDeq_bits_vsGrowth_3           (_slideAddressGen_indexDeq_bits_vsGrowth_3),
    .indexDeq_bits_executeGroup         (_slideAddressGen_indexDeq_bits_executeGroup),
    .indexDeq_bits_readDataOffset       (_slideAddressGen_indexDeq_bits_readDataOffset),
    .indexDeq_bits_last                 (_slideAddressGen_indexDeq_bits_last),
    .slideGroupOut                      (_slideAddressGen_slideGroupOut),
    .slideMaskInput                     (_GEN_140[_slideAddressGen_slideGroupOut[10:0]])
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) accessCountQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(accessCountQueue_enq_ready & accessCountQueue_enq_valid)),
    .pop_req_n    (~(accessCountQueue_deq_ready & ~_accessCountQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (accessCountQueue_dataIn),
    .empty        (_accessCountQueue_fifo_empty),
    .almost_empty (accessCountQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (accessCountQueue_almostFull),
    .full         (_accessCountQueue_fifo_full),
    .error        (_accessCountQueue_fifo_error),
    .data_out     (_accessCountQueue_fifo_data_out)
  );
  MaskUnitReadCrossBar readCrossBar (
    .input_0_ready            (_readCrossBar_input_0_ready),
    .input_0_valid            (readCrossBar_input_0_valid),
    .input_0_bits_vs          (selectExecuteReq_0_bits_vs),
    .input_0_bits_offset      (selectExecuteReq_0_bits_offset),
    .input_0_bits_readLane    (selectExecuteReq_0_bits_readLane),
    .input_0_bits_dataOffset  (selectExecuteReq_0_bits_dataOffset),
    .input_1_ready            (_readCrossBar_input_1_ready),
    .input_1_valid            (readCrossBar_input_1_valid),
    .input_1_bits_vs          (selectExecuteReq_1_bits_vs),
    .input_1_bits_offset      (selectExecuteReq_1_bits_offset),
    .input_1_bits_readLane    (selectExecuteReq_1_bits_readLane),
    .input_1_bits_dataOffset  (selectExecuteReq_1_bits_dataOffset),
    .input_2_ready            (_readCrossBar_input_2_ready),
    .input_2_valid            (readCrossBar_input_2_valid),
    .input_2_bits_vs          (selectExecuteReq_2_bits_vs),
    .input_2_bits_offset      (selectExecuteReq_2_bits_offset),
    .input_2_bits_readLane    (selectExecuteReq_2_bits_readLane),
    .input_2_bits_dataOffset  (selectExecuteReq_2_bits_dataOffset),
    .input_3_ready            (_readCrossBar_input_3_ready),
    .input_3_valid            (readCrossBar_input_3_valid),
    .input_3_bits_vs          (selectExecuteReq_3_bits_vs),
    .input_3_bits_offset      (selectExecuteReq_3_bits_offset),
    .input_3_bits_readLane    (selectExecuteReq_3_bits_readLane),
    .input_3_bits_dataOffset  (selectExecuteReq_3_bits_dataOffset),
    .output_0_ready           (readChannel_0_ready_0 & readMessageQueue_enq_ready),
    .output_0_valid           (_readCrossBar_output_0_valid),
    .output_0_bits_vs         (_readCrossBar_output_0_bits_vs),
    .output_0_bits_offset     (_readCrossBar_output_0_bits_offset),
    .output_0_bits_writeIndex (_readCrossBar_output_0_bits_writeIndex),
    .output_0_bits_dataOffset (readMessageQueue_enq_bits_dataOffset),
    .output_1_ready           (readChannel_1_ready_0 & readMessageQueue_1_enq_ready),
    .output_1_valid           (_readCrossBar_output_1_valid),
    .output_1_bits_vs         (_readCrossBar_output_1_bits_vs),
    .output_1_bits_offset     (_readCrossBar_output_1_bits_offset),
    .output_1_bits_writeIndex (_readCrossBar_output_1_bits_writeIndex),
    .output_1_bits_dataOffset (readMessageQueue_1_enq_bits_dataOffset),
    .output_2_ready           (readChannel_2_ready_0 & readMessageQueue_2_enq_ready),
    .output_2_valid           (_readCrossBar_output_2_valid),
    .output_2_bits_vs         (_readCrossBar_output_2_bits_vs),
    .output_2_bits_offset     (_readCrossBar_output_2_bits_offset),
    .output_2_bits_writeIndex (_readCrossBar_output_2_bits_writeIndex),
    .output_2_bits_dataOffset (readMessageQueue_2_enq_bits_dataOffset),
    .output_3_ready           (readChannel_3_ready_0 & readMessageQueue_3_enq_ready),
    .output_3_valid           (_readCrossBar_output_3_valid),
    .output_3_bits_vs         (_readCrossBar_output_3_bits_vs),
    .output_3_bits_offset     (_readCrossBar_output_3_bits_offset),
    .output_3_bits_writeIndex (_readCrossBar_output_3_bits_writeIndex),
    .output_3_bits_dataOffset (readMessageQueue_3_enq_bits_dataOffset)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(25)
  ) readWaitQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readWaitQueue_enq_ready & readWaitQueue_enq_valid)),
    .pop_req_n    (~(readWaitQueue_deq_ready & ~_readWaitQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (readWaitQueue_dataIn),
    .empty        (_readWaitQueue_fifo_empty),
    .almost_empty (readWaitQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readWaitQueue_almostFull),
    .full         (_readWaitQueue_fifo_full),
    .error        (_readWaitQueue_fifo_error),
    .data_out     (_readWaitQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(159)
  ) compressUnitResultQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(compressUnitResultQueue_enq_ready & compressUnitResultQueue_enq_valid & ~(_compressUnitResultQueue_fifo_empty & compressUnitResultQueue_deq_ready))),
    .pop_req_n    (~(compressUnitResultQueue_deq_ready & ~_compressUnitResultQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (compressUnitResultQueue_dataIn),
    .empty        (_compressUnitResultQueue_fifo_empty),
    .almost_empty (compressUnitResultQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (compressUnitResultQueue_almostFull),
    .full         (_compressUnitResultQueue_fifo_full),
    .error        (_compressUnitResultQueue_fifo_error),
    .data_out     (_compressUnitResultQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(36)
  ) reorderQueueVec_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_0_enq_ready & reorderQueueVec_0_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_0_deq_ready & ~_reorderQueueVec_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn),
    .empty        (_reorderQueueVec_fifo_empty),
    .almost_empty (reorderQueueVec_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_0_almostFull),
    .full         (_reorderQueueVec_fifo_full),
    .error        (_reorderQueueVec_fifo_error),
    .data_out     (_reorderQueueVec_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(36)
  ) reorderQueueVec_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_1_enq_ready & reorderQueueVec_1_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_1_deq_ready & ~_reorderQueueVec_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_1),
    .empty        (_reorderQueueVec_fifo_1_empty),
    .almost_empty (reorderQueueVec_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_1_almostFull),
    .full         (_reorderQueueVec_fifo_1_full),
    .error        (_reorderQueueVec_fifo_1_error),
    .data_out     (_reorderQueueVec_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(36)
  ) reorderQueueVec_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_2_enq_ready & reorderQueueVec_2_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_2_deq_ready & ~_reorderQueueVec_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_2),
    .empty        (_reorderQueueVec_fifo_2_empty),
    .almost_empty (reorderQueueVec_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_2_almostFull),
    .full         (_reorderQueueVec_fifo_2_full),
    .error        (_reorderQueueVec_fifo_2_error),
    .data_out     (_reorderQueueVec_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(36)
  ) reorderQueueVec_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_3_enq_ready & reorderQueueVec_3_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_3_deq_ready & ~_reorderQueueVec_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_3),
    .empty        (_reorderQueueVec_fifo_3_empty),
    .almost_empty (reorderQueueVec_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_3_almostFull),
    .full         (_reorderQueueVec_fifo_3_full),
    .error        (_reorderQueueVec_fifo_3_error),
    .data_out     (_reorderQueueVec_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(6)
  ) readMessageQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_enq_ready & readMessageQueue_enq_valid)),
    .pop_req_n    (~(readMessageQueue_deq_ready & ~_readMessageQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn),
    .empty        (_readMessageQueue_fifo_empty),
    .almost_empty (readMessageQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_almostFull),
    .full         (_readMessageQueue_fifo_full),
    .error        (_readMessageQueue_fifo_error),
    .data_out     (_readMessageQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(6)
  ) readMessageQueue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_1_enq_ready & readMessageQueue_1_enq_valid)),
    .pop_req_n    (~(readMessageQueue_1_deq_ready & ~_readMessageQueue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_1),
    .empty        (_readMessageQueue_fifo_1_empty),
    .almost_empty (readMessageQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_1_almostFull),
    .full         (_readMessageQueue_fifo_1_full),
    .error        (_readMessageQueue_fifo_1_error),
    .data_out     (_readMessageQueue_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(6)
  ) readMessageQueue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_2_enq_ready & readMessageQueue_2_enq_valid)),
    .pop_req_n    (~(readMessageQueue_2_deq_ready & ~_readMessageQueue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_2),
    .empty        (_readMessageQueue_fifo_2_empty),
    .almost_empty (readMessageQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_2_almostFull),
    .full         (_readMessageQueue_fifo_2_full),
    .error        (_readMessageQueue_fifo_2_error),
    .data_out     (_readMessageQueue_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(6)
  ) readMessageQueue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_3_enq_ready & readMessageQueue_3_enq_valid)),
    .pop_req_n    (~(readMessageQueue_3_deq_ready & ~_readMessageQueue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_3),
    .empty        (_readMessageQueue_fifo_3_empty),
    .almost_empty (readMessageQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_3_almostFull),
    .full         (_readMessageQueue_fifo_3_full),
    .error        (_readMessageQueue_fifo_3_error),
    .data_out     (_readMessageQueue_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_enq_ready & readData_readDataQueue_enq_valid & ~(_readData_readDataQueue_fifo_empty & readData_readDataQueue_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_deq_ready & ~_readData_readDataQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_enq_bits),
    .empty        (_readData_readDataQueue_fifo_empty),
    .almost_empty (readData_readDataQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_almostFull),
    .full         (_readData_readDataQueue_fifo_full),
    .error        (_readData_readDataQueue_fifo_error),
    .data_out     (_readData_readDataQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_1_enq_ready & readData_readDataQueue_1_enq_valid & ~(_readData_readDataQueue_fifo_1_empty & readData_readDataQueue_1_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_1_deq_ready & ~_readData_readDataQueue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_1_enq_bits),
    .empty        (_readData_readDataQueue_fifo_1_empty),
    .almost_empty (readData_readDataQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_1_almostFull),
    .full         (_readData_readDataQueue_fifo_1_full),
    .error        (_readData_readDataQueue_fifo_1_error),
    .data_out     (_readData_readDataQueue_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_2_enq_ready & readData_readDataQueue_2_enq_valid & ~(_readData_readDataQueue_fifo_2_empty & readData_readDataQueue_2_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_2_deq_ready & ~_readData_readDataQueue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_2_enq_bits),
    .empty        (_readData_readDataQueue_fifo_2_empty),
    .almost_empty (readData_readDataQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_2_almostFull),
    .full         (_readData_readDataQueue_fifo_2_full),
    .error        (_readData_readDataQueue_fifo_2_error),
    .data_out     (_readData_readDataQueue_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_3_enq_ready & readData_readDataQueue_3_enq_valid & ~(_readData_readDataQueue_fifo_3_empty & readData_readDataQueue_3_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_3_deq_ready & ~_readData_readDataQueue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_3_enq_bits),
    .empty        (_readData_readDataQueue_fifo_3_empty),
    .almost_empty (readData_readDataQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_3_almostFull),
    .full         (_readData_readDataQueue_fifo_3_full),
    .error        (_readData_readDataQueue_fifo_3_error),
    .data_out     (_readData_readDataQueue_fifo_3_data_out)
  );
  MaskCompress compressUnit (
    .clock                  (clock),
    .reset                  (reset),
    .in_valid               (viotaCounterAdd),
    .in_bits_maskType       (instReg_maskType),
    .in_bits_eew            (instReg_sew),
    .in_bits_uop            (instReg_decodeResult_topUop[2:0]),
    .in_bits_readFromScalar (instReg_readFromScala),
    .in_bits_source1        (source1Select),
    .in_bits_mask           ({16'h0, executeElementMask}),
    .in_bits_source2        (source2),
    .in_bits_pipeData       (source1),
    .in_bits_groupCounter   (requestCounter),
    .in_bits_ffoInput       ({view__in_bits_ffoInput_hi, view__in_bits_ffoInput_lo}),
    .in_bits_validInput     ({view__in_bits_validInput_hi, view__in_bits_validInput_lo}),
    .in_bits_lastCompress   (lastGroup),
    .out_data               (compressUnitResultQueue_enq_bits_data),
    .out_mask               (compressUnitResultQueue_enq_bits_mask),
    .out_groupCounter       (compressUnitResultQueue_enq_bits_groupCounter),
    .out_ffoOutput          (compressUnitResultQueue_enq_bits_ffoOutput),
    .out_compressValid      (_compressUnit_out_compressValid),
    .newInstruction         (instReq_valid),
    .ffoInstruction         (&(instReq_bits_decodeResult_topUop[2:1])),
    .writeData              (_compressUnit_writeData),
    .stageValid             (_compressUnit_stageValid)
  );
  MaskReduce reduceUnit (
    .clock               (clock),
    .reset               (reset),
    .in_ready            (_reduceUnit_in_ready),
    .in_valid            (reduceUnit_in_valid),
    .in_bits_maskType    (instReg_maskType),
    .in_bits_eew         (instReg_sew),
    .in_bits_uop         (instReg_decodeResult_topUop[2:0]),
    .in_bits_readVS1     (readVS1Reg_data),
    .in_bits_source2     (source2),
    .in_bits_sourceValid ({view__in_bits_sourceValid_hi, view__in_bits_sourceValid_lo}),
    .in_bits_lastGroup   (lastGroup),
    .in_bits_vxrm        (instReg_vxrm),
    .in_bits_aluUop      (instReg_decodeResult_uop),
    .in_bits_sign        (~instReg_decodeResult_unsigned1),
    .out_valid           (_reduceUnit_out_valid),
    .out_bits_data       (_reduceUnit_out_bits_data),
    .out_bits_mask       (_reduceUnit_out_bits_mask),
    .firstGroup          (~readVS1Reg_sendToExecution & _view__firstGroup_T_1),
    .newInstruction      (instReq_valid),
    .validInst           (|instReg_vl),
    .pop                 (instReg_decodeResult_popCount)
  );
  MaskExtend extendUnit (
    .in_eew          (instReg_sew),
    .in_uop          (instReg_decodeResult_topUop[2:0]),
    .in_source2      (source2),
    .in_groupCounter (extendGroupCount[9:0]),
    .out             (_extendUnit_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(55)
  ) writeQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_0_enq_ready & writeQueue_0_enq_valid)),
    .pop_req_n    (~(writeQueue_0_deq_ready & ~_writeQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn),
    .empty        (_writeQueue_fifo_empty),
    .almost_empty (writeQueue_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_0_almostFull),
    .full         (_writeQueue_fifo_full),
    .error        (_writeQueue_fifo_error),
    .data_out     (_writeQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(55)
  ) writeQueue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_1_enq_ready & writeQueue_1_enq_valid)),
    .pop_req_n    (~(writeQueue_1_deq_ready & ~_writeQueue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_1),
    .empty        (_writeQueue_fifo_1_empty),
    .almost_empty (writeQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_1_almostFull),
    .full         (_writeQueue_fifo_1_full),
    .error        (_writeQueue_fifo_1_error),
    .data_out     (_writeQueue_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(55)
  ) writeQueue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_2_enq_ready & writeQueue_2_enq_valid)),
    .pop_req_n    (~(writeQueue_2_deq_ready & ~_writeQueue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_2),
    .empty        (_writeQueue_fifo_2_empty),
    .almost_empty (writeQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_2_almostFull),
    .full         (_writeQueue_fifo_2_full),
    .error        (_writeQueue_fifo_2_error),
    .data_out     (_writeQueue_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(55)
  ) writeQueue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_3_enq_ready & writeQueue_3_enq_valid)),
    .pop_req_n    (~(writeQueue_3_deq_ready & ~_writeQueue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_3),
    .empty        (_writeQueue_fifo_3_empty),
    .almost_empty (writeQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_3_almostFull),
    .full         (_writeQueue_fifo_3_full),
    .error        (_writeQueue_fifo_3_error),
    .data_out     (_writeQueue_fifo_3_data_out)
  );
  assign exeResp_0_valid = exeResp_0_valid_0;
  assign exeResp_0_bits_vd = exeResp_0_bits_vd_0;
  assign exeResp_0_bits_offset = exeResp_0_bits_offset_0;
  assign exeResp_0_bits_mask = exeResp_0_bits_mask_0;
  assign exeResp_0_bits_data = exeResp_0_bits_data_0;
  assign exeResp_0_bits_instructionIndex = exeResp_0_bits_instructionIndex_0;
  assign exeResp_1_valid = exeResp_1_valid_0;
  assign exeResp_1_bits_vd = exeResp_1_bits_vd_0;
  assign exeResp_1_bits_offset = exeResp_1_bits_offset_0;
  assign exeResp_1_bits_mask = exeResp_1_bits_mask_0;
  assign exeResp_1_bits_data = exeResp_1_bits_data_0;
  assign exeResp_1_bits_instructionIndex = exeResp_1_bits_instructionIndex_0;
  assign exeResp_2_valid = exeResp_2_valid_0;
  assign exeResp_2_bits_vd = exeResp_2_bits_vd_0;
  assign exeResp_2_bits_offset = exeResp_2_bits_offset_0;
  assign exeResp_2_bits_mask = exeResp_2_bits_mask_0;
  assign exeResp_2_bits_data = exeResp_2_bits_data_0;
  assign exeResp_2_bits_instructionIndex = exeResp_2_bits_instructionIndex_0;
  assign exeResp_3_valid = exeResp_3_valid_0;
  assign exeResp_3_bits_vd = exeResp_3_bits_vd_0;
  assign exeResp_3_bits_offset = exeResp_3_bits_offset_0;
  assign exeResp_3_bits_mask = exeResp_3_bits_mask_0;
  assign exeResp_3_bits_data = exeResp_3_bits_data_0;
  assign exeResp_3_bits_instructionIndex = exeResp_3_bits_instructionIndex_0;
  assign tokenIO_0_maskRequestRelease = tokenIO_0_maskRequestRelease_0;
  assign tokenIO_1_maskRequestRelease = tokenIO_1_maskRequestRelease_0;
  assign tokenIO_2_maskRequestRelease = tokenIO_2_maskRequestRelease_0;
  assign tokenIO_3_maskRequestRelease = tokenIO_3_maskRequestRelease_0;
  assign readChannel_0_valid = readChannel_0_valid_0;
  assign readChannel_0_bits_vs = readChannel_0_bits_vs_0;
  assign readChannel_0_bits_offset = readChannel_0_bits_offset_0;
  assign readChannel_0_bits_instructionIndex = readChannel_0_bits_instructionIndex_0;
  assign readChannel_1_valid = readChannel_1_valid_0;
  assign readChannel_1_bits_vs = readChannel_1_bits_vs_0;
  assign readChannel_1_bits_offset = readChannel_1_bits_offset_0;
  assign readChannel_1_bits_instructionIndex = readChannel_1_bits_instructionIndex_0;
  assign readChannel_2_valid = readChannel_2_valid_0;
  assign readChannel_2_bits_vs = readChannel_2_bits_vs_0;
  assign readChannel_2_bits_offset = readChannel_2_bits_offset_0;
  assign readChannel_2_bits_instructionIndex = readChannel_2_bits_instructionIndex_0;
  assign readChannel_3_valid = readChannel_3_valid_0;
  assign readChannel_3_bits_vs = readChannel_3_bits_vs_0;
  assign readChannel_3_bits_offset = readChannel_3_bits_offset_0;
  assign readChannel_3_bits_instructionIndex = readChannel_3_bits_instructionIndex_0;
  assign lastReport = _lastReport_output;
  assign laneMaskInput_0 = _GEN_127[laneMaskSelect_0[5:0]];
  assign laneMaskInput_1 = _GEN_128[laneMaskSelect_1[5:0]];
  assign laneMaskInput_2 = _GEN_129[laneMaskSelect_2[5:0]];
  assign laneMaskInput_3 = _GEN_130[laneMaskSelect_3[5:0]];
  assign writeRDData = instReg_decodeResult_popCount ? _reduceUnit_out_bits_data : _compressUnit_writeData;
  assign gatherData_valid = gatherData_valid_0;
  assign gatherData_bits = gatherData_bits_0;
endmodule

